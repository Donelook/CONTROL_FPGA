// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Oct 16 2025 00:42:38

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    s4_phy,
    rgb_g,
    start_stop,
    s2_phy,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output s4_phy;
    output rgb_g;
    input start_stop;
    output s2_phy;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__21137;
    wire N__21136;
    wire N__21135;
    wire N__21126;
    wire N__21125;
    wire N__21124;
    wire N__21117;
    wire N__21116;
    wire N__21115;
    wire N__21108;
    wire N__21107;
    wire N__21106;
    wire N__21099;
    wire N__21098;
    wire N__21097;
    wire N__21090;
    wire N__21089;
    wire N__21088;
    wire N__21081;
    wire N__21080;
    wire N__21079;
    wire N__21072;
    wire N__21071;
    wire N__21070;
    wire N__21063;
    wire N__21062;
    wire N__21061;
    wire N__21054;
    wire N__21053;
    wire N__21052;
    wire N__21045;
    wire N__21044;
    wire N__21043;
    wire N__21036;
    wire N__21035;
    wire N__21034;
    wire N__21027;
    wire N__21026;
    wire N__21025;
    wire N__21008;
    wire N__21005;
    wire N__21004;
    wire N__21003;
    wire N__21000;
    wire N__20997;
    wire N__20994;
    wire N__20987;
    wire N__20984;
    wire N__20983;
    wire N__20982;
    wire N__20979;
    wire N__20976;
    wire N__20973;
    wire N__20966;
    wire N__20965;
    wire N__20964;
    wire N__20959;
    wire N__20956;
    wire N__20955;
    wire N__20950;
    wire N__20947;
    wire N__20942;
    wire N__20941;
    wire N__20940;
    wire N__20939;
    wire N__20938;
    wire N__20937;
    wire N__20936;
    wire N__20935;
    wire N__20934;
    wire N__20933;
    wire N__20932;
    wire N__20931;
    wire N__20930;
    wire N__20929;
    wire N__20928;
    wire N__20927;
    wire N__20926;
    wire N__20925;
    wire N__20924;
    wire N__20923;
    wire N__20922;
    wire N__20921;
    wire N__20920;
    wire N__20919;
    wire N__20918;
    wire N__20917;
    wire N__20916;
    wire N__20915;
    wire N__20914;
    wire N__20913;
    wire N__20912;
    wire N__20911;
    wire N__20910;
    wire N__20909;
    wire N__20908;
    wire N__20907;
    wire N__20906;
    wire N__20905;
    wire N__20904;
    wire N__20903;
    wire N__20902;
    wire N__20901;
    wire N__20900;
    wire N__20899;
    wire N__20898;
    wire N__20897;
    wire N__20896;
    wire N__20895;
    wire N__20894;
    wire N__20893;
    wire N__20892;
    wire N__20891;
    wire N__20890;
    wire N__20889;
    wire N__20888;
    wire N__20887;
    wire N__20886;
    wire N__20885;
    wire N__20884;
    wire N__20883;
    wire N__20882;
    wire N__20881;
    wire N__20880;
    wire N__20879;
    wire N__20878;
    wire N__20877;
    wire N__20876;
    wire N__20875;
    wire N__20874;
    wire N__20873;
    wire N__20872;
    wire N__20871;
    wire N__20870;
    wire N__20869;
    wire N__20868;
    wire N__20867;
    wire N__20866;
    wire N__20865;
    wire N__20864;
    wire N__20705;
    wire N__20702;
    wire N__20699;
    wire N__20696;
    wire N__20693;
    wire N__20692;
    wire N__20689;
    wire N__20686;
    wire N__20681;
    wire N__20680;
    wire N__20679;
    wire N__20674;
    wire N__20671;
    wire N__20668;
    wire N__20663;
    wire N__20660;
    wire N__20659;
    wire N__20658;
    wire N__20655;
    wire N__20652;
    wire N__20651;
    wire N__20648;
    wire N__20643;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20631;
    wire N__20628;
    wire N__20625;
    wire N__20622;
    wire N__20615;
    wire N__20614;
    wire N__20613;
    wire N__20612;
    wire N__20609;
    wire N__20602;
    wire N__20597;
    wire N__20596;
    wire N__20595;
    wire N__20594;
    wire N__20593;
    wire N__20592;
    wire N__20591;
    wire N__20590;
    wire N__20589;
    wire N__20588;
    wire N__20587;
    wire N__20586;
    wire N__20585;
    wire N__20584;
    wire N__20583;
    wire N__20582;
    wire N__20581;
    wire N__20580;
    wire N__20579;
    wire N__20578;
    wire N__20569;
    wire N__20560;
    wire N__20551;
    wire N__20542;
    wire N__20533;
    wire N__20532;
    wire N__20531;
    wire N__20530;
    wire N__20529;
    wire N__20528;
    wire N__20527;
    wire N__20526;
    wire N__20525;
    wire N__20524;
    wire N__20523;
    wire N__20518;
    wire N__20511;
    wire N__20506;
    wire N__20497;
    wire N__20488;
    wire N__20479;
    wire N__20476;
    wire N__20473;
    wire N__20468;
    wire N__20467;
    wire N__20466;
    wire N__20465;
    wire N__20464;
    wire N__20463;
    wire N__20462;
    wire N__20461;
    wire N__20458;
    wire N__20455;
    wire N__20452;
    wire N__20447;
    wire N__20444;
    wire N__20441;
    wire N__20438;
    wire N__20435;
    wire N__20432;
    wire N__20429;
    wire N__20426;
    wire N__20425;
    wire N__20424;
    wire N__20423;
    wire N__20422;
    wire N__20421;
    wire N__20420;
    wire N__20419;
    wire N__20418;
    wire N__20417;
    wire N__20416;
    wire N__20415;
    wire N__20414;
    wire N__20413;
    wire N__20412;
    wire N__20411;
    wire N__20410;
    wire N__20409;
    wire N__20408;
    wire N__20407;
    wire N__20406;
    wire N__20405;
    wire N__20402;
    wire N__20401;
    wire N__20400;
    wire N__20399;
    wire N__20398;
    wire N__20397;
    wire N__20396;
    wire N__20395;
    wire N__20394;
    wire N__20393;
    wire N__20392;
    wire N__20391;
    wire N__20390;
    wire N__20389;
    wire N__20386;
    wire N__20385;
    wire N__20384;
    wire N__20383;
    wire N__20382;
    wire N__20381;
    wire N__20380;
    wire N__20379;
    wire N__20378;
    wire N__20377;
    wire N__20376;
    wire N__20375;
    wire N__20374;
    wire N__20373;
    wire N__20372;
    wire N__20371;
    wire N__20370;
    wire N__20369;
    wire N__20368;
    wire N__20367;
    wire N__20366;
    wire N__20363;
    wire N__20362;
    wire N__20361;
    wire N__20360;
    wire N__20357;
    wire N__20356;
    wire N__20355;
    wire N__20354;
    wire N__20353;
    wire N__20352;
    wire N__20351;
    wire N__20350;
    wire N__20347;
    wire N__20346;
    wire N__20201;
    wire N__20198;
    wire N__20195;
    wire N__20192;
    wire N__20191;
    wire N__20190;
    wire N__20189;
    wire N__20188;
    wire N__20185;
    wire N__20182;
    wire N__20181;
    wire N__20178;
    wire N__20175;
    wire N__20172;
    wire N__20171;
    wire N__20168;
    wire N__20165;
    wire N__20162;
    wire N__20159;
    wire N__20156;
    wire N__20153;
    wire N__20150;
    wire N__20147;
    wire N__20144;
    wire N__20141;
    wire N__20136;
    wire N__20131;
    wire N__20128;
    wire N__20125;
    wire N__20122;
    wire N__20117;
    wire N__20114;
    wire N__20107;
    wire N__20102;
    wire N__20101;
    wire N__20098;
    wire N__20095;
    wire N__20090;
    wire N__20089;
    wire N__20088;
    wire N__20085;
    wire N__20082;
    wire N__20079;
    wire N__20072;
    wire N__20071;
    wire N__20070;
    wire N__20069;
    wire N__20066;
    wire N__20063;
    wire N__20060;
    wire N__20057;
    wire N__20048;
    wire N__20045;
    wire N__20042;
    wire N__20039;
    wire N__20036;
    wire N__20033;
    wire N__20030;
    wire N__20027;
    wire N__20024;
    wire N__20021;
    wire N__20018;
    wire N__20015;
    wire N__20012;
    wire N__20011;
    wire N__20010;
    wire N__20009;
    wire N__20006;
    wire N__20003;
    wire N__19998;
    wire N__19991;
    wire N__19990;
    wire N__19989;
    wire N__19986;
    wire N__19983;
    wire N__19980;
    wire N__19973;
    wire N__19972;
    wire N__19971;
    wire N__19968;
    wire N__19965;
    wire N__19962;
    wire N__19955;
    wire N__19952;
    wire N__19949;
    wire N__19946;
    wire N__19943;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19928;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19915;
    wire N__19914;
    wire N__19911;
    wire N__19910;
    wire N__19907;
    wire N__19904;
    wire N__19901;
    wire N__19898;
    wire N__19893;
    wire N__19888;
    wire N__19883;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19868;
    wire N__19865;
    wire N__19862;
    wire N__19859;
    wire N__19856;
    wire N__19853;
    wire N__19850;
    wire N__19847;
    wire N__19844;
    wire N__19841;
    wire N__19838;
    wire N__19835;
    wire N__19832;
    wire N__19829;
    wire N__19828;
    wire N__19827;
    wire N__19826;
    wire N__19825;
    wire N__19824;
    wire N__19823;
    wire N__19822;
    wire N__19821;
    wire N__19810;
    wire N__19801;
    wire N__19798;
    wire N__19795;
    wire N__19790;
    wire N__19787;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19769;
    wire N__19766;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19754;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19735;
    wire N__19734;
    wire N__19731;
    wire N__19728;
    wire N__19725;
    wire N__19720;
    wire N__19715;
    wire N__19712;
    wire N__19711;
    wire N__19710;
    wire N__19707;
    wire N__19704;
    wire N__19701;
    wire N__19696;
    wire N__19691;
    wire N__19688;
    wire N__19687;
    wire N__19686;
    wire N__19683;
    wire N__19680;
    wire N__19677;
    wire N__19670;
    wire N__19667;
    wire N__19666;
    wire N__19665;
    wire N__19662;
    wire N__19659;
    wire N__19656;
    wire N__19649;
    wire N__19646;
    wire N__19645;
    wire N__19642;
    wire N__19639;
    wire N__19634;
    wire N__19633;
    wire N__19632;
    wire N__19629;
    wire N__19626;
    wire N__19623;
    wire N__19618;
    wire N__19613;
    wire N__19610;
    wire N__19609;
    wire N__19606;
    wire N__19603;
    wire N__19598;
    wire N__19597;
    wire N__19596;
    wire N__19593;
    wire N__19590;
    wire N__19587;
    wire N__19582;
    wire N__19577;
    wire N__19574;
    wire N__19571;
    wire N__19570;
    wire N__19569;
    wire N__19568;
    wire N__19567;
    wire N__19566;
    wire N__19563;
    wire N__19562;
    wire N__19561;
    wire N__19560;
    wire N__19559;
    wire N__19558;
    wire N__19557;
    wire N__19554;
    wire N__19553;
    wire N__19546;
    wire N__19543;
    wire N__19532;
    wire N__19527;
    wire N__19524;
    wire N__19521;
    wire N__19516;
    wire N__19509;
    wire N__19504;
    wire N__19501;
    wire N__19496;
    wire N__19495;
    wire N__19494;
    wire N__19493;
    wire N__19492;
    wire N__19481;
    wire N__19478;
    wire N__19475;
    wire N__19474;
    wire N__19473;
    wire N__19470;
    wire N__19465;
    wire N__19460;
    wire N__19459;
    wire N__19458;
    wire N__19455;
    wire N__19452;
    wire N__19449;
    wire N__19446;
    wire N__19441;
    wire N__19436;
    wire N__19433;
    wire N__19430;
    wire N__19429;
    wire N__19428;
    wire N__19425;
    wire N__19422;
    wire N__19419;
    wire N__19414;
    wire N__19409;
    wire N__19408;
    wire N__19405;
    wire N__19404;
    wire N__19401;
    wire N__19398;
    wire N__19395;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19379;
    wire N__19376;
    wire N__19375;
    wire N__19374;
    wire N__19371;
    wire N__19368;
    wire N__19365;
    wire N__19360;
    wire N__19355;
    wire N__19354;
    wire N__19351;
    wire N__19348;
    wire N__19347;
    wire N__19342;
    wire N__19339;
    wire N__19334;
    wire N__19331;
    wire N__19328;
    wire N__19327;
    wire N__19326;
    wire N__19323;
    wire N__19320;
    wire N__19317;
    wire N__19310;
    wire N__19309;
    wire N__19308;
    wire N__19305;
    wire N__19302;
    wire N__19299;
    wire N__19296;
    wire N__19293;
    wire N__19288;
    wire N__19283;
    wire N__19280;
    wire N__19277;
    wire N__19276;
    wire N__19275;
    wire N__19272;
    wire N__19269;
    wire N__19266;
    wire N__19259;
    wire N__19256;
    wire N__19255;
    wire N__19254;
    wire N__19251;
    wire N__19248;
    wire N__19245;
    wire N__19240;
    wire N__19235;
    wire N__19232;
    wire N__19231;
    wire N__19230;
    wire N__19227;
    wire N__19224;
    wire N__19221;
    wire N__19216;
    wire N__19211;
    wire N__19208;
    wire N__19207;
    wire N__19206;
    wire N__19203;
    wire N__19198;
    wire N__19193;
    wire N__19190;
    wire N__19189;
    wire N__19188;
    wire N__19185;
    wire N__19180;
    wire N__19175;
    wire N__19174;
    wire N__19173;
    wire N__19170;
    wire N__19167;
    wire N__19164;
    wire N__19159;
    wire N__19154;
    wire N__19153;
    wire N__19150;
    wire N__19147;
    wire N__19146;
    wire N__19145;
    wire N__19144;
    wire N__19141;
    wire N__19136;
    wire N__19131;
    wire N__19128;
    wire N__19125;
    wire N__19122;
    wire N__19117;
    wire N__19114;
    wire N__19109;
    wire N__19106;
    wire N__19105;
    wire N__19104;
    wire N__19101;
    wire N__19098;
    wire N__19095;
    wire N__19090;
    wire N__19085;
    wire N__19084;
    wire N__19081;
    wire N__19078;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19063;
    wire N__19062;
    wire N__19059;
    wire N__19056;
    wire N__19053;
    wire N__19046;
    wire N__19045;
    wire N__19042;
    wire N__19039;
    wire N__19036;
    wire N__19033;
    wire N__19028;
    wire N__19025;
    wire N__19024;
    wire N__19023;
    wire N__19020;
    wire N__19017;
    wire N__19014;
    wire N__19007;
    wire N__19004;
    wire N__19003;
    wire N__19000;
    wire N__18997;
    wire N__18992;
    wire N__18989;
    wire N__18986;
    wire N__18985;
    wire N__18984;
    wire N__18981;
    wire N__18978;
    wire N__18975;
    wire N__18970;
    wire N__18965;
    wire N__18964;
    wire N__18961;
    wire N__18958;
    wire N__18955;
    wire N__18952;
    wire N__18949;
    wire N__18946;
    wire N__18941;
    wire N__18938;
    wire N__18937;
    wire N__18936;
    wire N__18933;
    wire N__18930;
    wire N__18927;
    wire N__18922;
    wire N__18917;
    wire N__18916;
    wire N__18915;
    wire N__18912;
    wire N__18911;
    wire N__18910;
    wire N__18907;
    wire N__18902;
    wire N__18899;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18885;
    wire N__18882;
    wire N__18877;
    wire N__18872;
    wire N__18869;
    wire N__18868;
    wire N__18867;
    wire N__18864;
    wire N__18859;
    wire N__18854;
    wire N__18853;
    wire N__18852;
    wire N__18851;
    wire N__18846;
    wire N__18845;
    wire N__18840;
    wire N__18839;
    wire N__18838;
    wire N__18837;
    wire N__18834;
    wire N__18831;
    wire N__18828;
    wire N__18825;
    wire N__18820;
    wire N__18815;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18799;
    wire N__18796;
    wire N__18791;
    wire N__18788;
    wire N__18787;
    wire N__18782;
    wire N__18779;
    wire N__18778;
    wire N__18777;
    wire N__18776;
    wire N__18775;
    wire N__18774;
    wire N__18773;
    wire N__18772;
    wire N__18759;
    wire N__18754;
    wire N__18749;
    wire N__18748;
    wire N__18745;
    wire N__18742;
    wire N__18741;
    wire N__18736;
    wire N__18733;
    wire N__18728;
    wire N__18725;
    wire N__18722;
    wire N__18721;
    wire N__18718;
    wire N__18717;
    wire N__18714;
    wire N__18711;
    wire N__18708;
    wire N__18707;
    wire N__18704;
    wire N__18699;
    wire N__18696;
    wire N__18689;
    wire N__18688;
    wire N__18687;
    wire N__18684;
    wire N__18683;
    wire N__18682;
    wire N__18681;
    wire N__18680;
    wire N__18679;
    wire N__18678;
    wire N__18677;
    wire N__18676;
    wire N__18673;
    wire N__18670;
    wire N__18667;
    wire N__18664;
    wire N__18649;
    wire N__18648;
    wire N__18647;
    wire N__18644;
    wire N__18641;
    wire N__18634;
    wire N__18629;
    wire N__18620;
    wire N__18617;
    wire N__18616;
    wire N__18613;
    wire N__18612;
    wire N__18609;
    wire N__18606;
    wire N__18603;
    wire N__18600;
    wire N__18593;
    wire N__18592;
    wire N__18591;
    wire N__18590;
    wire N__18583;
    wire N__18580;
    wire N__18579;
    wire N__18578;
    wire N__18577;
    wire N__18576;
    wire N__18575;
    wire N__18570;
    wire N__18567;
    wire N__18558;
    wire N__18551;
    wire N__18548;
    wire N__18547;
    wire N__18546;
    wire N__18543;
    wire N__18540;
    wire N__18537;
    wire N__18534;
    wire N__18531;
    wire N__18528;
    wire N__18527;
    wire N__18520;
    wire N__18517;
    wire N__18514;
    wire N__18511;
    wire N__18506;
    wire N__18505;
    wire N__18502;
    wire N__18501;
    wire N__18498;
    wire N__18495;
    wire N__18492;
    wire N__18485;
    wire N__18484;
    wire N__18483;
    wire N__18480;
    wire N__18477;
    wire N__18474;
    wire N__18467;
    wire N__18464;
    wire N__18463;
    wire N__18462;
    wire N__18459;
    wire N__18454;
    wire N__18449;
    wire N__18446;
    wire N__18443;
    wire N__18442;
    wire N__18441;
    wire N__18438;
    wire N__18435;
    wire N__18432;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18416;
    wire N__18415;
    wire N__18412;
    wire N__18409;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18397;
    wire N__18396;
    wire N__18393;
    wire N__18390;
    wire N__18387;
    wire N__18382;
    wire N__18377;
    wire N__18374;
    wire N__18373;
    wire N__18370;
    wire N__18367;
    wire N__18362;
    wire N__18359;
    wire N__18356;
    wire N__18355;
    wire N__18354;
    wire N__18351;
    wire N__18348;
    wire N__18345;
    wire N__18340;
    wire N__18335;
    wire N__18332;
    wire N__18331;
    wire N__18330;
    wire N__18327;
    wire N__18326;
    wire N__18321;
    wire N__18318;
    wire N__18315;
    wire N__18312;
    wire N__18307;
    wire N__18304;
    wire N__18299;
    wire N__18296;
    wire N__18295;
    wire N__18294;
    wire N__18291;
    wire N__18286;
    wire N__18281;
    wire N__18278;
    wire N__18277;
    wire N__18274;
    wire N__18271;
    wire N__18268;
    wire N__18265;
    wire N__18262;
    wire N__18259;
    wire N__18254;
    wire N__18251;
    wire N__18250;
    wire N__18249;
    wire N__18246;
    wire N__18241;
    wire N__18236;
    wire N__18235;
    wire N__18232;
    wire N__18229;
    wire N__18226;
    wire N__18223;
    wire N__18220;
    wire N__18217;
    wire N__18214;
    wire N__18211;
    wire N__18206;
    wire N__18203;
    wire N__18200;
    wire N__18197;
    wire N__18196;
    wire N__18195;
    wire N__18194;
    wire N__18193;
    wire N__18192;
    wire N__18179;
    wire N__18176;
    wire N__18173;
    wire N__18170;
    wire N__18167;
    wire N__18164;
    wire N__18161;
    wire N__18158;
    wire N__18155;
    wire N__18152;
    wire N__18151;
    wire N__18150;
    wire N__18149;
    wire N__18148;
    wire N__18147;
    wire N__18136;
    wire N__18133;
    wire N__18128;
    wire N__18127;
    wire N__18126;
    wire N__18123;
    wire N__18122;
    wire N__18115;
    wire N__18112;
    wire N__18107;
    wire N__18106;
    wire N__18105;
    wire N__18102;
    wire N__18099;
    wire N__18096;
    wire N__18093;
    wire N__18090;
    wire N__18089;
    wire N__18086;
    wire N__18081;
    wire N__18078;
    wire N__18077;
    wire N__18074;
    wire N__18069;
    wire N__18066;
    wire N__18059;
    wire N__18058;
    wire N__18057;
    wire N__18056;
    wire N__18053;
    wire N__18050;
    wire N__18047;
    wire N__18044;
    wire N__18043;
    wire N__18040;
    wire N__18035;
    wire N__18030;
    wire N__18023;
    wire N__18022;
    wire N__18019;
    wire N__18018;
    wire N__18015;
    wire N__18012;
    wire N__18009;
    wire N__18006;
    wire N__18005;
    wire N__18002;
    wire N__17999;
    wire N__17996;
    wire N__17993;
    wire N__17984;
    wire N__17981;
    wire N__17978;
    wire N__17977;
    wire N__17974;
    wire N__17971;
    wire N__17970;
    wire N__17967;
    wire N__17964;
    wire N__17961;
    wire N__17960;
    wire N__17957;
    wire N__17952;
    wire N__17949;
    wire N__17942;
    wire N__17941;
    wire N__17940;
    wire N__17939;
    wire N__17938;
    wire N__17937;
    wire N__17932;
    wire N__17927;
    wire N__17922;
    wire N__17921;
    wire N__17920;
    wire N__17913;
    wire N__17908;
    wire N__17903;
    wire N__17902;
    wire N__17901;
    wire N__17900;
    wire N__17899;
    wire N__17896;
    wire N__17893;
    wire N__17882;
    wire N__17879;
    wire N__17878;
    wire N__17875;
    wire N__17872;
    wire N__17871;
    wire N__17866;
    wire N__17863;
    wire N__17858;
    wire N__17855;
    wire N__17852;
    wire N__17851;
    wire N__17850;
    wire N__17849;
    wire N__17846;
    wire N__17843;
    wire N__17840;
    wire N__17837;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17825;
    wire N__17820;
    wire N__17817;
    wire N__17810;
    wire N__17809;
    wire N__17804;
    wire N__17801;
    wire N__17798;
    wire N__17795;
    wire N__17792;
    wire N__17789;
    wire N__17788;
    wire N__17787;
    wire N__17784;
    wire N__17779;
    wire N__17774;
    wire N__17773;
    wire N__17770;
    wire N__17769;
    wire N__17766;
    wire N__17763;
    wire N__17760;
    wire N__17757;
    wire N__17750;
    wire N__17747;
    wire N__17746;
    wire N__17745;
    wire N__17742;
    wire N__17739;
    wire N__17736;
    wire N__17729;
    wire N__17726;
    wire N__17723;
    wire N__17720;
    wire N__17717;
    wire N__17716;
    wire N__17713;
    wire N__17710;
    wire N__17707;
    wire N__17704;
    wire N__17701;
    wire N__17696;
    wire N__17695;
    wire N__17692;
    wire N__17689;
    wire N__17686;
    wire N__17683;
    wire N__17680;
    wire N__17675;
    wire N__17674;
    wire N__17671;
    wire N__17668;
    wire N__17665;
    wire N__17662;
    wire N__17657;
    wire N__17654;
    wire N__17653;
    wire N__17650;
    wire N__17647;
    wire N__17644;
    wire N__17641;
    wire N__17636;
    wire N__17633;
    wire N__17630;
    wire N__17627;
    wire N__17624;
    wire N__17621;
    wire N__17618;
    wire N__17615;
    wire N__17612;
    wire N__17609;
    wire N__17606;
    wire N__17603;
    wire N__17600;
    wire N__17597;
    wire N__17594;
    wire N__17591;
    wire N__17588;
    wire N__17585;
    wire N__17582;
    wire N__17579;
    wire N__17576;
    wire N__17573;
    wire N__17570;
    wire N__17567;
    wire N__17566;
    wire N__17565;
    wire N__17564;
    wire N__17563;
    wire N__17562;
    wire N__17561;
    wire N__17560;
    wire N__17559;
    wire N__17558;
    wire N__17557;
    wire N__17556;
    wire N__17555;
    wire N__17554;
    wire N__17553;
    wire N__17552;
    wire N__17551;
    wire N__17550;
    wire N__17549;
    wire N__17548;
    wire N__17547;
    wire N__17546;
    wire N__17545;
    wire N__17544;
    wire N__17543;
    wire N__17542;
    wire N__17533;
    wire N__17532;
    wire N__17531;
    wire N__17530;
    wire N__17529;
    wire N__17524;
    wire N__17515;
    wire N__17506;
    wire N__17497;
    wire N__17488;
    wire N__17479;
    wire N__17476;
    wire N__17467;
    wire N__17464;
    wire N__17459;
    wire N__17452;
    wire N__17441;
    wire N__17438;
    wire N__17435;
    wire N__17432;
    wire N__17429;
    wire N__17428;
    wire N__17425;
    wire N__17422;
    wire N__17417;
    wire N__17414;
    wire N__17413;
    wire N__17410;
    wire N__17407;
    wire N__17402;
    wire N__17399;
    wire N__17396;
    wire N__17395;
    wire N__17392;
    wire N__17389;
    wire N__17388;
    wire N__17383;
    wire N__17380;
    wire N__17375;
    wire N__17372;
    wire N__17371;
    wire N__17368;
    wire N__17365;
    wire N__17362;
    wire N__17359;
    wire N__17356;
    wire N__17353;
    wire N__17348;
    wire N__17345;
    wire N__17344;
    wire N__17341;
    wire N__17338;
    wire N__17337;
    wire N__17332;
    wire N__17329;
    wire N__17324;
    wire N__17321;
    wire N__17318;
    wire N__17315;
    wire N__17312;
    wire N__17309;
    wire N__17306;
    wire N__17303;
    wire N__17300;
    wire N__17297;
    wire N__17294;
    wire N__17291;
    wire N__17288;
    wire N__17285;
    wire N__17282;
    wire N__17279;
    wire N__17276;
    wire N__17273;
    wire N__17270;
    wire N__17267;
    wire N__17266;
    wire N__17265;
    wire N__17264;
    wire N__17261;
    wire N__17258;
    wire N__17255;
    wire N__17252;
    wire N__17243;
    wire N__17240;
    wire N__17237;
    wire N__17234;
    wire N__17233;
    wire N__17232;
    wire N__17229;
    wire N__17226;
    wire N__17223;
    wire N__17216;
    wire N__17213;
    wire N__17212;
    wire N__17211;
    wire N__17208;
    wire N__17205;
    wire N__17202;
    wire N__17195;
    wire N__17194;
    wire N__17193;
    wire N__17192;
    wire N__17191;
    wire N__17180;
    wire N__17177;
    wire N__17174;
    wire N__17171;
    wire N__17168;
    wire N__17165;
    wire N__17162;
    wire N__17159;
    wire N__17156;
    wire N__17153;
    wire N__17150;
    wire N__17147;
    wire N__17144;
    wire N__17141;
    wire N__17138;
    wire N__17135;
    wire N__17132;
    wire N__17129;
    wire N__17126;
    wire N__17123;
    wire N__17120;
    wire N__17117;
    wire N__17114;
    wire N__17111;
    wire N__17110;
    wire N__17107;
    wire N__17104;
    wire N__17099;
    wire N__17096;
    wire N__17093;
    wire N__17092;
    wire N__17089;
    wire N__17086;
    wire N__17085;
    wire N__17082;
    wire N__17079;
    wire N__17076;
    wire N__17069;
    wire N__17068;
    wire N__17065;
    wire N__17062;
    wire N__17061;
    wire N__17058;
    wire N__17055;
    wire N__17052;
    wire N__17049;
    wire N__17044;
    wire N__17039;
    wire N__17038;
    wire N__17035;
    wire N__17032;
    wire N__17031;
    wire N__17026;
    wire N__17023;
    wire N__17022;
    wire N__17017;
    wire N__17016;
    wire N__17013;
    wire N__17010;
    wire N__17007;
    wire N__17000;
    wire N__16999;
    wire N__16998;
    wire N__16997;
    wire N__16996;
    wire N__16995;
    wire N__16994;
    wire N__16987;
    wire N__16984;
    wire N__16979;
    wire N__16976;
    wire N__16973;
    wire N__16966;
    wire N__16965;
    wire N__16964;
    wire N__16963;
    wire N__16960;
    wire N__16957;
    wire N__16952;
    wire N__16949;
    wire N__16942;
    wire N__16939;
    wire N__16934;
    wire N__16931;
    wire N__16928;
    wire N__16927;
    wire N__16924;
    wire N__16921;
    wire N__16920;
    wire N__16915;
    wire N__16912;
    wire N__16907;
    wire N__16904;
    wire N__16901;
    wire N__16898;
    wire N__16895;
    wire N__16892;
    wire N__16891;
    wire N__16890;
    wire N__16889;
    wire N__16886;
    wire N__16883;
    wire N__16880;
    wire N__16877;
    wire N__16874;
    wire N__16869;
    wire N__16866;
    wire N__16859;
    wire N__16856;
    wire N__16853;
    wire N__16850;
    wire N__16847;
    wire N__16844;
    wire N__16841;
    wire N__16838;
    wire N__16835;
    wire N__16832;
    wire N__16829;
    wire N__16826;
    wire N__16823;
    wire N__16820;
    wire N__16819;
    wire N__16816;
    wire N__16813;
    wire N__16808;
    wire N__16807;
    wire N__16804;
    wire N__16801;
    wire N__16796;
    wire N__16793;
    wire N__16792;
    wire N__16789;
    wire N__16786;
    wire N__16783;
    wire N__16782;
    wire N__16779;
    wire N__16778;
    wire N__16775;
    wire N__16772;
    wire N__16769;
    wire N__16766;
    wire N__16761;
    wire N__16754;
    wire N__16751;
    wire N__16750;
    wire N__16747;
    wire N__16744;
    wire N__16741;
    wire N__16738;
    wire N__16737;
    wire N__16736;
    wire N__16733;
    wire N__16730;
    wire N__16727;
    wire N__16724;
    wire N__16715;
    wire N__16712;
    wire N__16711;
    wire N__16708;
    wire N__16705;
    wire N__16702;
    wire N__16699;
    wire N__16698;
    wire N__16697;
    wire N__16694;
    wire N__16691;
    wire N__16688;
    wire N__16685;
    wire N__16676;
    wire N__16673;
    wire N__16672;
    wire N__16669;
    wire N__16666;
    wire N__16665;
    wire N__16660;
    wire N__16657;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16645;
    wire N__16642;
    wire N__16639;
    wire N__16638;
    wire N__16635;
    wire N__16632;
    wire N__16629;
    wire N__16622;
    wire N__16619;
    wire N__16618;
    wire N__16615;
    wire N__16612;
    wire N__16611;
    wire N__16606;
    wire N__16603;
    wire N__16600;
    wire N__16597;
    wire N__16592;
    wire N__16589;
    wire N__16588;
    wire N__16585;
    wire N__16582;
    wire N__16577;
    wire N__16576;
    wire N__16573;
    wire N__16570;
    wire N__16565;
    wire N__16564;
    wire N__16561;
    wire N__16558;
    wire N__16555;
    wire N__16552;
    wire N__16549;
    wire N__16548;
    wire N__16543;
    wire N__16540;
    wire N__16535;
    wire N__16532;
    wire N__16531;
    wire N__16528;
    wire N__16525;
    wire N__16522;
    wire N__16519;
    wire N__16516;
    wire N__16515;
    wire N__16510;
    wire N__16507;
    wire N__16504;
    wire N__16501;
    wire N__16496;
    wire N__16493;
    wire N__16490;
    wire N__16487;
    wire N__16484;
    wire N__16483;
    wire N__16480;
    wire N__16477;
    wire N__16474;
    wire N__16471;
    wire N__16466;
    wire N__16463;
    wire N__16460;
    wire N__16457;
    wire N__16456;
    wire N__16453;
    wire N__16450;
    wire N__16449;
    wire N__16446;
    wire N__16443;
    wire N__16440;
    wire N__16437;
    wire N__16432;
    wire N__16429;
    wire N__16426;
    wire N__16421;
    wire N__16420;
    wire N__16417;
    wire N__16414;
    wire N__16411;
    wire N__16408;
    wire N__16405;
    wire N__16402;
    wire N__16401;
    wire N__16398;
    wire N__16395;
    wire N__16392;
    wire N__16389;
    wire N__16386;
    wire N__16383;
    wire N__16376;
    wire N__16375;
    wire N__16374;
    wire N__16371;
    wire N__16368;
    wire N__16365;
    wire N__16360;
    wire N__16355;
    wire N__16352;
    wire N__16351;
    wire N__16350;
    wire N__16347;
    wire N__16344;
    wire N__16341;
    wire N__16336;
    wire N__16331;
    wire N__16328;
    wire N__16327;
    wire N__16326;
    wire N__16323;
    wire N__16320;
    wire N__16317;
    wire N__16310;
    wire N__16307;
    wire N__16306;
    wire N__16305;
    wire N__16302;
    wire N__16299;
    wire N__16296;
    wire N__16289;
    wire N__16286;
    wire N__16285;
    wire N__16282;
    wire N__16279;
    wire N__16274;
    wire N__16273;
    wire N__16272;
    wire N__16269;
    wire N__16266;
    wire N__16263;
    wire N__16258;
    wire N__16253;
    wire N__16250;
    wire N__16249;
    wire N__16246;
    wire N__16243;
    wire N__16238;
    wire N__16237;
    wire N__16236;
    wire N__16233;
    wire N__16230;
    wire N__16227;
    wire N__16222;
    wire N__16217;
    wire N__16214;
    wire N__16211;
    wire N__16210;
    wire N__16209;
    wire N__16206;
    wire N__16203;
    wire N__16200;
    wire N__16195;
    wire N__16190;
    wire N__16187;
    wire N__16186;
    wire N__16185;
    wire N__16182;
    wire N__16179;
    wire N__16176;
    wire N__16171;
    wire N__16166;
    wire N__16163;
    wire N__16162;
    wire N__16161;
    wire N__16158;
    wire N__16155;
    wire N__16152;
    wire N__16145;
    wire N__16142;
    wire N__16141;
    wire N__16140;
    wire N__16137;
    wire N__16134;
    wire N__16131;
    wire N__16124;
    wire N__16121;
    wire N__16120;
    wire N__16119;
    wire N__16116;
    wire N__16113;
    wire N__16110;
    wire N__16105;
    wire N__16100;
    wire N__16097;
    wire N__16096;
    wire N__16095;
    wire N__16092;
    wire N__16089;
    wire N__16086;
    wire N__16081;
    wire N__16076;
    wire N__16073;
    wire N__16072;
    wire N__16071;
    wire N__16068;
    wire N__16063;
    wire N__16058;
    wire N__16055;
    wire N__16054;
    wire N__16053;
    wire N__16050;
    wire N__16045;
    wire N__16040;
    wire N__16037;
    wire N__16036;
    wire N__16035;
    wire N__16032;
    wire N__16027;
    wire N__16022;
    wire N__16019;
    wire N__16018;
    wire N__16017;
    wire N__16014;
    wire N__16011;
    wire N__16008;
    wire N__16003;
    wire N__15998;
    wire N__15995;
    wire N__15994;
    wire N__15993;
    wire N__15990;
    wire N__15987;
    wire N__15984;
    wire N__15979;
    wire N__15974;
    wire N__15971;
    wire N__15970;
    wire N__15969;
    wire N__15966;
    wire N__15963;
    wire N__15960;
    wire N__15953;
    wire N__15950;
    wire N__15949;
    wire N__15948;
    wire N__15945;
    wire N__15942;
    wire N__15939;
    wire N__15932;
    wire N__15929;
    wire N__15928;
    wire N__15927;
    wire N__15924;
    wire N__15921;
    wire N__15918;
    wire N__15913;
    wire N__15908;
    wire N__15905;
    wire N__15904;
    wire N__15903;
    wire N__15900;
    wire N__15897;
    wire N__15894;
    wire N__15889;
    wire N__15884;
    wire N__15881;
    wire N__15880;
    wire N__15879;
    wire N__15876;
    wire N__15871;
    wire N__15866;
    wire N__15863;
    wire N__15862;
    wire N__15861;
    wire N__15858;
    wire N__15853;
    wire N__15848;
    wire N__15845;
    wire N__15844;
    wire N__15843;
    wire N__15836;
    wire N__15833;
    wire N__15832;
    wire N__15831;
    wire N__15830;
    wire N__15829;
    wire N__15828;
    wire N__15827;
    wire N__15816;
    wire N__15813;
    wire N__15810;
    wire N__15803;
    wire N__15802;
    wire N__15801;
    wire N__15800;
    wire N__15799;
    wire N__15798;
    wire N__15791;
    wire N__15786;
    wire N__15783;
    wire N__15776;
    wire N__15773;
    wire N__15772;
    wire N__15771;
    wire N__15768;
    wire N__15765;
    wire N__15762;
    wire N__15759;
    wire N__15756;
    wire N__15753;
    wire N__15746;
    wire N__15743;
    wire N__15740;
    wire N__15739;
    wire N__15736;
    wire N__15733;
    wire N__15732;
    wire N__15729;
    wire N__15726;
    wire N__15723;
    wire N__15720;
    wire N__15717;
    wire N__15714;
    wire N__15707;
    wire N__15706;
    wire N__15703;
    wire N__15700;
    wire N__15699;
    wire N__15696;
    wire N__15695;
    wire N__15692;
    wire N__15689;
    wire N__15686;
    wire N__15683;
    wire N__15678;
    wire N__15671;
    wire N__15668;
    wire N__15665;
    wire N__15662;
    wire N__15659;
    wire N__15658;
    wire N__15657;
    wire N__15654;
    wire N__15651;
    wire N__15648;
    wire N__15643;
    wire N__15638;
    wire N__15635;
    wire N__15634;
    wire N__15633;
    wire N__15630;
    wire N__15627;
    wire N__15624;
    wire N__15619;
    wire N__15614;
    wire N__15611;
    wire N__15610;
    wire N__15609;
    wire N__15606;
    wire N__15601;
    wire N__15596;
    wire N__15593;
    wire N__15590;
    wire N__15589;
    wire N__15584;
    wire N__15581;
    wire N__15578;
    wire N__15575;
    wire N__15572;
    wire N__15569;
    wire N__15566;
    wire N__15563;
    wire N__15560;
    wire N__15559;
    wire N__15554;
    wire N__15551;
    wire N__15548;
    wire N__15545;
    wire N__15542;
    wire N__15539;
    wire N__15538;
    wire N__15537;
    wire N__15534;
    wire N__15533;
    wire N__15532;
    wire N__15531;
    wire N__15530;
    wire N__15529;
    wire N__15524;
    wire N__15517;
    wire N__15512;
    wire N__15509;
    wire N__15500;
    wire N__15499;
    wire N__15498;
    wire N__15495;
    wire N__15492;
    wire N__15489;
    wire N__15482;
    wire N__15479;
    wire N__15478;
    wire N__15475;
    wire N__15472;
    wire N__15471;
    wire N__15470;
    wire N__15469;
    wire N__15468;
    wire N__15467;
    wire N__15466;
    wire N__15463;
    wire N__15460;
    wire N__15459;
    wire N__15458;
    wire N__15457;
    wire N__15456;
    wire N__15455;
    wire N__15454;
    wire N__15453;
    wire N__15452;
    wire N__15451;
    wire N__15440;
    wire N__15437;
    wire N__15436;
    wire N__15435;
    wire N__15434;
    wire N__15433;
    wire N__15432;
    wire N__15429;
    wire N__15426;
    wire N__15421;
    wire N__15420;
    wire N__15405;
    wire N__15402;
    wire N__15399;
    wire N__15398;
    wire N__15395;
    wire N__15392;
    wire N__15385;
    wire N__15382;
    wire N__15377;
    wire N__15374;
    wire N__15367;
    wire N__15364;
    wire N__15347;
    wire N__15346;
    wire N__15345;
    wire N__15344;
    wire N__15343;
    wire N__15342;
    wire N__15341;
    wire N__15338;
    wire N__15337;
    wire N__15336;
    wire N__15335;
    wire N__15334;
    wire N__15331;
    wire N__15330;
    wire N__15327;
    wire N__15324;
    wire N__15321;
    wire N__15320;
    wire N__15319;
    wire N__15318;
    wire N__15317;
    wire N__15316;
    wire N__15313;
    wire N__15310;
    wire N__15307;
    wire N__15306;
    wire N__15305;
    wire N__15304;
    wire N__15303;
    wire N__15300;
    wire N__15297;
    wire N__15294;
    wire N__15291;
    wire N__15286;
    wire N__15285;
    wire N__15282;
    wire N__15275;
    wire N__15262;
    wire N__15259;
    wire N__15242;
    wire N__15239;
    wire N__15236;
    wire N__15235;
    wire N__15230;
    wire N__15227;
    wire N__15222;
    wire N__15221;
    wire N__15218;
    wire N__15215;
    wire N__15212;
    wire N__15209;
    wire N__15204;
    wire N__15201;
    wire N__15196;
    wire N__15185;
    wire N__15184;
    wire N__15181;
    wire N__15178;
    wire N__15177;
    wire N__15172;
    wire N__15169;
    wire N__15168;
    wire N__15167;
    wire N__15164;
    wire N__15161;
    wire N__15156;
    wire N__15149;
    wire N__15148;
    wire N__15147;
    wire N__15146;
    wire N__15145;
    wire N__15144;
    wire N__15143;
    wire N__15142;
    wire N__15141;
    wire N__15140;
    wire N__15137;
    wire N__15136;
    wire N__15135;
    wire N__15134;
    wire N__15133;
    wire N__15132;
    wire N__15131;
    wire N__15130;
    wire N__15129;
    wire N__15124;
    wire N__15111;
    wire N__15108;
    wire N__15107;
    wire N__15106;
    wire N__15105;
    wire N__15104;
    wire N__15103;
    wire N__15100;
    wire N__15083;
    wire N__15078;
    wire N__15075;
    wire N__15074;
    wire N__15071;
    wire N__15068;
    wire N__15063;
    wire N__15060;
    wire N__15051;
    wire N__15048;
    wire N__15035;
    wire N__15034;
    wire N__15031;
    wire N__15028;
    wire N__15025;
    wire N__15022;
    wire N__15017;
    wire N__15014;
    wire N__15011;
    wire N__15008;
    wire N__15005;
    wire N__15002;
    wire N__15001;
    wire N__15000;
    wire N__14997;
    wire N__14992;
    wire N__14987;
    wire N__14984;
    wire N__14983;
    wire N__14980;
    wire N__14977;
    wire N__14974;
    wire N__14969;
    wire N__14966;
    wire N__14963;
    wire N__14960;
    wire N__14959;
    wire N__14956;
    wire N__14953;
    wire N__14950;
    wire N__14945;
    wire N__14942;
    wire N__14939;
    wire N__14936;
    wire N__14935;
    wire N__14932;
    wire N__14929;
    wire N__14926;
    wire N__14921;
    wire N__14918;
    wire N__14915;
    wire N__14912;
    wire N__14911;
    wire N__14908;
    wire N__14905;
    wire N__14902;
    wire N__14897;
    wire N__14894;
    wire N__14891;
    wire N__14888;
    wire N__14887;
    wire N__14884;
    wire N__14881;
    wire N__14880;
    wire N__14879;
    wire N__14876;
    wire N__14873;
    wire N__14868;
    wire N__14865;
    wire N__14862;
    wire N__14859;
    wire N__14852;
    wire N__14849;
    wire N__14848;
    wire N__14847;
    wire N__14846;
    wire N__14843;
    wire N__14836;
    wire N__14831;
    wire N__14828;
    wire N__14827;
    wire N__14826;
    wire N__14825;
    wire N__14824;
    wire N__14823;
    wire N__14816;
    wire N__14815;
    wire N__14814;
    wire N__14807;
    wire N__14804;
    wire N__14801;
    wire N__14800;
    wire N__14799;
    wire N__14798;
    wire N__14795;
    wire N__14794;
    wire N__14791;
    wire N__14788;
    wire N__14775;
    wire N__14772;
    wire N__14769;
    wire N__14766;
    wire N__14759;
    wire N__14758;
    wire N__14757;
    wire N__14756;
    wire N__14751;
    wire N__14746;
    wire N__14745;
    wire N__14742;
    wire N__14739;
    wire N__14736;
    wire N__14729;
    wire N__14726;
    wire N__14723;
    wire N__14722;
    wire N__14721;
    wire N__14720;
    wire N__14719;
    wire N__14718;
    wire N__14717;
    wire N__14716;
    wire N__14709;
    wire N__14698;
    wire N__14697;
    wire N__14696;
    wire N__14695;
    wire N__14694;
    wire N__14693;
    wire N__14692;
    wire N__14691;
    wire N__14690;
    wire N__14687;
    wire N__14684;
    wire N__14667;
    wire N__14664;
    wire N__14661;
    wire N__14658;
    wire N__14651;
    wire N__14650;
    wire N__14647;
    wire N__14644;
    wire N__14641;
    wire N__14636;
    wire N__14633;
    wire N__14630;
    wire N__14627;
    wire N__14624;
    wire N__14621;
    wire N__14620;
    wire N__14617;
    wire N__14614;
    wire N__14611;
    wire N__14606;
    wire N__14603;
    wire N__14600;
    wire N__14597;
    wire N__14596;
    wire N__14593;
    wire N__14590;
    wire N__14587;
    wire N__14582;
    wire N__14579;
    wire N__14576;
    wire N__14573;
    wire N__14570;
    wire N__14569;
    wire N__14566;
    wire N__14563;
    wire N__14560;
    wire N__14555;
    wire N__14552;
    wire N__14549;
    wire N__14546;
    wire N__14543;
    wire N__14542;
    wire N__14539;
    wire N__14536;
    wire N__14533;
    wire N__14528;
    wire N__14525;
    wire N__14522;
    wire N__14519;
    wire N__14516;
    wire N__14515;
    wire N__14512;
    wire N__14509;
    wire N__14506;
    wire N__14501;
    wire N__14498;
    wire N__14495;
    wire N__14492;
    wire N__14491;
    wire N__14488;
    wire N__14485;
    wire N__14482;
    wire N__14477;
    wire N__14474;
    wire N__14471;
    wire N__14468;
    wire N__14465;
    wire N__14464;
    wire N__14461;
    wire N__14458;
    wire N__14455;
    wire N__14450;
    wire N__14447;
    wire N__14444;
    wire N__14441;
    wire N__14440;
    wire N__14437;
    wire N__14434;
    wire N__14433;
    wire N__14430;
    wire N__14427;
    wire N__14424;
    wire N__14417;
    wire N__14414;
    wire N__14411;
    wire N__14408;
    wire N__14405;
    wire N__14402;
    wire N__14399;
    wire N__14398;
    wire N__14395;
    wire N__14392;
    wire N__14387;
    wire N__14384;
    wire N__14381;
    wire N__14378;
    wire N__14375;
    wire N__14372;
    wire N__14369;
    wire N__14368;
    wire N__14365;
    wire N__14362;
    wire N__14357;
    wire N__14354;
    wire N__14351;
    wire N__14348;
    wire N__14345;
    wire N__14342;
    wire N__14339;
    wire N__14336;
    wire N__14333;
    wire N__14330;
    wire N__14327;
    wire N__14324;
    wire N__14321;
    wire N__14320;
    wire N__14317;
    wire N__14314;
    wire N__14309;
    wire N__14306;
    wire N__14303;
    wire N__14300;
    wire N__14297;
    wire N__14294;
    wire N__14291;
    wire N__14288;
    wire N__14287;
    wire N__14284;
    wire N__14281;
    wire N__14276;
    wire N__14273;
    wire N__14270;
    wire N__14267;
    wire N__14264;
    wire N__14261;
    wire N__14258;
    wire N__14255;
    wire N__14254;
    wire N__14251;
    wire N__14248;
    wire N__14243;
    wire N__14240;
    wire N__14237;
    wire N__14234;
    wire N__14231;
    wire N__14228;
    wire N__14225;
    wire N__14224;
    wire N__14221;
    wire N__14218;
    wire N__14215;
    wire N__14210;
    wire N__14207;
    wire N__14204;
    wire N__14201;
    wire N__14198;
    wire N__14195;
    wire N__14192;
    wire N__14189;
    wire N__14186;
    wire N__14183;
    wire N__14180;
    wire N__14177;
    wire N__14174;
    wire N__14173;
    wire N__14172;
    wire N__14171;
    wire N__14162;
    wire N__14159;
    wire N__14156;
    wire N__14153;
    wire N__14150;
    wire N__14147;
    wire N__14144;
    wire N__14141;
    wire N__14138;
    wire N__14135;
    wire N__14132;
    wire N__14129;
    wire N__14126;
    wire N__14123;
    wire N__14120;
    wire N__14117;
    wire N__14114;
    wire N__14111;
    wire N__14108;
    wire N__14105;
    wire N__14102;
    wire N__14099;
    wire N__14096;
    wire N__14095;
    wire N__14092;
    wire N__14089;
    wire N__14088;
    wire N__14085;
    wire N__14082;
    wire N__14079;
    wire N__14076;
    wire N__14071;
    wire N__14066;
    wire N__14063;
    wire N__14062;
    wire N__14061;
    wire N__14058;
    wire N__14055;
    wire N__14054;
    wire N__14051;
    wire N__14048;
    wire N__14045;
    wire N__14042;
    wire N__14039;
    wire N__14032;
    wire N__14029;
    wire N__14024;
    wire N__14021;
    wire N__14020;
    wire N__14019;
    wire N__14016;
    wire N__14015;
    wire N__14012;
    wire N__14009;
    wire N__14006;
    wire N__14003;
    wire N__14000;
    wire N__13997;
    wire N__13994;
    wire N__13991;
    wire N__13986;
    wire N__13979;
    wire N__13976;
    wire N__13975;
    wire N__13974;
    wire N__13973;
    wire N__13970;
    wire N__13967;
    wire N__13966;
    wire N__13961;
    wire N__13958;
    wire N__13955;
    wire N__13952;
    wire N__13949;
    wire N__13942;
    wire N__13939;
    wire N__13934;
    wire N__13933;
    wire N__13930;
    wire N__13927;
    wire N__13926;
    wire N__13923;
    wire N__13922;
    wire N__13919;
    wire N__13916;
    wire N__13913;
    wire N__13910;
    wire N__13907;
    wire N__13904;
    wire N__13901;
    wire N__13898;
    wire N__13893;
    wire N__13888;
    wire N__13883;
    wire N__13882;
    wire N__13881;
    wire N__13878;
    wire N__13875;
    wire N__13872;
    wire N__13871;
    wire N__13868;
    wire N__13863;
    wire N__13860;
    wire N__13857;
    wire N__13854;
    wire N__13847;
    wire N__13846;
    wire N__13843;
    wire N__13842;
    wire N__13839;
    wire N__13838;
    wire N__13835;
    wire N__13832;
    wire N__13829;
    wire N__13826;
    wire N__13823;
    wire N__13820;
    wire N__13817;
    wire N__13808;
    wire N__13805;
    wire N__13802;
    wire N__13799;
    wire N__13798;
    wire N__13795;
    wire N__13792;
    wire N__13791;
    wire N__13788;
    wire N__13785;
    wire N__13782;
    wire N__13775;
    wire N__13772;
    wire N__13769;
    wire N__13768;
    wire N__13765;
    wire N__13762;
    wire N__13761;
    wire N__13758;
    wire N__13755;
    wire N__13752;
    wire N__13745;
    wire N__13742;
    wire N__13741;
    wire N__13738;
    wire N__13735;
    wire N__13732;
    wire N__13729;
    wire N__13726;
    wire N__13725;
    wire N__13722;
    wire N__13719;
    wire N__13716;
    wire N__13713;
    wire N__13708;
    wire N__13703;
    wire N__13700;
    wire N__13699;
    wire N__13696;
    wire N__13693;
    wire N__13692;
    wire N__13689;
    wire N__13686;
    wire N__13683;
    wire N__13676;
    wire N__13673;
    wire N__13672;
    wire N__13671;
    wire N__13670;
    wire N__13669;
    wire N__13666;
    wire N__13655;
    wire N__13652;
    wire N__13649;
    wire N__13648;
    wire N__13645;
    wire N__13642;
    wire N__13639;
    wire N__13636;
    wire N__13633;
    wire N__13630;
    wire N__13627;
    wire N__13624;
    wire N__13619;
    wire N__13618;
    wire N__13615;
    wire N__13612;
    wire N__13611;
    wire N__13608;
    wire N__13605;
    wire N__13602;
    wire N__13599;
    wire N__13594;
    wire N__13589;
    wire N__13586;
    wire N__13585;
    wire N__13584;
    wire N__13581;
    wire N__13578;
    wire N__13575;
    wire N__13572;
    wire N__13569;
    wire N__13566;
    wire N__13559;
    wire N__13556;
    wire N__13555;
    wire N__13554;
    wire N__13553;
    wire N__13552;
    wire N__13551;
    wire N__13550;
    wire N__13543;
    wire N__13542;
    wire N__13541;
    wire N__13540;
    wire N__13537;
    wire N__13530;
    wire N__13527;
    wire N__13522;
    wire N__13517;
    wire N__13514;
    wire N__13507;
    wire N__13502;
    wire N__13499;
    wire N__13498;
    wire N__13495;
    wire N__13492;
    wire N__13491;
    wire N__13490;
    wire N__13487;
    wire N__13484;
    wire N__13481;
    wire N__13478;
    wire N__13475;
    wire N__13472;
    wire N__13469;
    wire N__13466;
    wire N__13463;
    wire N__13458;
    wire N__13455;
    wire N__13452;
    wire N__13445;
    wire N__13442;
    wire N__13439;
    wire N__13436;
    wire N__13433;
    wire N__13430;
    wire N__13427;
    wire N__13424;
    wire N__13421;
    wire N__13418;
    wire N__13417;
    wire N__13416;
    wire N__13413;
    wire N__13410;
    wire N__13407;
    wire N__13404;
    wire N__13401;
    wire N__13398;
    wire N__13395;
    wire N__13392;
    wire N__13389;
    wire N__13382;
    wire N__13379;
    wire N__13378;
    wire N__13377;
    wire N__13374;
    wire N__13371;
    wire N__13368;
    wire N__13365;
    wire N__13362;
    wire N__13359;
    wire N__13356;
    wire N__13353;
    wire N__13350;
    wire N__13343;
    wire N__13340;
    wire N__13339;
    wire N__13336;
    wire N__13333;
    wire N__13332;
    wire N__13329;
    wire N__13326;
    wire N__13323;
    wire N__13320;
    wire N__13317;
    wire N__13314;
    wire N__13307;
    wire N__13306;
    wire N__13303;
    wire N__13302;
    wire N__13297;
    wire N__13294;
    wire N__13289;
    wire N__13288;
    wire N__13283;
    wire N__13282;
    wire N__13281;
    wire N__13278;
    wire N__13275;
    wire N__13272;
    wire N__13267;
    wire N__13262;
    wire N__13259;
    wire N__13256;
    wire N__13253;
    wire N__13250;
    wire N__13247;
    wire N__13244;
    wire N__13241;
    wire N__13238;
    wire N__13235;
    wire N__13232;
    wire N__13229;
    wire N__13226;
    wire N__13223;
    wire N__13220;
    wire N__13217;
    wire N__13216;
    wire N__13213;
    wire N__13210;
    wire N__13205;
    wire N__13204;
    wire N__13201;
    wire N__13198;
    wire N__13193;
    wire N__13190;
    wire N__13187;
    wire N__13184;
    wire N__13181;
    wire N__13178;
    wire N__13175;
    wire N__13172;
    wire N__13169;
    wire N__13166;
    wire N__13163;
    wire N__13160;
    wire N__13159;
    wire N__13154;
    wire N__13151;
    wire N__13150;
    wire N__13147;
    wire N__13144;
    wire N__13139;
    wire N__13138;
    wire N__13133;
    wire N__13130;
    wire N__13127;
    wire N__13126;
    wire N__13125;
    wire N__13122;
    wire N__13119;
    wire N__13116;
    wire N__13113;
    wire N__13106;
    wire N__13105;
    wire N__13102;
    wire N__13099;
    wire N__13094;
    wire N__13093;
    wire N__13088;
    wire N__13085;
    wire N__13084;
    wire N__13083;
    wire N__13078;
    wire N__13075;
    wire N__13072;
    wire N__13071;
    wire N__13068;
    wire N__13065;
    wire N__13062;
    wire N__13059;
    wire N__13058;
    wire N__13057;
    wire N__13052;
    wire N__13049;
    wire N__13046;
    wire N__13043;
    wire N__13040;
    wire N__13035;
    wire N__13032;
    wire N__13025;
    wire N__13022;
    wire N__13019;
    wire N__13016;
    wire N__13015;
    wire N__13014;
    wire N__13011;
    wire N__13008;
    wire N__13005;
    wire N__13002;
    wire N__12997;
    wire N__12992;
    wire N__12989;
    wire N__12986;
    wire N__12983;
    wire N__12980;
    wire N__12977;
    wire N__12974;
    wire N__12971;
    wire N__12968;
    wire N__12965;
    wire N__12962;
    wire N__12961;
    wire N__12960;
    wire N__12955;
    wire N__12952;
    wire N__12947;
    wire N__12944;
    wire N__12941;
    wire N__12940;
    wire N__12937;
    wire N__12936;
    wire N__12931;
    wire N__12928;
    wire N__12927;
    wire N__12924;
    wire N__12919;
    wire N__12914;
    wire N__12913;
    wire N__12912;
    wire N__12911;
    wire N__12910;
    wire N__12909;
    wire N__12908;
    wire N__12907;
    wire N__12906;
    wire N__12905;
    wire N__12904;
    wire N__12903;
    wire N__12902;
    wire N__12899;
    wire N__12896;
    wire N__12893;
    wire N__12892;
    wire N__12889;
    wire N__12888;
    wire N__12885;
    wire N__12882;
    wire N__12881;
    wire N__12880;
    wire N__12879;
    wire N__12878;
    wire N__12875;
    wire N__12872;
    wire N__12869;
    wire N__12866;
    wire N__12863;
    wire N__12862;
    wire N__12861;
    wire N__12858;
    wire N__12855;
    wire N__12854;
    wire N__12853;
    wire N__12844;
    wire N__12835;
    wire N__12818;
    wire N__12813;
    wire N__12810;
    wire N__12803;
    wire N__12800;
    wire N__12799;
    wire N__12794;
    wire N__12791;
    wire N__12786;
    wire N__12783;
    wire N__12780;
    wire N__12777;
    wire N__12774;
    wire N__12769;
    wire N__12764;
    wire N__12755;
    wire N__12752;
    wire N__12749;
    wire N__12746;
    wire N__12743;
    wire N__12740;
    wire N__12737;
    wire N__12736;
    wire N__12735;
    wire N__12728;
    wire N__12727;
    wire N__12726;
    wire N__12725;
    wire N__12724;
    wire N__12723;
    wire N__12722;
    wire N__12721;
    wire N__12718;
    wire N__12707;
    wire N__12702;
    wire N__12695;
    wire N__12692;
    wire N__12689;
    wire N__12686;
    wire N__12683;
    wire N__12680;
    wire N__12677;
    wire N__12674;
    wire N__12671;
    wire N__12668;
    wire N__12667;
    wire N__12666;
    wire N__12663;
    wire N__12660;
    wire N__12657;
    wire N__12652;
    wire N__12649;
    wire N__12646;
    wire N__12641;
    wire N__12638;
    wire N__12635;
    wire N__12632;
    wire N__12629;
    wire N__12626;
    wire N__12623;
    wire N__12620;
    wire N__12617;
    wire N__12614;
    wire N__12611;
    wire N__12608;
    wire N__12605;
    wire N__12602;
    wire N__12599;
    wire N__12596;
    wire N__12593;
    wire N__12590;
    wire N__12587;
    wire N__12584;
    wire N__12581;
    wire N__12578;
    wire N__12575;
    wire N__12572;
    wire N__12569;
    wire N__12566;
    wire N__12563;
    wire N__12560;
    wire N__12557;
    wire N__12554;
    wire N__12551;
    wire N__12548;
    wire N__12545;
    wire N__12542;
    wire N__12539;
    wire N__12536;
    wire N__12533;
    wire N__12530;
    wire N__12527;
    wire N__12524;
    wire N__12521;
    wire N__12518;
    wire N__12515;
    wire N__12512;
    wire N__12509;
    wire N__12506;
    wire N__12503;
    wire N__12500;
    wire N__12497;
    wire N__12494;
    wire N__12491;
    wire N__12488;
    wire N__12485;
    wire N__12482;
    wire N__12479;
    wire N__12476;
    wire N__12473;
    wire N__12470;
    wire N__12467;
    wire N__12464;
    wire N__12461;
    wire N__12458;
    wire N__12455;
    wire N__12452;
    wire N__12449;
    wire N__12446;
    wire N__12443;
    wire N__12440;
    wire N__12437;
    wire N__12434;
    wire N__12431;
    wire N__12428;
    wire N__12425;
    wire N__12422;
    wire N__12419;
    wire N__12416;
    wire N__12413;
    wire N__12410;
    wire N__12407;
    wire N__12404;
    wire N__12401;
    wire N__12398;
    wire N__12395;
    wire N__12392;
    wire N__12389;
    wire N__12386;
    wire N__12383;
    wire N__12380;
    wire N__12379;
    wire N__12378;
    wire N__12375;
    wire N__12372;
    wire N__12369;
    wire N__12364;
    wire N__12359;
    wire N__12358;
    wire N__12355;
    wire N__12352;
    wire N__12347;
    wire N__12346;
    wire N__12341;
    wire N__12340;
    wire N__12339;
    wire N__12336;
    wire N__12333;
    wire N__12330;
    wire N__12323;
    wire N__12322;
    wire N__12321;
    wire N__12318;
    wire N__12315;
    wire N__12314;
    wire N__12311;
    wire N__12308;
    wire N__12305;
    wire N__12302;
    wire N__12295;
    wire N__12290;
    wire N__12287;
    wire N__12286;
    wire N__12285;
    wire N__12284;
    wire N__12281;
    wire N__12278;
    wire N__12277;
    wire N__12272;
    wire N__12267;
    wire N__12264;
    wire N__12257;
    wire N__12256;
    wire N__12253;
    wire N__12250;
    wire N__12245;
    wire N__12244;
    wire N__12243;
    wire N__12242;
    wire N__12241;
    wire N__12238;
    wire N__12235;
    wire N__12232;
    wire N__12231;
    wire N__12230;
    wire N__12229;
    wire N__12228;
    wire N__12227;
    wire N__12226;
    wire N__12225;
    wire N__12224;
    wire N__12223;
    wire N__12222;
    wire N__12221;
    wire N__12220;
    wire N__12217;
    wire N__12214;
    wire N__12199;
    wire N__12196;
    wire N__12193;
    wire N__12190;
    wire N__12187;
    wire N__12186;
    wire N__12185;
    wire N__12184;
    wire N__12183;
    wire N__12180;
    wire N__12177;
    wire N__12174;
    wire N__12171;
    wire N__12170;
    wire N__12169;
    wire N__12164;
    wire N__12161;
    wire N__12144;
    wire N__12137;
    wire N__12134;
    wire N__12131;
    wire N__12128;
    wire N__12127;
    wire N__12124;
    wire N__12115;
    wire N__12110;
    wire N__12107;
    wire N__12104;
    wire N__12101;
    wire N__12098;
    wire N__12089;
    wire N__12086;
    wire N__12083;
    wire N__12080;
    wire N__12077;
    wire N__12074;
    wire N__12071;
    wire N__12068;
    wire N__12065;
    wire N__12062;
    wire N__12059;
    wire N__12056;
    wire N__12053;
    wire N__12050;
    wire N__12047;
    wire N__12044;
    wire N__12043;
    wire N__12042;
    wire N__12039;
    wire N__12036;
    wire N__12035;
    wire N__12032;
    wire N__12027;
    wire N__12024;
    wire N__12021;
    wire N__12016;
    wire N__12013;
    wire N__12010;
    wire N__12007;
    wire N__12004;
    wire N__11999;
    wire N__11996;
    wire N__11993;
    wire N__11992;
    wire N__11991;
    wire N__11988;
    wire N__11985;
    wire N__11982;
    wire N__11975;
    wire N__11972;
    wire N__11969;
    wire N__11966;
    wire N__11965;
    wire N__11964;
    wire N__11963;
    wire N__11962;
    wire N__11959;
    wire N__11954;
    wire N__11949;
    wire N__11942;
    wire N__11941;
    wire N__11940;
    wire N__11939;
    wire N__11938;
    wire N__11937;
    wire N__11936;
    wire N__11935;
    wire N__11934;
    wire N__11933;
    wire N__11932;
    wire N__11929;
    wire N__11928;
    wire N__11925;
    wire N__11922;
    wire N__11919;
    wire N__11916;
    wire N__11915;
    wire N__11914;
    wire N__11913;
    wire N__11912;
    wire N__11911;
    wire N__11908;
    wire N__11905;
    wire N__11904;
    wire N__11903;
    wire N__11902;
    wire N__11901;
    wire N__11898;
    wire N__11895;
    wire N__11892;
    wire N__11889;
    wire N__11888;
    wire N__11883;
    wire N__11882;
    wire N__11881;
    wire N__11866;
    wire N__11861;
    wire N__11856;
    wire N__11839;
    wire N__11836;
    wire N__11833;
    wire N__11828;
    wire N__11825;
    wire N__11820;
    wire N__11817;
    wire N__11814;
    wire N__11809;
    wire N__11806;
    wire N__11803;
    wire N__11800;
    wire N__11795;
    wire N__11786;
    wire N__11783;
    wire N__11780;
    wire N__11777;
    wire N__11774;
    wire N__11771;
    wire N__11768;
    wire N__11765;
    wire N__11762;
    wire N__11759;
    wire N__11756;
    wire N__11753;
    wire N__11750;
    wire N__11749;
    wire N__11746;
    wire N__11743;
    wire N__11742;
    wire N__11739;
    wire N__11736;
    wire N__11733;
    wire N__11726;
    wire N__11723;
    wire N__11720;
    wire N__11717;
    wire N__11714;
    wire N__11713;
    wire N__11712;
    wire N__11709;
    wire N__11708;
    wire N__11707;
    wire N__11706;
    wire N__11703;
    wire N__11702;
    wire N__11701;
    wire N__11700;
    wire N__11699;
    wire N__11696;
    wire N__11687;
    wire N__11676;
    wire N__11671;
    wire N__11668;
    wire N__11663;
    wire N__11660;
    wire N__11657;
    wire N__11654;
    wire N__11651;
    wire N__11650;
    wire N__11645;
    wire N__11644;
    wire N__11643;
    wire N__11640;
    wire N__11635;
    wire N__11634;
    wire N__11631;
    wire N__11628;
    wire N__11625;
    wire N__11618;
    wire N__11615;
    wire N__11612;
    wire N__11609;
    wire N__11606;
    wire N__11603;
    wire N__11600;
    wire N__11597;
    wire N__11594;
    wire N__11591;
    wire N__11588;
    wire N__11585;
    wire N__11582;
    wire N__11579;
    wire N__11576;
    wire N__11573;
    wire N__11570;
    wire N__11567;
    wire N__11564;
    wire N__11561;
    wire N__11558;
    wire N__11557;
    wire N__11556;
    wire N__11555;
    wire N__11550;
    wire N__11545;
    wire N__11542;
    wire N__11539;
    wire N__11534;
    wire N__11531;
    wire N__11528;
    wire N__11525;
    wire N__11522;
    wire N__11519;
    wire N__11518;
    wire N__11517;
    wire N__11516;
    wire N__11515;
    wire N__11514;
    wire N__11501;
    wire N__11498;
    wire N__11495;
    wire N__11494;
    wire N__11493;
    wire N__11492;
    wire N__11491;
    wire N__11490;
    wire N__11489;
    wire N__11486;
    wire N__11473;
    wire N__11468;
    wire N__11467;
    wire N__11464;
    wire N__11461;
    wire N__11458;
    wire N__11455;
    wire N__11450;
    wire N__11447;
    wire N__11444;
    wire N__11443;
    wire N__11442;
    wire N__11441;
    wire N__11440;
    wire N__11439;
    wire N__11438;
    wire N__11435;
    wire N__11434;
    wire N__11429;
    wire N__11416;
    wire N__11415;
    wire N__11414;
    wire N__11409;
    wire N__11408;
    wire N__11405;
    wire N__11404;
    wire N__11403;
    wire N__11402;
    wire N__11401;
    wire N__11398;
    wire N__11397;
    wire N__11394;
    wire N__11377;
    wire N__11372;
    wire N__11369;
    wire N__11366;
    wire N__11363;
    wire N__11360;
    wire N__11357;
    wire N__11354;
    wire N__11351;
    wire N__11348;
    wire N__11345;
    wire N__11342;
    wire N__11339;
    wire N__11336;
    wire N__11333;
    wire N__11330;
    wire N__11327;
    wire N__11324;
    wire N__11321;
    wire N__11318;
    wire N__11315;
    wire N__11312;
    wire N__11309;
    wire N__11306;
    wire N__11303;
    wire N__11300;
    wire N__11297;
    wire N__11294;
    wire N__11291;
    wire N__11288;
    wire N__11285;
    wire N__11282;
    wire N__11279;
    wire N__11276;
    wire N__11273;
    wire N__11270;
    wire N__11269;
    wire N__11266;
    wire N__11263;
    wire N__11262;
    wire N__11259;
    wire N__11256;
    wire N__11253;
    wire N__11250;
    wire N__11247;
    wire N__11244;
    wire N__11237;
    wire N__11234;
    wire N__11231;
    wire N__11228;
    wire N__11225;
    wire N__11222;
    wire N__11219;
    wire N__11216;
    wire N__11213;
    wire N__11210;
    wire N__11207;
    wire N__11204;
    wire N__11201;
    wire N__11198;
    wire N__11195;
    wire N__11192;
    wire N__11189;
    wire N__11186;
    wire N__11183;
    wire N__11180;
    wire N__11177;
    wire N__11174;
    wire N__11171;
    wire N__11168;
    wire N__11165;
    wire N__11162;
    wire N__11159;
    wire N__11156;
    wire N__11153;
    wire N__11150;
    wire N__11147;
    wire N__11146;
    wire N__11145;
    wire N__11142;
    wire N__11139;
    wire N__11136;
    wire N__11133;
    wire N__11130;
    wire N__11127;
    wire N__11120;
    wire N__11117;
    wire N__11116;
    wire N__11115;
    wire N__11110;
    wire N__11107;
    wire N__11104;
    wire N__11101;
    wire N__11098;
    wire N__11093;
    wire N__11090;
    wire N__11087;
    wire N__11084;
    wire N__11081;
    wire N__11080;
    wire N__11077;
    wire N__11076;
    wire N__11075;
    wire N__11072;
    wire N__11071;
    wire N__11068;
    wire N__11063;
    wire N__11060;
    wire N__11057;
    wire N__11050;
    wire N__11045;
    wire N__11044;
    wire N__11043;
    wire N__11042;
    wire N__11041;
    wire N__11038;
    wire N__11033;
    wire N__11028;
    wire N__11021;
    wire N__11018;
    wire N__11015;
    wire N__11012;
    wire N__11009;
    wire N__11006;
    wire N__11005;
    wire N__11004;
    wire N__11001;
    wire N__10998;
    wire N__10995;
    wire N__10988;
    wire N__10985;
    wire N__10982;
    wire N__10979;
    wire N__10976;
    wire N__10973;
    wire N__10970;
    wire N__10967;
    wire N__10964;
    wire N__10961;
    wire N__10958;
    wire N__10955;
    wire N__10952;
    wire N__10949;
    wire N__10946;
    wire N__10943;
    wire N__10940;
    wire N__10937;
    wire N__10934;
    wire N__10931;
    wire N__10928;
    wire N__10925;
    wire N__10922;
    wire N__10919;
    wire N__10916;
    wire N__10913;
    wire N__10910;
    wire N__10907;
    wire N__10904;
    wire N__10901;
    wire N__10898;
    wire N__10895;
    wire N__10892;
    wire N__10891;
    wire N__10890;
    wire N__10889;
    wire N__10888;
    wire N__10887;
    wire N__10886;
    wire N__10885;
    wire N__10884;
    wire N__10883;
    wire N__10882;
    wire N__10881;
    wire N__10880;
    wire N__10879;
    wire N__10876;
    wire N__10875;
    wire N__10874;
    wire N__10873;
    wire N__10872;
    wire N__10871;
    wire N__10870;
    wire N__10853;
    wire N__10846;
    wire N__10843;
    wire N__10842;
    wire N__10825;
    wire N__10822;
    wire N__10819;
    wire N__10818;
    wire N__10817;
    wire N__10816;
    wire N__10811;
    wire N__10806;
    wire N__10803;
    wire N__10800;
    wire N__10797;
    wire N__10794;
    wire N__10781;
    wire N__10780;
    wire N__10779;
    wire N__10778;
    wire N__10777;
    wire N__10776;
    wire N__10775;
    wire N__10774;
    wire N__10773;
    wire N__10772;
    wire N__10771;
    wire N__10770;
    wire N__10769;
    wire N__10768;
    wire N__10767;
    wire N__10766;
    wire N__10765;
    wire N__10764;
    wire N__10763;
    wire N__10746;
    wire N__10729;
    wire N__10722;
    wire N__10721;
    wire N__10720;
    wire N__10715;
    wire N__10712;
    wire N__10711;
    wire N__10710;
    wire N__10709;
    wire N__10704;
    wire N__10699;
    wire N__10696;
    wire N__10693;
    wire N__10690;
    wire N__10679;
    wire N__10676;
    wire N__10673;
    wire N__10670;
    wire N__10667;
    wire N__10664;
    wire N__10661;
    wire N__10658;
    wire N__10655;
    wire N__10652;
    wire N__10649;
    wire N__10646;
    wire N__10643;
    wire N__10640;
    wire N__10637;
    wire N__10634;
    wire N__10631;
    wire N__10628;
    wire N__10625;
    wire N__10622;
    wire N__10619;
    wire N__10618;
    wire N__10615;
    wire N__10612;
    wire N__10609;
    wire N__10604;
    wire N__10601;
    wire N__10598;
    wire N__10595;
    wire N__10594;
    wire N__10591;
    wire N__10588;
    wire N__10585;
    wire N__10580;
    wire N__10577;
    wire N__10574;
    wire N__10571;
    wire N__10570;
    wire N__10567;
    wire N__10564;
    wire N__10561;
    wire N__10556;
    wire N__10553;
    wire N__10550;
    wire N__10547;
    wire N__10546;
    wire N__10543;
    wire N__10540;
    wire N__10537;
    wire N__10532;
    wire N__10529;
    wire N__10526;
    wire N__10523;
    wire N__10522;
    wire N__10519;
    wire N__10516;
    wire N__10511;
    wire N__10508;
    wire N__10505;
    wire N__10502;
    wire N__10501;
    wire N__10498;
    wire N__10495;
    wire N__10490;
    wire N__10487;
    wire N__10484;
    wire N__10481;
    wire N__10480;
    wire N__10477;
    wire N__10474;
    wire N__10469;
    wire N__10466;
    wire N__10463;
    wire N__10460;
    wire N__10459;
    wire N__10456;
    wire N__10453;
    wire N__10448;
    wire N__10445;
    wire N__10442;
    wire N__10439;
    wire N__10438;
    wire N__10435;
    wire N__10432;
    wire N__10427;
    wire N__10424;
    wire N__10421;
    wire N__10418;
    wire N__10417;
    wire N__10414;
    wire N__10411;
    wire N__10406;
    wire N__10403;
    wire N__10400;
    wire N__10397;
    wire N__10396;
    wire N__10393;
    wire N__10390;
    wire N__10385;
    wire N__10382;
    wire N__10379;
    wire N__10376;
    wire N__10373;
    wire N__10372;
    wire N__10369;
    wire N__10366;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10352;
    wire N__10349;
    wire N__10348;
    wire N__10345;
    wire N__10342;
    wire N__10337;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10325;
    wire N__10324;
    wire N__10321;
    wire N__10318;
    wire N__10313;
    wire N__10310;
    wire N__10307;
    wire N__10304;
    wire N__10303;
    wire N__10300;
    wire N__10297;
    wire N__10294;
    wire N__10291;
    wire N__10286;
    wire N__10283;
    wire N__10280;
    wire N__10277;
    wire N__10274;
    wire N__10271;
    wire N__10268;
    wire N__10265;
    wire N__10262;
    wire N__10259;
    wire N__10256;
    wire N__10253;
    wire N__10250;
    wire N__10247;
    wire N__10244;
    wire N__10241;
    wire N__10240;
    wire N__10237;
    wire N__10236;
    wire N__10233;
    wire N__10230;
    wire N__10227;
    wire N__10220;
    wire N__10217;
    wire N__10214;
    wire N__10211;
    wire N__10210;
    wire N__10207;
    wire N__10204;
    wire N__10199;
    wire N__10196;
    wire N__10193;
    wire N__10192;
    wire N__10189;
    wire N__10186;
    wire N__10181;
    wire N__10178;
    wire N__10175;
    wire N__10172;
    wire N__10171;
    wire N__10168;
    wire N__10165;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10151;
    wire N__10148;
    wire N__10145;
    wire N__10142;
    wire N__10139;
    wire N__10136;
    wire N__10133;
    wire N__10130;
    wire N__10129;
    wire N__10126;
    wire N__10125;
    wire N__10122;
    wire N__10119;
    wire N__10116;
    wire N__10109;
    wire N__10106;
    wire N__10103;
    wire N__10100;
    wire N__10097;
    wire N__10094;
    wire N__10091;
    wire N__10088;
    wire N__10085;
    wire N__10082;
    wire N__10079;
    wire N__10076;
    wire N__10073;
    wire N__10070;
    wire N__10067;
    wire N__10064;
    wire N__10061;
    wire N__10058;
    wire N__10057;
    wire N__10054;
    wire N__10051;
    wire N__10046;
    wire N__10043;
    wire N__10040;
    wire N__10037;
    wire N__10036;
    wire N__10033;
    wire N__10030;
    wire N__10025;
    wire N__10022;
    wire N__10019;
    wire N__10016;
    wire N__10015;
    wire N__10012;
    wire N__10009;
    wire N__10004;
    wire N__10001;
    wire N__9998;
    wire N__9995;
    wire N__9994;
    wire N__9991;
    wire N__9988;
    wire N__9983;
    wire N__9980;
    wire N__9977;
    wire N__9974;
    wire N__9971;
    wire N__9968;
    wire N__9967;
    wire N__9964;
    wire N__9961;
    wire N__9956;
    wire N__9953;
    wire N__9950;
    wire N__9947;
    wire N__9944;
    wire N__9941;
    wire N__9940;
    wire N__9937;
    wire N__9934;
    wire N__9929;
    wire N__9926;
    wire N__9923;
    wire N__9920;
    wire N__9917;
    wire N__9914;
    wire N__9913;
    wire N__9910;
    wire N__9907;
    wire N__9902;
    wire N__9899;
    wire N__9896;
    wire N__9893;
    wire N__9892;
    wire N__9889;
    wire N__9886;
    wire N__9881;
    wire N__9878;
    wire N__9875;
    wire N__9872;
    wire N__9871;
    wire N__9868;
    wire N__9865;
    wire N__9860;
    wire N__9857;
    wire N__9854;
    wire N__9851;
    wire N__9850;
    wire N__9847;
    wire N__9844;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9830;
    wire N__9829;
    wire N__9826;
    wire N__9823;
    wire N__9818;
    wire N__9815;
    wire N__9812;
    wire N__9809;
    wire N__9808;
    wire N__9805;
    wire N__9802;
    wire N__9797;
    wire N__9794;
    wire N__9791;
    wire N__9788;
    wire N__9787;
    wire N__9784;
    wire N__9781;
    wire N__9776;
    wire N__9773;
    wire N__9770;
    wire N__9767;
    wire N__9766;
    wire N__9763;
    wire N__9760;
    wire N__9757;
    wire N__9752;
    wire N__9749;
    wire N__9746;
    wire N__9743;
    wire N__9742;
    wire N__9739;
    wire N__9736;
    wire N__9731;
    wire N__9728;
    wire N__9725;
    wire N__9722;
    wire N__9721;
    wire N__9720;
    wire N__9717;
    wire N__9714;
    wire N__9711;
    wire N__9710;
    wire N__9709;
    wire N__9708;
    wire N__9707;
    wire N__9706;
    wire N__9705;
    wire N__9704;
    wire N__9703;
    wire N__9702;
    wire N__9701;
    wire N__9700;
    wire N__9699;
    wire N__9698;
    wire N__9697;
    wire N__9696;
    wire N__9695;
    wire N__9688;
    wire N__9679;
    wire N__9678;
    wire N__9677;
    wire N__9668;
    wire N__9651;
    wire N__9646;
    wire N__9645;
    wire N__9644;
    wire N__9643;
    wire N__9638;
    wire N__9631;
    wire N__9626;
    wire N__9623;
    wire N__9614;
    wire N__9613;
    wire N__9612;
    wire N__9611;
    wire N__9610;
    wire N__9609;
    wire N__9608;
    wire N__9607;
    wire N__9606;
    wire N__9605;
    wire N__9604;
    wire N__9603;
    wire N__9602;
    wire N__9601;
    wire N__9600;
    wire N__9599;
    wire N__9598;
    wire N__9595;
    wire N__9594;
    wire N__9593;
    wire N__9592;
    wire N__9575;
    wire N__9560;
    wire N__9557;
    wire N__9556;
    wire N__9547;
    wire N__9542;
    wire N__9541;
    wire N__9540;
    wire N__9539;
    wire N__9534;
    wire N__9531;
    wire N__9528;
    wire N__9523;
    wire N__9520;
    wire N__9509;
    wire N__9508;
    wire N__9507;
    wire N__9506;
    wire N__9505;
    wire N__9504;
    wire N__9503;
    wire N__9494;
    wire N__9493;
    wire N__9492;
    wire N__9491;
    wire N__9490;
    wire N__9489;
    wire N__9488;
    wire N__9487;
    wire N__9486;
    wire N__9485;
    wire N__9484;
    wire N__9483;
    wire N__9482;
    wire N__9481;
    wire N__9480;
    wire N__9479;
    wire N__9476;
    wire N__9475;
    wire N__9474;
    wire N__9469;
    wire N__9466;
    wire N__9449;
    wire N__9434;
    wire N__9431;
    wire N__9426;
    wire N__9413;
    wire N__9412;
    wire N__9411;
    wire N__9410;
    wire N__9409;
    wire N__9408;
    wire N__9407;
    wire N__9406;
    wire N__9403;
    wire N__9400;
    wire N__9397;
    wire N__9394;
    wire N__9393;
    wire N__9392;
    wire N__9391;
    wire N__9390;
    wire N__9387;
    wire N__9384;
    wire N__9381;
    wire N__9378;
    wire N__9377;
    wire N__9376;
    wire N__9375;
    wire N__9374;
    wire N__9373;
    wire N__9372;
    wire N__9371;
    wire N__9370;
    wire N__9369;
    wire N__9360;
    wire N__9351;
    wire N__9350;
    wire N__9349;
    wire N__9348;
    wire N__9339;
    wire N__9334;
    wire N__9325;
    wire N__9318;
    wire N__9313;
    wire N__9310;
    wire N__9305;
    wire N__9290;
    wire N__9287;
    wire N__9284;
    wire N__9281;
    wire N__9278;
    wire N__9277;
    wire N__9274;
    wire N__9271;
    wire N__9266;
    wire N__9263;
    wire N__9260;
    wire N__9257;
    wire N__9254;
    wire N__9253;
    wire N__9250;
    wire N__9247;
    wire N__9242;
    wire N__9239;
    wire N__9236;
    wire N__9233;
    wire N__9232;
    wire N__9229;
    wire N__9226;
    wire N__9221;
    wire N__9218;
    wire N__9215;
    wire N__9212;
    wire N__9211;
    wire N__9208;
    wire N__9205;
    wire N__9200;
    wire N__9197;
    wire N__9194;
    wire N__9191;
    wire N__9190;
    wire N__9187;
    wire N__9184;
    wire N__9179;
    wire N__9176;
    wire N__9173;
    wire N__9170;
    wire N__9167;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9157;
    wire N__9154;
    wire N__9151;
    wire N__9146;
    wire N__9143;
    wire N__9140;
    wire N__9137;
    wire N__9136;
    wire N__9133;
    wire N__9130;
    wire N__9125;
    wire N__9122;
    wire N__9119;
    wire N__9116;
    wire N__9113;
    wire N__9110;
    wire N__9107;
    wire N__9104;
    wire N__9101;
    wire N__9098;
    wire N__9095;
    wire N__9092;
    wire N__9089;
    wire N__9086;
    wire N__9083;
    wire N__9082;
    wire N__9079;
    wire N__9076;
    wire N__9071;
    wire N__9068;
    wire N__9065;
    wire N__9062;
    wire N__9061;
    wire N__9058;
    wire N__9055;
    wire N__9050;
    wire N__9047;
    wire N__9044;
    wire N__9041;
    wire N__9040;
    wire N__9037;
    wire N__9034;
    wire N__9029;
    wire N__9026;
    wire N__9023;
    wire N__9020;
    wire N__9019;
    wire N__9016;
    wire N__9013;
    wire N__9008;
    wire N__9005;
    wire N__9002;
    wire N__8999;
    wire N__8998;
    wire N__8995;
    wire N__8992;
    wire N__8987;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8977;
    wire N__8974;
    wire N__8971;
    wire N__8966;
    wire N__8963;
    wire N__8960;
    wire N__8957;
    wire N__8956;
    wire N__8953;
    wire N__8950;
    wire N__8945;
    wire N__8942;
    wire N__8939;
    wire N__8936;
    wire N__8935;
    wire N__8932;
    wire N__8929;
    wire N__8924;
    wire N__8921;
    wire N__8918;
    wire N__8915;
    wire N__8914;
    wire N__8911;
    wire N__8910;
    wire N__8907;
    wire N__8904;
    wire N__8901;
    wire N__8894;
    wire N__8891;
    wire N__8888;
    wire N__8885;
    wire N__8884;
    wire N__8881;
    wire N__8878;
    wire N__8873;
    wire N__8870;
    wire N__8867;
    wire N__8864;
    wire N__8863;
    wire N__8860;
    wire N__8857;
    wire N__8852;
    wire N__8849;
    wire N__8846;
    wire N__8843;
    wire N__8842;
    wire N__8839;
    wire N__8836;
    wire N__8831;
    wire N__8828;
    wire N__8825;
    wire N__8822;
    wire N__8821;
    wire N__8818;
    wire N__8815;
    wire N__8810;
    wire N__8807;
    wire N__8804;
    wire N__8801;
    wire N__8800;
    wire N__8797;
    wire N__8794;
    wire N__8789;
    wire N__8786;
    wire N__8783;
    wire N__8780;
    wire N__8779;
    wire N__8776;
    wire N__8773;
    wire N__8768;
    wire N__8765;
    wire N__8762;
    wire N__8759;
    wire N__8756;
    wire N__8753;
    wire N__8750;
    wire N__8747;
    wire N__8744;
    wire N__8741;
    wire N__8738;
    wire N__8735;
    wire N__8732;
    wire N__8729;
    wire N__8726;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8711;
    wire N__8708;
    wire N__8705;
    wire N__8702;
    wire N__8699;
    wire N__8696;
    wire N__8693;
    wire N__8690;
    wire N__8687;
    wire N__8684;
    wire N__8681;
    wire N__8678;
    wire N__8675;
    wire N__8672;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8618;
    wire N__8615;
    wire N__8612;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8600;
    wire N__8597;
    wire N__8594;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire N__8570;
    wire N__8567;
    wire N__8564;
    wire N__8561;
    wire N__8558;
    wire N__8555;
    wire N__8552;
    wire N__8549;
    wire N__8546;
    wire N__8543;
    wire N__8540;
    wire N__8537;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8525;
    wire N__8522;
    wire N__8519;
    wire N__8516;
    wire N__8513;
    wire N__8510;
    wire N__8507;
    wire N__8504;
    wire N__8501;
    wire N__8498;
    wire N__8495;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8474;
    wire N__8471;
    wire N__8468;
    wire N__8465;
    wire N__8462;
    wire N__8459;
    wire N__8456;
    wire N__8453;
    wire N__8450;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8438;
    wire N__8435;
    wire N__8432;
    wire N__8429;
    wire N__8426;
    wire N__8423;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8408;
    wire N__8405;
    wire N__8402;
    wire N__8399;
    wire N__8396;
    wire N__8393;
    wire N__8390;
    wire N__8387;
    wire N__8384;
    wire N__8381;
    wire N__8378;
    wire N__8375;
    wire N__8372;
    wire N__8369;
    wire N__8366;
    wire N__8363;
    wire N__8360;
    wire N__8357;
    wire N__8354;
    wire N__8351;
    wire N__8348;
    wire N__8345;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8333;
    wire N__8330;
    wire N__8327;
    wire N__8324;
    wire N__8321;
    wire N__8318;
    wire N__8315;
    wire N__8312;
    wire N__8309;
    wire N__8306;
    wire N__8303;
    wire N__8302;
    wire N__8301;
    wire N__8300;
    wire N__8297;
    wire N__8294;
    wire N__8291;
    wire N__8288;
    wire N__8279;
    wire N__8276;
    wire N__8273;
    wire N__8270;
    wire N__8267;
    wire N__8264;
    wire N__8261;
    wire N__8258;
    wire N__8255;
    wire N__8252;
    wire N__8249;
    wire N__8246;
    wire N__8243;
    wire N__8240;
    wire N__8237;
    wire N__8234;
    wire N__8231;
    wire N__8228;
    wire N__8225;
    wire N__8222;
    wire N__8219;
    wire N__8216;
    wire N__8213;
    wire N__8210;
    wire N__8207;
    wire N__8204;
    wire N__8201;
    wire N__8198;
    wire GNDG0;
    wire VCCG0;
    wire bfn_1_14_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ;
    wire bfn_1_15_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ;
    wire bfn_1_16_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ;
    wire bfn_1_17_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ;
    wire bfn_1_18_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ;
    wire bfn_1_19_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ;
    wire CONSTANT_ONE_NET;
    wire rgb_drv_RNOZ0;
    wire N_39_i_i;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0 ;
    wire \phase_controller_inst1.stoper_tr.time_passed11_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ;
    wire \phase_controller_inst1.stoper_hc.time_passed11_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ;
    wire bfn_2_23_0_;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7 ;
    wire bfn_2_24_0_;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15 ;
    wire bfn_2_25_0_;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11 ;
    wire \phase_controller_slave.stoper_hc.time_passed11_cascade_ ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire bfn_3_15_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire bfn_3_16_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_17 ;
    wire bfn_3_17_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ;
    wire \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_3_19_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_3_20_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_17 ;
    wire bfn_3_21_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_1 ;
    wire bfn_3_25_0_;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_9 ;
    wire bfn_3_26_0_;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_16 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_17 ;
    wire bfn_3_27_0_;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_ ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ;
    wire \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ;
    wire \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ;
    wire \phase_controller_inst1.stoper_tr.time_passed11 ;
    wire \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ;
    wire \phase_controller_inst1.stoper_hc.time_passed11 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ;
    wire \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_4Z0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_3Z0Z_3_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.N_144_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_0Z0Z_6_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2Z0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2Z0Z_9_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_time_6_i_o2Z0Z_15_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_1Z0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_ ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.N_122 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a3_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.N_144 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2Z0Z_6 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_0Z0Z_6 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2Z0Z_9 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.target_time_6_i_o2Z0Z_15 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ;
    wire \phase_controller_slave.stoper_hc.time_passed11 ;
    wire \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire \phase_controller_inst1.N_110 ;
    wire \phase_controller_inst1.N_112 ;
    wire \phase_controller_inst1.tr_time_passed ;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire \phase_controller_inst1.hc_time_passed ;
    wire \phase_controller_inst1.stateZ0Z_4 ;
    wire \phase_controller_inst1.N_107 ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_1 ;
    wire bfn_5_17_0_;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_9 ;
    wire bfn_5_18_0_;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_17 ;
    wire bfn_5_19_0_;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_ ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.N_38 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ;
    wire \phase_controller_slave.start_timer_tr_0_sqmuxa ;
    wire \phase_controller_slave.tr_time_passed ;
    wire \phase_controller_slave.stateZ0Z_0 ;
    wire \phase_controller_slave.state_RNIVDE2Z0Z_0 ;
    wire start_stop_c;
    wire shift_flag_start;
    wire il_max_comp2_c;
    wire il_max_comp2_D1;
    wire \phase_controller_slave.state_RNO_0Z0Z_3 ;
    wire il_max_comp2_D2;
    wire \phase_controller_slave.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_slave.stateZ0Z_4 ;
    wire \phase_controller_slave.start_timer_hcZ0 ;
    wire \phase_controller_slave.stateZ0Z_2 ;
    wire \phase_controller_slave.hc_time_passed ;
    wire \phase_controller_slave.start_timer_hc_RNOZ0Z_0 ;
    wire il_max_comp1_c;
    wire il_min_comp2_c;
    wire il_max_comp1_D1;
    wire il_max_comp1_D2;
    wire \phase_controller_inst1.start_timer_hc_0_sqmuxa ;
    wire il_min_comp1_c;
    wire il_min_comp1_D1;
    wire il_min_comp1_D2;
    wire \phase_controller_inst1.T01_0_sqmuxa ;
    wire \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa ;
    wire il_min_comp2_D1;
    wire il_min_comp2_D2;
    wire measured_delay_hc_5;
    wire measured_delay_hc_2;
    wire measured_delay_hc_11;
    wire measured_delay_hc_12;
    wire measured_delay_hc_3;
    wire measured_delay_hc_4;
    wire \delay_measurement_inst.delay_hc_reg_3_0_a2_0_6 ;
    wire measured_delay_hc_1;
    wire measured_delay_hc_10;
    wire measured_delay_hc_9;
    wire measured_delay_hc_15;
    wire measured_delay_hc_19;
    wire measured_delay_hc_6;
    wire measured_delay_hc_17;
    wire measured_delay_hc_16;
    wire measured_delay_hc_14;
    wire measured_delay_hc_18;
    wire measured_delay_hc_7;
    wire measured_delay_hc_8;
    wire bfn_8_13_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire bfn_8_14_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire bfn_8_15_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire bfn_8_16_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.N_256_i_g ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ;
    wire bfn_8_17_0_;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9 ;
    wire bfn_8_18_0_;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17 ;
    wire bfn_8_19_0_;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19 ;
    wire \phase_controller_inst1.stoper_tr.N_55 ;
    wire \phase_controller_slave.stoper_tr.time_passed11 ;
    wire \phase_controller_inst1.stoper_tr.N_50 ;
    wire \phase_controller_inst1.stoper_tr.N_32 ;
    wire \phase_controller_inst1.stoper_tr.N_32_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.N_33 ;
    wire \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ;
    wire \phase_controller_slave.start_timer_trZ0 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ;
    wire \delay_measurement_inst.elapsed_time_hc_1 ;
    wire \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_0_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_0_3 ;
    wire \delay_measurement_inst.elapsed_time_hc_2 ;
    wire \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_3_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.N_232_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_2 ;
    wire \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_6_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_0_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_7 ;
    wire \delay_measurement_inst.un3_elapsed_time_hc_0_i ;
    wire \delay_measurement_inst.un3_elapsed_time_hc_0_i_cascade_ ;
    wire \delay_measurement_inst.N_219 ;
    wire \delay_measurement_inst.delay_hc_timer.N_237_cascade_ ;
    wire \delay_measurement_inst.N_209 ;
    wire \delay_measurement_inst.N_207 ;
    wire \delay_measurement_inst.N_207_cascade_ ;
    wire \delay_measurement_inst.N_243 ;
    wire \delay_measurement_inst.N_247 ;
    wire \delay_measurement_inst.N_216_1 ;
    wire measured_delay_hc_13;
    wire \delay_measurement_inst.un3_elapsed_time_hc_0_i_0 ;
    wire \phase_controller_slave.stateZ0Z_1 ;
    wire s4_phy_c;
    wire bfn_9_13_0_;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire bfn_9_14_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire bfn_9_15_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire bfn_9_16_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire measured_delay_tr_1;
    wire measured_delay_tr_2;
    wire measured_delay_tr_3;
    wire measured_delay_tr_6;
    wire measured_delay_tr_18;
    wire measured_delay_tr_17;
    wire measured_delay_tr_16;
    wire measured_delay_tr_12;
    wire measured_delay_tr_11;
    wire measured_delay_tr_13;
    wire measured_delay_tr_10;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_0_6 ;
    wire measured_delay_tr_9;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_0_6_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_9 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_9_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_0_6 ;
    wire \phase_controller_inst1.stoper_tr.N_97 ;
    wire measured_delay_tr_4;
    wire measured_delay_tr_14;
    wire measured_delay_tr_15;
    wire measured_delay_tr_5;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3 ;
    wire \phase_controller_inst1.stateZ0Z_3 ;
    wire s1_phy_c;
    wire bfn_9_21_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire bfn_9_22_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire bfn_9_23_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire bfn_9_24_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \phase_controller_slave.stateZ0Z_3 ;
    wire s3_phy_c;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.N_255_i_g ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \delay_measurement_inst.elapsed_time_tr_5 ;
    wire \delay_measurement_inst.elapsed_time_tr_4 ;
    wire \delay_measurement_inst.elapsed_time_tr_3 ;
    wire \delay_measurement_inst.elapsed_time_tr_1 ;
    wire \delay_measurement_inst.elapsed_time_tr_2 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_177_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3_cascade_ ;
    wire \delay_measurement_inst.elapsed_time_tr_16 ;
    wire \delay_measurement_inst.elapsed_time_tr_17 ;
    wire \delay_measurement_inst.elapsed_time_tr_18 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire \delay_measurement_inst.elapsed_time_tr_12 ;
    wire \delay_measurement_inst.elapsed_time_tr_11 ;
    wire \delay_measurement_inst.elapsed_time_tr_13 ;
    wire \delay_measurement_inst.elapsed_time_tr_10 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19 ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6 ;
    wire \delay_measurement_inst.N_35_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_7 ;
    wire \delay_measurement_inst.N_164 ;
    wire \delay_measurement_inst.N_187 ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_7 ;
    wire \delay_measurement_inst.N_187_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_177 ;
    wire \delay_measurement_inst.un3_elapsed_time_tr_0_i_cascade_ ;
    wire \delay_measurement_inst.N_162_1 ;
    wire \delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10 ;
    wire \delay_measurement_inst.delay_tr_reg3lto9 ;
    wire \delay_measurement_inst.delay_tr_reg3lto14 ;
    wire \delay_measurement_inst.N_39 ;
    wire \delay_measurement_inst.delay_tr_timer.N_180_cascade_ ;
    wire \delay_measurement_inst.delay_tr_reg3lto6 ;
    wire \delay_measurement_inst.delay_tr_reg3lto15 ;
    wire \delay_measurement_inst.delay_tr_reg_5_0_a2_0_6 ;
    wire \delay_measurement_inst.elapsed_time_tr_7 ;
    wire measured_delay_tr_7;
    wire \delay_measurement_inst.un3_elapsed_time_tr_0_i ;
    wire \delay_measurement_inst.N_41 ;
    wire \delay_measurement_inst.elapsed_time_tr_8 ;
    wire measured_delay_tr_8;
    wire \delay_measurement_inst.elapsed_time_tr_31 ;
    wire \delay_measurement_inst.elapsed_time_tr_19 ;
    wire \delay_measurement_inst.N_35 ;
    wire measured_delay_tr_19;
    wire \delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.elapsed_time_hc_3 ;
    wire bfn_10_21_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.elapsed_time_hc_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.elapsed_time_hc_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_reg3lto6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.elapsed_time_hc_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.elapsed_time_hc_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_reg3lto9 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.elapsed_time_hc_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire \delay_measurement_inst.elapsed_time_hc_11 ;
    wire bfn_10_22_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.elapsed_time_hc_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.elapsed_time_hc_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_reg3lto14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_reg3lto15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.elapsed_time_hc_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.elapsed_time_hc_17 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.elapsed_time_hc_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire \delay_measurement_inst.elapsed_time_hc_19 ;
    wire bfn_10_23_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire bfn_10_24_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.elapsed_time_hc_31 ;
    wire \delay_measurement_inst.delay_hc_timer.N_253_i_g ;
    wire \delay_measurement_inst.delay_tr_timer.N_255_i ;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire s2_phy_c;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_7_19_cascade_ ;
    wire \delay_measurement_inst.N_276 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_6_19 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_0_19 ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.N_256_i ;
    wire delay_tr_input_c;
    wire delay_tr_d1;
    wire delay_tr_d2;
    wire \delay_measurement_inst.prev_tr_sigZ0 ;
    wire \delay_measurement_inst.tr_stateZ0Z_0 ;
    wire delay_hc_input_c;
    wire delay_hc_d1;
    wire \delay_measurement_inst.prev_hc_sigZ0 ;
    wire \delay_measurement_inst.hc_stateZ0Z_0 ;
    wire delay_hc_d2;
    wire clk_100mhz;
    wire \delay_measurement_inst.delay_hc_timer.N_253_i ;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.N_254_i_g ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire red_c_g;
    wire red_c_i;
    wire _gnd_net_;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__10667),
            .RESETB(N__20181),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clk_100mhz));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__21135),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__21137),
            .DIN(N__21136),
            .DOUT(N__21135),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__21137),
            .PADOUT(N__21136),
            .PADIN(N__21135),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__21126),
            .DIN(N__21125),
            .DOUT(N__21124),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__21126),
            .PADOUT(N__21125),
            .PADIN(N__21124),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__21117),
            .DIN(N__21116),
            .DOUT(N__21115),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__21117),
            .PADOUT(N__21116),
            .PADIN(N__21115),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__16859),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__21108),
            .DIN(N__21107),
            .DOUT(N__21106),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__21108),
            .PADOUT(N__21107),
            .PADIN(N__21106),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__15671),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__21099),
            .DIN(N__21098),
            .DOUT(N__21097),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__21099),
            .PADOUT(N__21098),
            .PADIN(N__21097),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__21090),
            .DIN(N__21089),
            .DOUT(N__21088),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__21090),
            .PADOUT(N__21089),
            .PADIN(N__21088),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__21081),
            .DIN(N__21080),
            .DOUT(N__21079),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__21081),
            .PADOUT(N__21080),
            .PADIN(N__21079),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__21072),
            .DIN(N__21071),
            .DOUT(N__21070),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__21072),
            .PADOUT(N__21071),
            .PADIN(N__21070),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__21063),
            .DIN(N__21062),
            .DOUT(N__21061),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__21063),
            .PADOUT(N__21062),
            .PADIN(N__21061),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__21054),
            .DIN(N__21053),
            .DOUT(N__21052),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__21054),
            .PADOUT(N__21053),
            .PADIN(N__21052),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__19883),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__21045),
            .DIN(N__21044),
            .DOUT(N__21043),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__21045),
            .PADOUT(N__21044),
            .PADIN(N__21043),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17243),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_iopad (
            .OE(N__21036),
            .DIN(N__21035),
            .DOUT(N__21034),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_preio (
            .PADOEN(N__21036),
            .PADOUT(N__21035),
            .PADIN(N__21034),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_iopad (
            .OE(N__21027),
            .DIN(N__21026),
            .DOUT(N__21025),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_preio (
            .PADOEN(N__21027),
            .PADOUT(N__21026),
            .PADIN(N__21025),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__4965 (
            .O(N__21008),
            .I(N__21005));
    LocalMux I__4964 (
            .O(N__21005),
            .I(N__21000));
    InMux I__4963 (
            .O(N__21004),
            .I(N__20997));
    InMux I__4962 (
            .O(N__21003),
            .I(N__20994));
    Odrv4 I__4961 (
            .O(N__21000),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    LocalMux I__4960 (
            .O(N__20997),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    LocalMux I__4959 (
            .O(N__20994),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    InMux I__4958 (
            .O(N__20987),
            .I(N__20984));
    LocalMux I__4957 (
            .O(N__20984),
            .I(N__20979));
    InMux I__4956 (
            .O(N__20983),
            .I(N__20976));
    InMux I__4955 (
            .O(N__20982),
            .I(N__20973));
    Odrv4 I__4954 (
            .O(N__20979),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    LocalMux I__4953 (
            .O(N__20976),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    LocalMux I__4952 (
            .O(N__20973),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    InMux I__4951 (
            .O(N__20966),
            .I(N__20959));
    InMux I__4950 (
            .O(N__20965),
            .I(N__20959));
    InMux I__4949 (
            .O(N__20964),
            .I(N__20956));
    LocalMux I__4948 (
            .O(N__20959),
            .I(N__20950));
    LocalMux I__4947 (
            .O(N__20956),
            .I(N__20950));
    InMux I__4946 (
            .O(N__20955),
            .I(N__20947));
    Odrv4 I__4945 (
            .O(N__20950),
            .I(delay_hc_d2));
    LocalMux I__4944 (
            .O(N__20947),
            .I(delay_hc_d2));
    ClkMux I__4943 (
            .O(N__20942),
            .I(N__20705));
    ClkMux I__4942 (
            .O(N__20941),
            .I(N__20705));
    ClkMux I__4941 (
            .O(N__20940),
            .I(N__20705));
    ClkMux I__4940 (
            .O(N__20939),
            .I(N__20705));
    ClkMux I__4939 (
            .O(N__20938),
            .I(N__20705));
    ClkMux I__4938 (
            .O(N__20937),
            .I(N__20705));
    ClkMux I__4937 (
            .O(N__20936),
            .I(N__20705));
    ClkMux I__4936 (
            .O(N__20935),
            .I(N__20705));
    ClkMux I__4935 (
            .O(N__20934),
            .I(N__20705));
    ClkMux I__4934 (
            .O(N__20933),
            .I(N__20705));
    ClkMux I__4933 (
            .O(N__20932),
            .I(N__20705));
    ClkMux I__4932 (
            .O(N__20931),
            .I(N__20705));
    ClkMux I__4931 (
            .O(N__20930),
            .I(N__20705));
    ClkMux I__4930 (
            .O(N__20929),
            .I(N__20705));
    ClkMux I__4929 (
            .O(N__20928),
            .I(N__20705));
    ClkMux I__4928 (
            .O(N__20927),
            .I(N__20705));
    ClkMux I__4927 (
            .O(N__20926),
            .I(N__20705));
    ClkMux I__4926 (
            .O(N__20925),
            .I(N__20705));
    ClkMux I__4925 (
            .O(N__20924),
            .I(N__20705));
    ClkMux I__4924 (
            .O(N__20923),
            .I(N__20705));
    ClkMux I__4923 (
            .O(N__20922),
            .I(N__20705));
    ClkMux I__4922 (
            .O(N__20921),
            .I(N__20705));
    ClkMux I__4921 (
            .O(N__20920),
            .I(N__20705));
    ClkMux I__4920 (
            .O(N__20919),
            .I(N__20705));
    ClkMux I__4919 (
            .O(N__20918),
            .I(N__20705));
    ClkMux I__4918 (
            .O(N__20917),
            .I(N__20705));
    ClkMux I__4917 (
            .O(N__20916),
            .I(N__20705));
    ClkMux I__4916 (
            .O(N__20915),
            .I(N__20705));
    ClkMux I__4915 (
            .O(N__20914),
            .I(N__20705));
    ClkMux I__4914 (
            .O(N__20913),
            .I(N__20705));
    ClkMux I__4913 (
            .O(N__20912),
            .I(N__20705));
    ClkMux I__4912 (
            .O(N__20911),
            .I(N__20705));
    ClkMux I__4911 (
            .O(N__20910),
            .I(N__20705));
    ClkMux I__4910 (
            .O(N__20909),
            .I(N__20705));
    ClkMux I__4909 (
            .O(N__20908),
            .I(N__20705));
    ClkMux I__4908 (
            .O(N__20907),
            .I(N__20705));
    ClkMux I__4907 (
            .O(N__20906),
            .I(N__20705));
    ClkMux I__4906 (
            .O(N__20905),
            .I(N__20705));
    ClkMux I__4905 (
            .O(N__20904),
            .I(N__20705));
    ClkMux I__4904 (
            .O(N__20903),
            .I(N__20705));
    ClkMux I__4903 (
            .O(N__20902),
            .I(N__20705));
    ClkMux I__4902 (
            .O(N__20901),
            .I(N__20705));
    ClkMux I__4901 (
            .O(N__20900),
            .I(N__20705));
    ClkMux I__4900 (
            .O(N__20899),
            .I(N__20705));
    ClkMux I__4899 (
            .O(N__20898),
            .I(N__20705));
    ClkMux I__4898 (
            .O(N__20897),
            .I(N__20705));
    ClkMux I__4897 (
            .O(N__20896),
            .I(N__20705));
    ClkMux I__4896 (
            .O(N__20895),
            .I(N__20705));
    ClkMux I__4895 (
            .O(N__20894),
            .I(N__20705));
    ClkMux I__4894 (
            .O(N__20893),
            .I(N__20705));
    ClkMux I__4893 (
            .O(N__20892),
            .I(N__20705));
    ClkMux I__4892 (
            .O(N__20891),
            .I(N__20705));
    ClkMux I__4891 (
            .O(N__20890),
            .I(N__20705));
    ClkMux I__4890 (
            .O(N__20889),
            .I(N__20705));
    ClkMux I__4889 (
            .O(N__20888),
            .I(N__20705));
    ClkMux I__4888 (
            .O(N__20887),
            .I(N__20705));
    ClkMux I__4887 (
            .O(N__20886),
            .I(N__20705));
    ClkMux I__4886 (
            .O(N__20885),
            .I(N__20705));
    ClkMux I__4885 (
            .O(N__20884),
            .I(N__20705));
    ClkMux I__4884 (
            .O(N__20883),
            .I(N__20705));
    ClkMux I__4883 (
            .O(N__20882),
            .I(N__20705));
    ClkMux I__4882 (
            .O(N__20881),
            .I(N__20705));
    ClkMux I__4881 (
            .O(N__20880),
            .I(N__20705));
    ClkMux I__4880 (
            .O(N__20879),
            .I(N__20705));
    ClkMux I__4879 (
            .O(N__20878),
            .I(N__20705));
    ClkMux I__4878 (
            .O(N__20877),
            .I(N__20705));
    ClkMux I__4877 (
            .O(N__20876),
            .I(N__20705));
    ClkMux I__4876 (
            .O(N__20875),
            .I(N__20705));
    ClkMux I__4875 (
            .O(N__20874),
            .I(N__20705));
    ClkMux I__4874 (
            .O(N__20873),
            .I(N__20705));
    ClkMux I__4873 (
            .O(N__20872),
            .I(N__20705));
    ClkMux I__4872 (
            .O(N__20871),
            .I(N__20705));
    ClkMux I__4871 (
            .O(N__20870),
            .I(N__20705));
    ClkMux I__4870 (
            .O(N__20869),
            .I(N__20705));
    ClkMux I__4869 (
            .O(N__20868),
            .I(N__20705));
    ClkMux I__4868 (
            .O(N__20867),
            .I(N__20705));
    ClkMux I__4867 (
            .O(N__20866),
            .I(N__20705));
    ClkMux I__4866 (
            .O(N__20865),
            .I(N__20705));
    ClkMux I__4865 (
            .O(N__20864),
            .I(N__20705));
    GlobalMux I__4864 (
            .O(N__20705),
            .I(clk_100mhz));
    IoInMux I__4863 (
            .O(N__20702),
            .I(N__20699));
    LocalMux I__4862 (
            .O(N__20699),
            .I(N__20696));
    Odrv12 I__4861 (
            .O(N__20696),
            .I(\delay_measurement_inst.delay_hc_timer.N_253_i ));
    InMux I__4860 (
            .O(N__20693),
            .I(N__20689));
    InMux I__4859 (
            .O(N__20692),
            .I(N__20686));
    LocalMux I__4858 (
            .O(N__20689),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    LocalMux I__4857 (
            .O(N__20686),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    InMux I__4856 (
            .O(N__20681),
            .I(N__20674));
    InMux I__4855 (
            .O(N__20680),
            .I(N__20674));
    InMux I__4854 (
            .O(N__20679),
            .I(N__20671));
    LocalMux I__4853 (
            .O(N__20674),
            .I(N__20668));
    LocalMux I__4852 (
            .O(N__20671),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    Odrv4 I__4851 (
            .O(N__20668),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    CEMux I__4850 (
            .O(N__20663),
            .I(N__20660));
    LocalMux I__4849 (
            .O(N__20660),
            .I(N__20655));
    CEMux I__4848 (
            .O(N__20659),
            .I(N__20652));
    CEMux I__4847 (
            .O(N__20658),
            .I(N__20648));
    Span4Mux_v I__4846 (
            .O(N__20655),
            .I(N__20643));
    LocalMux I__4845 (
            .O(N__20652),
            .I(N__20643));
    CEMux I__4844 (
            .O(N__20651),
            .I(N__20640));
    LocalMux I__4843 (
            .O(N__20648),
            .I(N__20637));
    Span4Mux_h I__4842 (
            .O(N__20643),
            .I(N__20634));
    LocalMux I__4841 (
            .O(N__20640),
            .I(N__20631));
    Span4Mux_v I__4840 (
            .O(N__20637),
            .I(N__20628));
    Span4Mux_h I__4839 (
            .O(N__20634),
            .I(N__20625));
    Sp12to4 I__4838 (
            .O(N__20631),
            .I(N__20622));
    Odrv4 I__4837 (
            .O(N__20628),
            .I(\delay_measurement_inst.delay_hc_timer.N_254_i_g ));
    Odrv4 I__4836 (
            .O(N__20625),
            .I(\delay_measurement_inst.delay_hc_timer.N_254_i_g ));
    Odrv12 I__4835 (
            .O(N__20622),
            .I(\delay_measurement_inst.delay_hc_timer.N_254_i_g ));
    InMux I__4834 (
            .O(N__20615),
            .I(N__20609));
    InMux I__4833 (
            .O(N__20614),
            .I(N__20602));
    InMux I__4832 (
            .O(N__20613),
            .I(N__20602));
    InMux I__4831 (
            .O(N__20612),
            .I(N__20602));
    LocalMux I__4830 (
            .O(N__20609),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__4829 (
            .O(N__20602),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    InMux I__4828 (
            .O(N__20597),
            .I(N__20569));
    InMux I__4827 (
            .O(N__20596),
            .I(N__20569));
    InMux I__4826 (
            .O(N__20595),
            .I(N__20569));
    InMux I__4825 (
            .O(N__20594),
            .I(N__20569));
    InMux I__4824 (
            .O(N__20593),
            .I(N__20560));
    InMux I__4823 (
            .O(N__20592),
            .I(N__20560));
    InMux I__4822 (
            .O(N__20591),
            .I(N__20560));
    InMux I__4821 (
            .O(N__20590),
            .I(N__20560));
    InMux I__4820 (
            .O(N__20589),
            .I(N__20551));
    InMux I__4819 (
            .O(N__20588),
            .I(N__20551));
    InMux I__4818 (
            .O(N__20587),
            .I(N__20551));
    InMux I__4817 (
            .O(N__20586),
            .I(N__20551));
    InMux I__4816 (
            .O(N__20585),
            .I(N__20542));
    InMux I__4815 (
            .O(N__20584),
            .I(N__20542));
    InMux I__4814 (
            .O(N__20583),
            .I(N__20542));
    InMux I__4813 (
            .O(N__20582),
            .I(N__20542));
    InMux I__4812 (
            .O(N__20581),
            .I(N__20533));
    InMux I__4811 (
            .O(N__20580),
            .I(N__20533));
    InMux I__4810 (
            .O(N__20579),
            .I(N__20533));
    InMux I__4809 (
            .O(N__20578),
            .I(N__20533));
    LocalMux I__4808 (
            .O(N__20569),
            .I(N__20518));
    LocalMux I__4807 (
            .O(N__20560),
            .I(N__20518));
    LocalMux I__4806 (
            .O(N__20551),
            .I(N__20511));
    LocalMux I__4805 (
            .O(N__20542),
            .I(N__20511));
    LocalMux I__4804 (
            .O(N__20533),
            .I(N__20511));
    InMux I__4803 (
            .O(N__20532),
            .I(N__20506));
    InMux I__4802 (
            .O(N__20531),
            .I(N__20506));
    InMux I__4801 (
            .O(N__20530),
            .I(N__20497));
    InMux I__4800 (
            .O(N__20529),
            .I(N__20497));
    InMux I__4799 (
            .O(N__20528),
            .I(N__20497));
    InMux I__4798 (
            .O(N__20527),
            .I(N__20497));
    InMux I__4797 (
            .O(N__20526),
            .I(N__20488));
    InMux I__4796 (
            .O(N__20525),
            .I(N__20488));
    InMux I__4795 (
            .O(N__20524),
            .I(N__20488));
    InMux I__4794 (
            .O(N__20523),
            .I(N__20488));
    Span4Mux_v I__4793 (
            .O(N__20518),
            .I(N__20479));
    Span4Mux_v I__4792 (
            .O(N__20511),
            .I(N__20479));
    LocalMux I__4791 (
            .O(N__20506),
            .I(N__20479));
    LocalMux I__4790 (
            .O(N__20497),
            .I(N__20479));
    LocalMux I__4789 (
            .O(N__20488),
            .I(N__20476));
    Span4Mux_h I__4788 (
            .O(N__20479),
            .I(N__20473));
    Odrv12 I__4787 (
            .O(N__20476),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__4786 (
            .O(N__20473),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    CascadeMux I__4785 (
            .O(N__20468),
            .I(N__20458));
    CascadeMux I__4784 (
            .O(N__20467),
            .I(N__20455));
    InMux I__4783 (
            .O(N__20466),
            .I(N__20452));
    InMux I__4782 (
            .O(N__20465),
            .I(N__20447));
    InMux I__4781 (
            .O(N__20464),
            .I(N__20447));
    InMux I__4780 (
            .O(N__20463),
            .I(N__20444));
    InMux I__4779 (
            .O(N__20462),
            .I(N__20441));
    InMux I__4778 (
            .O(N__20461),
            .I(N__20438));
    InMux I__4777 (
            .O(N__20458),
            .I(N__20435));
    InMux I__4776 (
            .O(N__20455),
            .I(N__20432));
    LocalMux I__4775 (
            .O(N__20452),
            .I(N__20429));
    LocalMux I__4774 (
            .O(N__20447),
            .I(N__20426));
    LocalMux I__4773 (
            .O(N__20444),
            .I(N__20402));
    LocalMux I__4772 (
            .O(N__20441),
            .I(N__20386));
    LocalMux I__4771 (
            .O(N__20438),
            .I(N__20363));
    LocalMux I__4770 (
            .O(N__20435),
            .I(N__20357));
    LocalMux I__4769 (
            .O(N__20432),
            .I(N__20347));
    Glb2LocalMux I__4768 (
            .O(N__20429),
            .I(N__20201));
    Glb2LocalMux I__4767 (
            .O(N__20426),
            .I(N__20201));
    SRMux I__4766 (
            .O(N__20425),
            .I(N__20201));
    SRMux I__4765 (
            .O(N__20424),
            .I(N__20201));
    SRMux I__4764 (
            .O(N__20423),
            .I(N__20201));
    SRMux I__4763 (
            .O(N__20422),
            .I(N__20201));
    SRMux I__4762 (
            .O(N__20421),
            .I(N__20201));
    SRMux I__4761 (
            .O(N__20420),
            .I(N__20201));
    SRMux I__4760 (
            .O(N__20419),
            .I(N__20201));
    SRMux I__4759 (
            .O(N__20418),
            .I(N__20201));
    SRMux I__4758 (
            .O(N__20417),
            .I(N__20201));
    SRMux I__4757 (
            .O(N__20416),
            .I(N__20201));
    SRMux I__4756 (
            .O(N__20415),
            .I(N__20201));
    SRMux I__4755 (
            .O(N__20414),
            .I(N__20201));
    SRMux I__4754 (
            .O(N__20413),
            .I(N__20201));
    SRMux I__4753 (
            .O(N__20412),
            .I(N__20201));
    SRMux I__4752 (
            .O(N__20411),
            .I(N__20201));
    SRMux I__4751 (
            .O(N__20410),
            .I(N__20201));
    SRMux I__4750 (
            .O(N__20409),
            .I(N__20201));
    SRMux I__4749 (
            .O(N__20408),
            .I(N__20201));
    SRMux I__4748 (
            .O(N__20407),
            .I(N__20201));
    SRMux I__4747 (
            .O(N__20406),
            .I(N__20201));
    SRMux I__4746 (
            .O(N__20405),
            .I(N__20201));
    Glb2LocalMux I__4745 (
            .O(N__20402),
            .I(N__20201));
    SRMux I__4744 (
            .O(N__20401),
            .I(N__20201));
    SRMux I__4743 (
            .O(N__20400),
            .I(N__20201));
    SRMux I__4742 (
            .O(N__20399),
            .I(N__20201));
    SRMux I__4741 (
            .O(N__20398),
            .I(N__20201));
    SRMux I__4740 (
            .O(N__20397),
            .I(N__20201));
    SRMux I__4739 (
            .O(N__20396),
            .I(N__20201));
    SRMux I__4738 (
            .O(N__20395),
            .I(N__20201));
    SRMux I__4737 (
            .O(N__20394),
            .I(N__20201));
    SRMux I__4736 (
            .O(N__20393),
            .I(N__20201));
    SRMux I__4735 (
            .O(N__20392),
            .I(N__20201));
    SRMux I__4734 (
            .O(N__20391),
            .I(N__20201));
    SRMux I__4733 (
            .O(N__20390),
            .I(N__20201));
    SRMux I__4732 (
            .O(N__20389),
            .I(N__20201));
    Glb2LocalMux I__4731 (
            .O(N__20386),
            .I(N__20201));
    SRMux I__4730 (
            .O(N__20385),
            .I(N__20201));
    SRMux I__4729 (
            .O(N__20384),
            .I(N__20201));
    SRMux I__4728 (
            .O(N__20383),
            .I(N__20201));
    SRMux I__4727 (
            .O(N__20382),
            .I(N__20201));
    SRMux I__4726 (
            .O(N__20381),
            .I(N__20201));
    SRMux I__4725 (
            .O(N__20380),
            .I(N__20201));
    SRMux I__4724 (
            .O(N__20379),
            .I(N__20201));
    SRMux I__4723 (
            .O(N__20378),
            .I(N__20201));
    SRMux I__4722 (
            .O(N__20377),
            .I(N__20201));
    SRMux I__4721 (
            .O(N__20376),
            .I(N__20201));
    SRMux I__4720 (
            .O(N__20375),
            .I(N__20201));
    SRMux I__4719 (
            .O(N__20374),
            .I(N__20201));
    SRMux I__4718 (
            .O(N__20373),
            .I(N__20201));
    SRMux I__4717 (
            .O(N__20372),
            .I(N__20201));
    SRMux I__4716 (
            .O(N__20371),
            .I(N__20201));
    SRMux I__4715 (
            .O(N__20370),
            .I(N__20201));
    SRMux I__4714 (
            .O(N__20369),
            .I(N__20201));
    SRMux I__4713 (
            .O(N__20368),
            .I(N__20201));
    SRMux I__4712 (
            .O(N__20367),
            .I(N__20201));
    SRMux I__4711 (
            .O(N__20366),
            .I(N__20201));
    Glb2LocalMux I__4710 (
            .O(N__20363),
            .I(N__20201));
    SRMux I__4709 (
            .O(N__20362),
            .I(N__20201));
    SRMux I__4708 (
            .O(N__20361),
            .I(N__20201));
    SRMux I__4707 (
            .O(N__20360),
            .I(N__20201));
    Glb2LocalMux I__4706 (
            .O(N__20357),
            .I(N__20201));
    SRMux I__4705 (
            .O(N__20356),
            .I(N__20201));
    SRMux I__4704 (
            .O(N__20355),
            .I(N__20201));
    SRMux I__4703 (
            .O(N__20354),
            .I(N__20201));
    SRMux I__4702 (
            .O(N__20353),
            .I(N__20201));
    SRMux I__4701 (
            .O(N__20352),
            .I(N__20201));
    SRMux I__4700 (
            .O(N__20351),
            .I(N__20201));
    SRMux I__4699 (
            .O(N__20350),
            .I(N__20201));
    Glb2LocalMux I__4698 (
            .O(N__20347),
            .I(N__20201));
    SRMux I__4697 (
            .O(N__20346),
            .I(N__20201));
    GlobalMux I__4696 (
            .O(N__20201),
            .I(N__20198));
    gio2CtrlBuf I__4695 (
            .O(N__20198),
            .I(red_c_g));
    CEMux I__4694 (
            .O(N__20195),
            .I(N__20192));
    LocalMux I__4693 (
            .O(N__20192),
            .I(N__20185));
    CEMux I__4692 (
            .O(N__20191),
            .I(N__20182));
    CEMux I__4691 (
            .O(N__20190),
            .I(N__20178));
    CEMux I__4690 (
            .O(N__20189),
            .I(N__20175));
    CEMux I__4689 (
            .O(N__20188),
            .I(N__20172));
    Span4Mux_v I__4688 (
            .O(N__20185),
            .I(N__20168));
    LocalMux I__4687 (
            .O(N__20182),
            .I(N__20165));
    IoInMux I__4686 (
            .O(N__20181),
            .I(N__20162));
    LocalMux I__4685 (
            .O(N__20178),
            .I(N__20159));
    LocalMux I__4684 (
            .O(N__20175),
            .I(N__20156));
    LocalMux I__4683 (
            .O(N__20172),
            .I(N__20153));
    CEMux I__4682 (
            .O(N__20171),
            .I(N__20150));
    Span4Mux_v I__4681 (
            .O(N__20168),
            .I(N__20147));
    Span4Mux_h I__4680 (
            .O(N__20165),
            .I(N__20144));
    LocalMux I__4679 (
            .O(N__20162),
            .I(N__20141));
    Span4Mux_h I__4678 (
            .O(N__20159),
            .I(N__20136));
    Span4Mux_h I__4677 (
            .O(N__20156),
            .I(N__20136));
    Span4Mux_v I__4676 (
            .O(N__20153),
            .I(N__20131));
    LocalMux I__4675 (
            .O(N__20150),
            .I(N__20131));
    Span4Mux_h I__4674 (
            .O(N__20147),
            .I(N__20128));
    Span4Mux_h I__4673 (
            .O(N__20144),
            .I(N__20125));
    IoSpan4Mux I__4672 (
            .O(N__20141),
            .I(N__20122));
    Span4Mux_h I__4671 (
            .O(N__20136),
            .I(N__20117));
    Span4Mux_v I__4670 (
            .O(N__20131),
            .I(N__20117));
    Span4Mux_h I__4669 (
            .O(N__20128),
            .I(N__20114));
    Span4Mux_h I__4668 (
            .O(N__20125),
            .I(N__20107));
    Span4Mux_s2_v I__4667 (
            .O(N__20122),
            .I(N__20107));
    Span4Mux_v I__4666 (
            .O(N__20117),
            .I(N__20107));
    Odrv4 I__4665 (
            .O(N__20114),
            .I(red_c_i));
    Odrv4 I__4664 (
            .O(N__20107),
            .I(red_c_i));
    InMux I__4663 (
            .O(N__20102),
            .I(N__20098));
    InMux I__4662 (
            .O(N__20101),
            .I(N__20095));
    LocalMux I__4661 (
            .O(N__20098),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    LocalMux I__4660 (
            .O(N__20095),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    InMux I__4659 (
            .O(N__20090),
            .I(N__20085));
    InMux I__4658 (
            .O(N__20089),
            .I(N__20082));
    InMux I__4657 (
            .O(N__20088),
            .I(N__20079));
    LocalMux I__4656 (
            .O(N__20085),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    LocalMux I__4655 (
            .O(N__20082),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    LocalMux I__4654 (
            .O(N__20079),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    InMux I__4653 (
            .O(N__20072),
            .I(N__20066));
    InMux I__4652 (
            .O(N__20071),
            .I(N__20063));
    InMux I__4651 (
            .O(N__20070),
            .I(N__20060));
    InMux I__4650 (
            .O(N__20069),
            .I(N__20057));
    LocalMux I__4649 (
            .O(N__20066),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__4648 (
            .O(N__20063),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__4647 (
            .O(N__20060),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__4646 (
            .O(N__20057),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    IoInMux I__4645 (
            .O(N__20048),
            .I(N__20045));
    LocalMux I__4644 (
            .O(N__20045),
            .I(N__20042));
    Span12Mux_s5_v I__4643 (
            .O(N__20042),
            .I(N__20039));
    Odrv12 I__4642 (
            .O(N__20039),
            .I(\delay_measurement_inst.delay_tr_timer.N_256_i ));
    InMux I__4641 (
            .O(N__20036),
            .I(N__20033));
    LocalMux I__4640 (
            .O(N__20033),
            .I(N__20030));
    Span4Mux_v I__4639 (
            .O(N__20030),
            .I(N__20027));
    Sp12to4 I__4638 (
            .O(N__20027),
            .I(N__20024));
    Span12Mux_s10_h I__4637 (
            .O(N__20024),
            .I(N__20021));
    Odrv12 I__4636 (
            .O(N__20021),
            .I(delay_tr_input_c));
    InMux I__4635 (
            .O(N__20018),
            .I(N__20015));
    LocalMux I__4634 (
            .O(N__20015),
            .I(delay_tr_d1));
    InMux I__4633 (
            .O(N__20012),
            .I(N__20006));
    InMux I__4632 (
            .O(N__20011),
            .I(N__20003));
    InMux I__4631 (
            .O(N__20010),
            .I(N__19998));
    InMux I__4630 (
            .O(N__20009),
            .I(N__19998));
    LocalMux I__4629 (
            .O(N__20006),
            .I(delay_tr_d2));
    LocalMux I__4628 (
            .O(N__20003),
            .I(delay_tr_d2));
    LocalMux I__4627 (
            .O(N__19998),
            .I(delay_tr_d2));
    InMux I__4626 (
            .O(N__19991),
            .I(N__19986));
    InMux I__4625 (
            .O(N__19990),
            .I(N__19983));
    InMux I__4624 (
            .O(N__19989),
            .I(N__19980));
    LocalMux I__4623 (
            .O(N__19986),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    LocalMux I__4622 (
            .O(N__19983),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    LocalMux I__4621 (
            .O(N__19980),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    InMux I__4620 (
            .O(N__19973),
            .I(N__19968));
    InMux I__4619 (
            .O(N__19972),
            .I(N__19965));
    InMux I__4618 (
            .O(N__19971),
            .I(N__19962));
    LocalMux I__4617 (
            .O(N__19968),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    LocalMux I__4616 (
            .O(N__19965),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    LocalMux I__4615 (
            .O(N__19962),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    InMux I__4614 (
            .O(N__19955),
            .I(N__19952));
    LocalMux I__4613 (
            .O(N__19952),
            .I(N__19949));
    Span12Mux_h I__4612 (
            .O(N__19949),
            .I(N__19946));
    Span12Mux_v I__4611 (
            .O(N__19946),
            .I(N__19943));
    Odrv12 I__4610 (
            .O(N__19943),
            .I(delay_hc_input_c));
    InMux I__4609 (
            .O(N__19940),
            .I(N__19937));
    LocalMux I__4608 (
            .O(N__19937),
            .I(delay_hc_d1));
    IoInMux I__4607 (
            .O(N__19934),
            .I(N__19931));
    LocalMux I__4606 (
            .O(N__19931),
            .I(N__19928));
    Span12Mux_s4_v I__4605 (
            .O(N__19928),
            .I(N__19925));
    Span12Mux_v I__4604 (
            .O(N__19925),
            .I(N__19922));
    Odrv12 I__4603 (
            .O(N__19922),
            .I(\delay_measurement_inst.delay_tr_timer.N_255_i ));
    InMux I__4602 (
            .O(N__19919),
            .I(N__19916));
    LocalMux I__4601 (
            .O(N__19916),
            .I(N__19911));
    CascadeMux I__4600 (
            .O(N__19915),
            .I(N__19907));
    CascadeMux I__4599 (
            .O(N__19914),
            .I(N__19904));
    Span4Mux_h I__4598 (
            .O(N__19911),
            .I(N__19901));
    InMux I__4597 (
            .O(N__19910),
            .I(N__19898));
    InMux I__4596 (
            .O(N__19907),
            .I(N__19893));
    InMux I__4595 (
            .O(N__19904),
            .I(N__19893));
    Span4Mux_v I__4594 (
            .O(N__19901),
            .I(N__19888));
    LocalMux I__4593 (
            .O(N__19898),
            .I(N__19888));
    LocalMux I__4592 (
            .O(N__19893),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__4591 (
            .O(N__19888),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    IoInMux I__4590 (
            .O(N__19883),
            .I(N__19880));
    LocalMux I__4589 (
            .O(N__19880),
            .I(N__19877));
    Span4Mux_s3_v I__4588 (
            .O(N__19877),
            .I(N__19874));
    Span4Mux_v I__4587 (
            .O(N__19874),
            .I(N__19871));
    Span4Mux_v I__4586 (
            .O(N__19871),
            .I(N__19868));
    Odrv4 I__4585 (
            .O(N__19868),
            .I(s2_phy_c));
    InMux I__4584 (
            .O(N__19865),
            .I(N__19862));
    LocalMux I__4583 (
            .O(N__19862),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__4582 (
            .O(N__19859),
            .I(N__19856));
    LocalMux I__4581 (
            .O(N__19856),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    CascadeMux I__4580 (
            .O(N__19853),
            .I(N__19850));
    InMux I__4579 (
            .O(N__19850),
            .I(N__19847));
    LocalMux I__4578 (
            .O(N__19847),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    InMux I__4577 (
            .O(N__19844),
            .I(N__19841));
    LocalMux I__4576 (
            .O(N__19841),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    InMux I__4575 (
            .O(N__19838),
            .I(N__19835));
    LocalMux I__4574 (
            .O(N__19835),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    CascadeMux I__4573 (
            .O(N__19832),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_7_19_cascade_ ));
    InMux I__4572 (
            .O(N__19829),
            .I(N__19810));
    InMux I__4571 (
            .O(N__19828),
            .I(N__19810));
    InMux I__4570 (
            .O(N__19827),
            .I(N__19810));
    InMux I__4569 (
            .O(N__19826),
            .I(N__19810));
    InMux I__4568 (
            .O(N__19825),
            .I(N__19810));
    InMux I__4567 (
            .O(N__19824),
            .I(N__19801));
    InMux I__4566 (
            .O(N__19823),
            .I(N__19801));
    InMux I__4565 (
            .O(N__19822),
            .I(N__19801));
    InMux I__4564 (
            .O(N__19821),
            .I(N__19801));
    LocalMux I__4563 (
            .O(N__19810),
            .I(N__19798));
    LocalMux I__4562 (
            .O(N__19801),
            .I(N__19795));
    Odrv12 I__4561 (
            .O(N__19798),
            .I(\delay_measurement_inst.N_276 ));
    Odrv4 I__4560 (
            .O(N__19795),
            .I(\delay_measurement_inst.N_276 ));
    InMux I__4559 (
            .O(N__19790),
            .I(N__19787));
    LocalMux I__4558 (
            .O(N__19787),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    InMux I__4557 (
            .O(N__19784),
            .I(N__19781));
    LocalMux I__4556 (
            .O(N__19781),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    CascadeMux I__4555 (
            .O(N__19778),
            .I(N__19775));
    InMux I__4554 (
            .O(N__19775),
            .I(N__19772));
    LocalMux I__4553 (
            .O(N__19772),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    InMux I__4552 (
            .O(N__19769),
            .I(N__19766));
    LocalMux I__4551 (
            .O(N__19766),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    InMux I__4550 (
            .O(N__19763),
            .I(N__19760));
    LocalMux I__4549 (
            .O(N__19760),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_6_19 ));
    InMux I__4548 (
            .O(N__19757),
            .I(N__19754));
    LocalMux I__4547 (
            .O(N__19754),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30 ));
    InMux I__4546 (
            .O(N__19751),
            .I(N__19748));
    LocalMux I__4545 (
            .O(N__19748),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    InMux I__4544 (
            .O(N__19745),
            .I(N__19742));
    LocalMux I__4543 (
            .O(N__19742),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_0_19 ));
    InMux I__4542 (
            .O(N__19739),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__4541 (
            .O(N__19736),
            .I(N__19731));
    CascadeMux I__4540 (
            .O(N__19735),
            .I(N__19728));
    InMux I__4539 (
            .O(N__19734),
            .I(N__19725));
    InMux I__4538 (
            .O(N__19731),
            .I(N__19720));
    InMux I__4537 (
            .O(N__19728),
            .I(N__19720));
    LocalMux I__4536 (
            .O(N__19725),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    LocalMux I__4535 (
            .O(N__19720),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__4534 (
            .O(N__19715),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__4533 (
            .O(N__19712),
            .I(N__19707));
    CascadeMux I__4532 (
            .O(N__19711),
            .I(N__19704));
    InMux I__4531 (
            .O(N__19710),
            .I(N__19701));
    InMux I__4530 (
            .O(N__19707),
            .I(N__19696));
    InMux I__4529 (
            .O(N__19704),
            .I(N__19696));
    LocalMux I__4528 (
            .O(N__19701),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    LocalMux I__4527 (
            .O(N__19696),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__4526 (
            .O(N__19691),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__4525 (
            .O(N__19688),
            .I(N__19683));
    InMux I__4524 (
            .O(N__19687),
            .I(N__19680));
    InMux I__4523 (
            .O(N__19686),
            .I(N__19677));
    LocalMux I__4522 (
            .O(N__19683),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    LocalMux I__4521 (
            .O(N__19680),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    LocalMux I__4520 (
            .O(N__19677),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__4519 (
            .O(N__19670),
            .I(bfn_10_24_0_));
    InMux I__4518 (
            .O(N__19667),
            .I(N__19662));
    InMux I__4517 (
            .O(N__19666),
            .I(N__19659));
    InMux I__4516 (
            .O(N__19665),
            .I(N__19656));
    LocalMux I__4515 (
            .O(N__19662),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    LocalMux I__4514 (
            .O(N__19659),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    LocalMux I__4513 (
            .O(N__19656),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__4512 (
            .O(N__19649),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__4511 (
            .O(N__19646),
            .I(N__19642));
    InMux I__4510 (
            .O(N__19645),
            .I(N__19639));
    LocalMux I__4509 (
            .O(N__19642),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    LocalMux I__4508 (
            .O(N__19639),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    CascadeMux I__4507 (
            .O(N__19634),
            .I(N__19629));
    CascadeMux I__4506 (
            .O(N__19633),
            .I(N__19626));
    InMux I__4505 (
            .O(N__19632),
            .I(N__19623));
    InMux I__4504 (
            .O(N__19629),
            .I(N__19618));
    InMux I__4503 (
            .O(N__19626),
            .I(N__19618));
    LocalMux I__4502 (
            .O(N__19623),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    LocalMux I__4501 (
            .O(N__19618),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    InMux I__4500 (
            .O(N__19613),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__4499 (
            .O(N__19610),
            .I(N__19606));
    InMux I__4498 (
            .O(N__19609),
            .I(N__19603));
    LocalMux I__4497 (
            .O(N__19606),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    LocalMux I__4496 (
            .O(N__19603),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    CascadeMux I__4495 (
            .O(N__19598),
            .I(N__19593));
    CascadeMux I__4494 (
            .O(N__19597),
            .I(N__19590));
    InMux I__4493 (
            .O(N__19596),
            .I(N__19587));
    InMux I__4492 (
            .O(N__19593),
            .I(N__19582));
    InMux I__4491 (
            .O(N__19590),
            .I(N__19582));
    LocalMux I__4490 (
            .O(N__19587),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    LocalMux I__4489 (
            .O(N__19582),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__4488 (
            .O(N__19577),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__4487 (
            .O(N__19574),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    CascadeMux I__4486 (
            .O(N__19571),
            .I(N__19563));
    CascadeMux I__4485 (
            .O(N__19570),
            .I(N__19554));
    InMux I__4484 (
            .O(N__19569),
            .I(N__19546));
    InMux I__4483 (
            .O(N__19568),
            .I(N__19546));
    InMux I__4482 (
            .O(N__19567),
            .I(N__19546));
    InMux I__4481 (
            .O(N__19566),
            .I(N__19543));
    InMux I__4480 (
            .O(N__19563),
            .I(N__19532));
    InMux I__4479 (
            .O(N__19562),
            .I(N__19532));
    InMux I__4478 (
            .O(N__19561),
            .I(N__19532));
    InMux I__4477 (
            .O(N__19560),
            .I(N__19532));
    InMux I__4476 (
            .O(N__19559),
            .I(N__19532));
    InMux I__4475 (
            .O(N__19558),
            .I(N__19527));
    InMux I__4474 (
            .O(N__19557),
            .I(N__19527));
    InMux I__4473 (
            .O(N__19554),
            .I(N__19524));
    InMux I__4472 (
            .O(N__19553),
            .I(N__19521));
    LocalMux I__4471 (
            .O(N__19546),
            .I(N__19516));
    LocalMux I__4470 (
            .O(N__19543),
            .I(N__19516));
    LocalMux I__4469 (
            .O(N__19532),
            .I(N__19509));
    LocalMux I__4468 (
            .O(N__19527),
            .I(N__19509));
    LocalMux I__4467 (
            .O(N__19524),
            .I(N__19509));
    LocalMux I__4466 (
            .O(N__19521),
            .I(N__19504));
    Span4Mux_v I__4465 (
            .O(N__19516),
            .I(N__19504));
    Span4Mux_h I__4464 (
            .O(N__19509),
            .I(N__19501));
    Odrv4 I__4463 (
            .O(N__19504),
            .I(\delay_measurement_inst.elapsed_time_hc_31 ));
    Odrv4 I__4462 (
            .O(N__19501),
            .I(\delay_measurement_inst.elapsed_time_hc_31 ));
    CEMux I__4461 (
            .O(N__19496),
            .I(N__19481));
    CEMux I__4460 (
            .O(N__19495),
            .I(N__19481));
    CEMux I__4459 (
            .O(N__19494),
            .I(N__19481));
    CEMux I__4458 (
            .O(N__19493),
            .I(N__19481));
    CEMux I__4457 (
            .O(N__19492),
            .I(N__19481));
    GlobalMux I__4456 (
            .O(N__19481),
            .I(N__19478));
    gio2CtrlBuf I__4455 (
            .O(N__19478),
            .I(\delay_measurement_inst.delay_hc_timer.N_253_i_g ));
    InMux I__4454 (
            .O(N__19475),
            .I(N__19470));
    InMux I__4453 (
            .O(N__19474),
            .I(N__19465));
    InMux I__4452 (
            .O(N__19473),
            .I(N__19465));
    LocalMux I__4451 (
            .O(N__19470),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    LocalMux I__4450 (
            .O(N__19465),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__4449 (
            .O(N__19460),
            .I(N__19455));
    InMux I__4448 (
            .O(N__19459),
            .I(N__19452));
    InMux I__4447 (
            .O(N__19458),
            .I(N__19449));
    LocalMux I__4446 (
            .O(N__19455),
            .I(N__19446));
    LocalMux I__4445 (
            .O(N__19452),
            .I(N__19441));
    LocalMux I__4444 (
            .O(N__19449),
            .I(N__19441));
    Span4Mux_v I__4443 (
            .O(N__19446),
            .I(N__19436));
    Span4Mux_v I__4442 (
            .O(N__19441),
            .I(N__19436));
    Odrv4 I__4441 (
            .O(N__19436),
            .I(\delay_measurement_inst.elapsed_time_hc_16 ));
    InMux I__4440 (
            .O(N__19433),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__4439 (
            .O(N__19430),
            .I(N__19425));
    CascadeMux I__4438 (
            .O(N__19429),
            .I(N__19422));
    InMux I__4437 (
            .O(N__19428),
            .I(N__19419));
    InMux I__4436 (
            .O(N__19425),
            .I(N__19414));
    InMux I__4435 (
            .O(N__19422),
            .I(N__19414));
    LocalMux I__4434 (
            .O(N__19419),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    LocalMux I__4433 (
            .O(N__19414),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    CascadeMux I__4432 (
            .O(N__19409),
            .I(N__19405));
    InMux I__4431 (
            .O(N__19408),
            .I(N__19401));
    InMux I__4430 (
            .O(N__19405),
            .I(N__19398));
    InMux I__4429 (
            .O(N__19404),
            .I(N__19395));
    LocalMux I__4428 (
            .O(N__19401),
            .I(N__19390));
    LocalMux I__4427 (
            .O(N__19398),
            .I(N__19390));
    LocalMux I__4426 (
            .O(N__19395),
            .I(N__19387));
    Span4Mux_h I__4425 (
            .O(N__19390),
            .I(N__19384));
    Odrv4 I__4424 (
            .O(N__19387),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    Odrv4 I__4423 (
            .O(N__19384),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    InMux I__4422 (
            .O(N__19379),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__4421 (
            .O(N__19376),
            .I(N__19371));
    CascadeMux I__4420 (
            .O(N__19375),
            .I(N__19368));
    InMux I__4419 (
            .O(N__19374),
            .I(N__19365));
    InMux I__4418 (
            .O(N__19371),
            .I(N__19360));
    InMux I__4417 (
            .O(N__19368),
            .I(N__19360));
    LocalMux I__4416 (
            .O(N__19365),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    LocalMux I__4415 (
            .O(N__19360),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__4414 (
            .O(N__19355),
            .I(N__19351));
    InMux I__4413 (
            .O(N__19354),
            .I(N__19348));
    LocalMux I__4412 (
            .O(N__19351),
            .I(N__19342));
    LocalMux I__4411 (
            .O(N__19348),
            .I(N__19342));
    InMux I__4410 (
            .O(N__19347),
            .I(N__19339));
    Span4Mux_v I__4409 (
            .O(N__19342),
            .I(N__19334));
    LocalMux I__4408 (
            .O(N__19339),
            .I(N__19334));
    Odrv4 I__4407 (
            .O(N__19334),
            .I(\delay_measurement_inst.elapsed_time_hc_18 ));
    InMux I__4406 (
            .O(N__19331),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__4405 (
            .O(N__19328),
            .I(N__19323));
    InMux I__4404 (
            .O(N__19327),
            .I(N__19320));
    InMux I__4403 (
            .O(N__19326),
            .I(N__19317));
    LocalMux I__4402 (
            .O(N__19323),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    LocalMux I__4401 (
            .O(N__19320),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    LocalMux I__4400 (
            .O(N__19317),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    CascadeMux I__4399 (
            .O(N__19310),
            .I(N__19305));
    InMux I__4398 (
            .O(N__19309),
            .I(N__19302));
    InMux I__4397 (
            .O(N__19308),
            .I(N__19299));
    InMux I__4396 (
            .O(N__19305),
            .I(N__19296));
    LocalMux I__4395 (
            .O(N__19302),
            .I(N__19293));
    LocalMux I__4394 (
            .O(N__19299),
            .I(N__19288));
    LocalMux I__4393 (
            .O(N__19296),
            .I(N__19288));
    Span4Mux_h I__4392 (
            .O(N__19293),
            .I(N__19283));
    Span4Mux_v I__4391 (
            .O(N__19288),
            .I(N__19283));
    Odrv4 I__4390 (
            .O(N__19283),
            .I(\delay_measurement_inst.elapsed_time_hc_19 ));
    InMux I__4389 (
            .O(N__19280),
            .I(bfn_10_23_0_));
    InMux I__4388 (
            .O(N__19277),
            .I(N__19272));
    InMux I__4387 (
            .O(N__19276),
            .I(N__19269));
    InMux I__4386 (
            .O(N__19275),
            .I(N__19266));
    LocalMux I__4385 (
            .O(N__19272),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    LocalMux I__4384 (
            .O(N__19269),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    LocalMux I__4383 (
            .O(N__19266),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__4382 (
            .O(N__19259),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__4381 (
            .O(N__19256),
            .I(N__19251));
    CascadeMux I__4380 (
            .O(N__19255),
            .I(N__19248));
    InMux I__4379 (
            .O(N__19254),
            .I(N__19245));
    InMux I__4378 (
            .O(N__19251),
            .I(N__19240));
    InMux I__4377 (
            .O(N__19248),
            .I(N__19240));
    LocalMux I__4376 (
            .O(N__19245),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    LocalMux I__4375 (
            .O(N__19240),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__4374 (
            .O(N__19235),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__4373 (
            .O(N__19232),
            .I(N__19227));
    CascadeMux I__4372 (
            .O(N__19231),
            .I(N__19224));
    InMux I__4371 (
            .O(N__19230),
            .I(N__19221));
    InMux I__4370 (
            .O(N__19227),
            .I(N__19216));
    InMux I__4369 (
            .O(N__19224),
            .I(N__19216));
    LocalMux I__4368 (
            .O(N__19221),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    LocalMux I__4367 (
            .O(N__19216),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__4366 (
            .O(N__19211),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__4365 (
            .O(N__19208),
            .I(N__19203));
    InMux I__4364 (
            .O(N__19207),
            .I(N__19198));
    InMux I__4363 (
            .O(N__19206),
            .I(N__19198));
    LocalMux I__4362 (
            .O(N__19203),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    LocalMux I__4361 (
            .O(N__19198),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__4360 (
            .O(N__19193),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__4359 (
            .O(N__19190),
            .I(N__19185));
    InMux I__4358 (
            .O(N__19189),
            .I(N__19180));
    InMux I__4357 (
            .O(N__19188),
            .I(N__19180));
    LocalMux I__4356 (
            .O(N__19185),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    LocalMux I__4355 (
            .O(N__19180),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    CascadeMux I__4354 (
            .O(N__19175),
            .I(N__19170));
    CascadeMux I__4353 (
            .O(N__19174),
            .I(N__19167));
    InMux I__4352 (
            .O(N__19173),
            .I(N__19164));
    InMux I__4351 (
            .O(N__19170),
            .I(N__19159));
    InMux I__4350 (
            .O(N__19167),
            .I(N__19159));
    LocalMux I__4349 (
            .O(N__19164),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    LocalMux I__4348 (
            .O(N__19159),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    CascadeMux I__4347 (
            .O(N__19154),
            .I(N__19150));
    CascadeMux I__4346 (
            .O(N__19153),
            .I(N__19147));
    InMux I__4345 (
            .O(N__19150),
            .I(N__19141));
    InMux I__4344 (
            .O(N__19147),
            .I(N__19136));
    InMux I__4343 (
            .O(N__19146),
            .I(N__19136));
    InMux I__4342 (
            .O(N__19145),
            .I(N__19131));
    InMux I__4341 (
            .O(N__19144),
            .I(N__19131));
    LocalMux I__4340 (
            .O(N__19141),
            .I(N__19128));
    LocalMux I__4339 (
            .O(N__19136),
            .I(N__19125));
    LocalMux I__4338 (
            .O(N__19131),
            .I(N__19122));
    Span4Mux_h I__4337 (
            .O(N__19128),
            .I(N__19117));
    Span4Mux_h I__4336 (
            .O(N__19125),
            .I(N__19117));
    Span4Mux_h I__4335 (
            .O(N__19122),
            .I(N__19114));
    Odrv4 I__4334 (
            .O(N__19117),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    Odrv4 I__4333 (
            .O(N__19114),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    InMux I__4332 (
            .O(N__19109),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__4331 (
            .O(N__19106),
            .I(N__19101));
    CascadeMux I__4330 (
            .O(N__19105),
            .I(N__19098));
    InMux I__4329 (
            .O(N__19104),
            .I(N__19095));
    InMux I__4328 (
            .O(N__19101),
            .I(N__19090));
    InMux I__4327 (
            .O(N__19098),
            .I(N__19090));
    LocalMux I__4326 (
            .O(N__19095),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    LocalMux I__4325 (
            .O(N__19090),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__4324 (
            .O(N__19085),
            .I(N__19081));
    InMux I__4323 (
            .O(N__19084),
            .I(N__19078));
    LocalMux I__4322 (
            .O(N__19081),
            .I(N__19073));
    LocalMux I__4321 (
            .O(N__19078),
            .I(N__19073));
    Span4Mux_h I__4320 (
            .O(N__19073),
            .I(N__19070));
    Odrv4 I__4319 (
            .O(N__19070),
            .I(\delay_measurement_inst.elapsed_time_hc_10 ));
    InMux I__4318 (
            .O(N__19067),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__4317 (
            .O(N__19064),
            .I(N__19059));
    InMux I__4316 (
            .O(N__19063),
            .I(N__19056));
    InMux I__4315 (
            .O(N__19062),
            .I(N__19053));
    LocalMux I__4314 (
            .O(N__19059),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    LocalMux I__4313 (
            .O(N__19056),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    LocalMux I__4312 (
            .O(N__19053),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__4311 (
            .O(N__19046),
            .I(N__19042));
    InMux I__4310 (
            .O(N__19045),
            .I(N__19039));
    LocalMux I__4309 (
            .O(N__19042),
            .I(N__19036));
    LocalMux I__4308 (
            .O(N__19039),
            .I(N__19033));
    Odrv12 I__4307 (
            .O(N__19036),
            .I(\delay_measurement_inst.elapsed_time_hc_11 ));
    Odrv4 I__4306 (
            .O(N__19033),
            .I(\delay_measurement_inst.elapsed_time_hc_11 ));
    InMux I__4305 (
            .O(N__19028),
            .I(bfn_10_22_0_));
    InMux I__4304 (
            .O(N__19025),
            .I(N__19020));
    InMux I__4303 (
            .O(N__19024),
            .I(N__19017));
    InMux I__4302 (
            .O(N__19023),
            .I(N__19014));
    LocalMux I__4301 (
            .O(N__19020),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    LocalMux I__4300 (
            .O(N__19017),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    LocalMux I__4299 (
            .O(N__19014),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__4298 (
            .O(N__19007),
            .I(N__19004));
    LocalMux I__4297 (
            .O(N__19004),
            .I(N__19000));
    InMux I__4296 (
            .O(N__19003),
            .I(N__18997));
    Span4Mux_h I__4295 (
            .O(N__19000),
            .I(N__18992));
    LocalMux I__4294 (
            .O(N__18997),
            .I(N__18992));
    Odrv4 I__4293 (
            .O(N__18992),
            .I(\delay_measurement_inst.elapsed_time_hc_12 ));
    InMux I__4292 (
            .O(N__18989),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__4291 (
            .O(N__18986),
            .I(N__18981));
    CascadeMux I__4290 (
            .O(N__18985),
            .I(N__18978));
    InMux I__4289 (
            .O(N__18984),
            .I(N__18975));
    InMux I__4288 (
            .O(N__18981),
            .I(N__18970));
    InMux I__4287 (
            .O(N__18978),
            .I(N__18970));
    LocalMux I__4286 (
            .O(N__18975),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    LocalMux I__4285 (
            .O(N__18970),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__4284 (
            .O(N__18965),
            .I(N__18961));
    CascadeMux I__4283 (
            .O(N__18964),
            .I(N__18958));
    LocalMux I__4282 (
            .O(N__18961),
            .I(N__18955));
    InMux I__4281 (
            .O(N__18958),
            .I(N__18952));
    Span4Mux_v I__4280 (
            .O(N__18955),
            .I(N__18949));
    LocalMux I__4279 (
            .O(N__18952),
            .I(N__18946));
    Odrv4 I__4278 (
            .O(N__18949),
            .I(\delay_measurement_inst.elapsed_time_hc_13 ));
    Odrv4 I__4277 (
            .O(N__18946),
            .I(\delay_measurement_inst.elapsed_time_hc_13 ));
    InMux I__4276 (
            .O(N__18941),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__4275 (
            .O(N__18938),
            .I(N__18933));
    CascadeMux I__4274 (
            .O(N__18937),
            .I(N__18930));
    InMux I__4273 (
            .O(N__18936),
            .I(N__18927));
    InMux I__4272 (
            .O(N__18933),
            .I(N__18922));
    InMux I__4271 (
            .O(N__18930),
            .I(N__18922));
    LocalMux I__4270 (
            .O(N__18927),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    LocalMux I__4269 (
            .O(N__18922),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    CascadeMux I__4268 (
            .O(N__18917),
            .I(N__18912));
    InMux I__4267 (
            .O(N__18916),
            .I(N__18907));
    InMux I__4266 (
            .O(N__18915),
            .I(N__18902));
    InMux I__4265 (
            .O(N__18912),
            .I(N__18902));
    InMux I__4264 (
            .O(N__18911),
            .I(N__18899));
    InMux I__4263 (
            .O(N__18910),
            .I(N__18896));
    LocalMux I__4262 (
            .O(N__18907),
            .I(N__18893));
    LocalMux I__4261 (
            .O(N__18902),
            .I(N__18890));
    LocalMux I__4260 (
            .O(N__18899),
            .I(N__18885));
    LocalMux I__4259 (
            .O(N__18896),
            .I(N__18885));
    Span4Mux_h I__4258 (
            .O(N__18893),
            .I(N__18882));
    Span4Mux_v I__4257 (
            .O(N__18890),
            .I(N__18877));
    Span4Mux_h I__4256 (
            .O(N__18885),
            .I(N__18877));
    Odrv4 I__4255 (
            .O(N__18882),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    Odrv4 I__4254 (
            .O(N__18877),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    InMux I__4253 (
            .O(N__18872),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__4252 (
            .O(N__18869),
            .I(N__18864));
    InMux I__4251 (
            .O(N__18868),
            .I(N__18859));
    InMux I__4250 (
            .O(N__18867),
            .I(N__18859));
    LocalMux I__4249 (
            .O(N__18864),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    LocalMux I__4248 (
            .O(N__18859),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__4247 (
            .O(N__18854),
            .I(N__18846));
    InMux I__4246 (
            .O(N__18853),
            .I(N__18846));
    InMux I__4245 (
            .O(N__18852),
            .I(N__18840));
    InMux I__4244 (
            .O(N__18851),
            .I(N__18840));
    LocalMux I__4243 (
            .O(N__18846),
            .I(N__18834));
    InMux I__4242 (
            .O(N__18845),
            .I(N__18831));
    LocalMux I__4241 (
            .O(N__18840),
            .I(N__18828));
    InMux I__4240 (
            .O(N__18839),
            .I(N__18825));
    InMux I__4239 (
            .O(N__18838),
            .I(N__18820));
    InMux I__4238 (
            .O(N__18837),
            .I(N__18820));
    Span4Mux_v I__4237 (
            .O(N__18834),
            .I(N__18815));
    LocalMux I__4236 (
            .O(N__18831),
            .I(N__18815));
    Span4Mux_v I__4235 (
            .O(N__18828),
            .I(N__18812));
    LocalMux I__4234 (
            .O(N__18825),
            .I(N__18809));
    LocalMux I__4233 (
            .O(N__18820),
            .I(N__18806));
    Span4Mux_v I__4232 (
            .O(N__18815),
            .I(N__18799));
    Span4Mux_h I__4231 (
            .O(N__18812),
            .I(N__18799));
    Span4Mux_v I__4230 (
            .O(N__18809),
            .I(N__18799));
    Span4Mux_h I__4229 (
            .O(N__18806),
            .I(N__18796));
    Odrv4 I__4228 (
            .O(N__18799),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    Odrv4 I__4227 (
            .O(N__18796),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    InMux I__4226 (
            .O(N__18791),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__4225 (
            .O(N__18788),
            .I(N__18782));
    InMux I__4224 (
            .O(N__18787),
            .I(N__18782));
    LocalMux I__4223 (
            .O(N__18782),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i ));
    InMux I__4222 (
            .O(N__18779),
            .I(N__18759));
    InMux I__4221 (
            .O(N__18778),
            .I(N__18759));
    InMux I__4220 (
            .O(N__18777),
            .I(N__18759));
    InMux I__4219 (
            .O(N__18776),
            .I(N__18759));
    InMux I__4218 (
            .O(N__18775),
            .I(N__18759));
    InMux I__4217 (
            .O(N__18774),
            .I(N__18759));
    InMux I__4216 (
            .O(N__18773),
            .I(N__18754));
    InMux I__4215 (
            .O(N__18772),
            .I(N__18754));
    LocalMux I__4214 (
            .O(N__18759),
            .I(\delay_measurement_inst.N_41 ));
    LocalMux I__4213 (
            .O(N__18754),
            .I(\delay_measurement_inst.N_41 ));
    InMux I__4212 (
            .O(N__18749),
            .I(N__18745));
    InMux I__4211 (
            .O(N__18748),
            .I(N__18742));
    LocalMux I__4210 (
            .O(N__18745),
            .I(N__18736));
    LocalMux I__4209 (
            .O(N__18742),
            .I(N__18736));
    InMux I__4208 (
            .O(N__18741),
            .I(N__18733));
    Span4Mux_v I__4207 (
            .O(N__18736),
            .I(N__18728));
    LocalMux I__4206 (
            .O(N__18733),
            .I(N__18728));
    Odrv4 I__4205 (
            .O(N__18728),
            .I(\delay_measurement_inst.elapsed_time_tr_8 ));
    InMux I__4204 (
            .O(N__18725),
            .I(N__18722));
    LocalMux I__4203 (
            .O(N__18722),
            .I(N__18718));
    CascadeMux I__4202 (
            .O(N__18721),
            .I(N__18714));
    Span4Mux_v I__4201 (
            .O(N__18718),
            .I(N__18711));
    InMux I__4200 (
            .O(N__18717),
            .I(N__18708));
    InMux I__4199 (
            .O(N__18714),
            .I(N__18704));
    Sp12to4 I__4198 (
            .O(N__18711),
            .I(N__18699));
    LocalMux I__4197 (
            .O(N__18708),
            .I(N__18699));
    InMux I__4196 (
            .O(N__18707),
            .I(N__18696));
    LocalMux I__4195 (
            .O(N__18704),
            .I(measured_delay_tr_8));
    Odrv12 I__4194 (
            .O(N__18699),
            .I(measured_delay_tr_8));
    LocalMux I__4193 (
            .O(N__18696),
            .I(measured_delay_tr_8));
    CascadeMux I__4192 (
            .O(N__18689),
            .I(N__18684));
    CascadeMux I__4191 (
            .O(N__18688),
            .I(N__18673));
    InMux I__4190 (
            .O(N__18687),
            .I(N__18670));
    InMux I__4189 (
            .O(N__18684),
            .I(N__18667));
    InMux I__4188 (
            .O(N__18683),
            .I(N__18664));
    InMux I__4187 (
            .O(N__18682),
            .I(N__18649));
    InMux I__4186 (
            .O(N__18681),
            .I(N__18649));
    InMux I__4185 (
            .O(N__18680),
            .I(N__18649));
    InMux I__4184 (
            .O(N__18679),
            .I(N__18649));
    InMux I__4183 (
            .O(N__18678),
            .I(N__18649));
    InMux I__4182 (
            .O(N__18677),
            .I(N__18649));
    InMux I__4181 (
            .O(N__18676),
            .I(N__18649));
    InMux I__4180 (
            .O(N__18673),
            .I(N__18644));
    LocalMux I__4179 (
            .O(N__18670),
            .I(N__18641));
    LocalMux I__4178 (
            .O(N__18667),
            .I(N__18634));
    LocalMux I__4177 (
            .O(N__18664),
            .I(N__18634));
    LocalMux I__4176 (
            .O(N__18649),
            .I(N__18634));
    InMux I__4175 (
            .O(N__18648),
            .I(N__18629));
    InMux I__4174 (
            .O(N__18647),
            .I(N__18629));
    LocalMux I__4173 (
            .O(N__18644),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    Odrv4 I__4172 (
            .O(N__18641),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    Odrv4 I__4171 (
            .O(N__18634),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    LocalMux I__4170 (
            .O(N__18629),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    InMux I__4169 (
            .O(N__18620),
            .I(N__18617));
    LocalMux I__4168 (
            .O(N__18617),
            .I(N__18613));
    CascadeMux I__4167 (
            .O(N__18616),
            .I(N__18609));
    Span4Mux_v I__4166 (
            .O(N__18613),
            .I(N__18606));
    InMux I__4165 (
            .O(N__18612),
            .I(N__18603));
    InMux I__4164 (
            .O(N__18609),
            .I(N__18600));
    Odrv4 I__4163 (
            .O(N__18606),
            .I(\delay_measurement_inst.elapsed_time_tr_19 ));
    LocalMux I__4162 (
            .O(N__18603),
            .I(\delay_measurement_inst.elapsed_time_tr_19 ));
    LocalMux I__4161 (
            .O(N__18600),
            .I(\delay_measurement_inst.elapsed_time_tr_19 ));
    InMux I__4160 (
            .O(N__18593),
            .I(N__18583));
    InMux I__4159 (
            .O(N__18592),
            .I(N__18583));
    InMux I__4158 (
            .O(N__18591),
            .I(N__18583));
    InMux I__4157 (
            .O(N__18590),
            .I(N__18580));
    LocalMux I__4156 (
            .O(N__18583),
            .I(N__18570));
    LocalMux I__4155 (
            .O(N__18580),
            .I(N__18570));
    InMux I__4154 (
            .O(N__18579),
            .I(N__18567));
    InMux I__4153 (
            .O(N__18578),
            .I(N__18558));
    InMux I__4152 (
            .O(N__18577),
            .I(N__18558));
    InMux I__4151 (
            .O(N__18576),
            .I(N__18558));
    InMux I__4150 (
            .O(N__18575),
            .I(N__18558));
    Odrv4 I__4149 (
            .O(N__18570),
            .I(\delay_measurement_inst.N_35 ));
    LocalMux I__4148 (
            .O(N__18567),
            .I(\delay_measurement_inst.N_35 ));
    LocalMux I__4147 (
            .O(N__18558),
            .I(\delay_measurement_inst.N_35 ));
    InMux I__4146 (
            .O(N__18551),
            .I(N__18548));
    LocalMux I__4145 (
            .O(N__18548),
            .I(N__18543));
    InMux I__4144 (
            .O(N__18547),
            .I(N__18540));
    CascadeMux I__4143 (
            .O(N__18546),
            .I(N__18537));
    Span4Mux_v I__4142 (
            .O(N__18543),
            .I(N__18534));
    LocalMux I__4141 (
            .O(N__18540),
            .I(N__18531));
    InMux I__4140 (
            .O(N__18537),
            .I(N__18528));
    Span4Mux_h I__4139 (
            .O(N__18534),
            .I(N__18520));
    Span4Mux_v I__4138 (
            .O(N__18531),
            .I(N__18520));
    LocalMux I__4137 (
            .O(N__18528),
            .I(N__18520));
    CascadeMux I__4136 (
            .O(N__18527),
            .I(N__18517));
    Span4Mux_h I__4135 (
            .O(N__18520),
            .I(N__18514));
    InMux I__4134 (
            .O(N__18517),
            .I(N__18511));
    Odrv4 I__4133 (
            .O(N__18514),
            .I(measured_delay_tr_19));
    LocalMux I__4132 (
            .O(N__18511),
            .I(measured_delay_tr_19));
    CEMux I__4131 (
            .O(N__18506),
            .I(N__18502));
    CEMux I__4130 (
            .O(N__18505),
            .I(N__18498));
    LocalMux I__4129 (
            .O(N__18502),
            .I(N__18495));
    CEMux I__4128 (
            .O(N__18501),
            .I(N__18492));
    LocalMux I__4127 (
            .O(N__18498),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ));
    Odrv12 I__4126 (
            .O(N__18495),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ));
    LocalMux I__4125 (
            .O(N__18492),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ));
    InMux I__4124 (
            .O(N__18485),
            .I(N__18480));
    InMux I__4123 (
            .O(N__18484),
            .I(N__18477));
    InMux I__4122 (
            .O(N__18483),
            .I(N__18474));
    LocalMux I__4121 (
            .O(N__18480),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__4120 (
            .O(N__18477),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__4119 (
            .O(N__18474),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    CascadeMux I__4118 (
            .O(N__18467),
            .I(N__18464));
    InMux I__4117 (
            .O(N__18464),
            .I(N__18459));
    InMux I__4116 (
            .O(N__18463),
            .I(N__18454));
    InMux I__4115 (
            .O(N__18462),
            .I(N__18454));
    LocalMux I__4114 (
            .O(N__18459),
            .I(N__18449));
    LocalMux I__4113 (
            .O(N__18454),
            .I(N__18449));
    Span4Mux_h I__4112 (
            .O(N__18449),
            .I(N__18446));
    Odrv4 I__4111 (
            .O(N__18446),
            .I(\delay_measurement_inst.elapsed_time_hc_3 ));
    InMux I__4110 (
            .O(N__18443),
            .I(N__18438));
    InMux I__4109 (
            .O(N__18442),
            .I(N__18435));
    InMux I__4108 (
            .O(N__18441),
            .I(N__18432));
    LocalMux I__4107 (
            .O(N__18438),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__4106 (
            .O(N__18435),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__4105 (
            .O(N__18432),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    CascadeMux I__4104 (
            .O(N__18425),
            .I(N__18422));
    InMux I__4103 (
            .O(N__18422),
            .I(N__18419));
    LocalMux I__4102 (
            .O(N__18419),
            .I(N__18416));
    Span4Mux_v I__4101 (
            .O(N__18416),
            .I(N__18412));
    InMux I__4100 (
            .O(N__18415),
            .I(N__18409));
    Sp12to4 I__4099 (
            .O(N__18412),
            .I(N__18404));
    LocalMux I__4098 (
            .O(N__18409),
            .I(N__18404));
    Odrv12 I__4097 (
            .O(N__18404),
            .I(\delay_measurement_inst.elapsed_time_hc_4 ));
    InMux I__4096 (
            .O(N__18401),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__4095 (
            .O(N__18398),
            .I(N__18393));
    CascadeMux I__4094 (
            .O(N__18397),
            .I(N__18390));
    InMux I__4093 (
            .O(N__18396),
            .I(N__18387));
    InMux I__4092 (
            .O(N__18393),
            .I(N__18382));
    InMux I__4091 (
            .O(N__18390),
            .I(N__18382));
    LocalMux I__4090 (
            .O(N__18387),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    LocalMux I__4089 (
            .O(N__18382),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__4088 (
            .O(N__18377),
            .I(N__18374));
    LocalMux I__4087 (
            .O(N__18374),
            .I(N__18370));
    InMux I__4086 (
            .O(N__18373),
            .I(N__18367));
    Span4Mux_v I__4085 (
            .O(N__18370),
            .I(N__18362));
    LocalMux I__4084 (
            .O(N__18367),
            .I(N__18362));
    Odrv4 I__4083 (
            .O(N__18362),
            .I(\delay_measurement_inst.elapsed_time_hc_5 ));
    InMux I__4082 (
            .O(N__18359),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__4081 (
            .O(N__18356),
            .I(N__18351));
    CascadeMux I__4080 (
            .O(N__18355),
            .I(N__18348));
    InMux I__4079 (
            .O(N__18354),
            .I(N__18345));
    InMux I__4078 (
            .O(N__18351),
            .I(N__18340));
    InMux I__4077 (
            .O(N__18348),
            .I(N__18340));
    LocalMux I__4076 (
            .O(N__18345),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    LocalMux I__4075 (
            .O(N__18340),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    CascadeMux I__4074 (
            .O(N__18335),
            .I(N__18332));
    InMux I__4073 (
            .O(N__18332),
            .I(N__18327));
    InMux I__4072 (
            .O(N__18331),
            .I(N__18321));
    InMux I__4071 (
            .O(N__18330),
            .I(N__18321));
    LocalMux I__4070 (
            .O(N__18327),
            .I(N__18318));
    InMux I__4069 (
            .O(N__18326),
            .I(N__18315));
    LocalMux I__4068 (
            .O(N__18321),
            .I(N__18312));
    Span4Mux_v I__4067 (
            .O(N__18318),
            .I(N__18307));
    LocalMux I__4066 (
            .O(N__18315),
            .I(N__18307));
    Span4Mux_h I__4065 (
            .O(N__18312),
            .I(N__18304));
    Odrv4 I__4064 (
            .O(N__18307),
            .I(\delay_measurement_inst.delay_hc_reg3lto6 ));
    Odrv4 I__4063 (
            .O(N__18304),
            .I(\delay_measurement_inst.delay_hc_reg3lto6 ));
    InMux I__4062 (
            .O(N__18299),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__4061 (
            .O(N__18296),
            .I(N__18291));
    InMux I__4060 (
            .O(N__18295),
            .I(N__18286));
    InMux I__4059 (
            .O(N__18294),
            .I(N__18286));
    LocalMux I__4058 (
            .O(N__18291),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    LocalMux I__4057 (
            .O(N__18286),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    CascadeMux I__4056 (
            .O(N__18281),
            .I(N__18278));
    InMux I__4055 (
            .O(N__18278),
            .I(N__18274));
    InMux I__4054 (
            .O(N__18277),
            .I(N__18271));
    LocalMux I__4053 (
            .O(N__18274),
            .I(N__18268));
    LocalMux I__4052 (
            .O(N__18271),
            .I(N__18265));
    Span4Mux_h I__4051 (
            .O(N__18268),
            .I(N__18262));
    Span4Mux_h I__4050 (
            .O(N__18265),
            .I(N__18259));
    Odrv4 I__4049 (
            .O(N__18262),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    Odrv4 I__4048 (
            .O(N__18259),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    InMux I__4047 (
            .O(N__18254),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__4046 (
            .O(N__18251),
            .I(N__18246));
    InMux I__4045 (
            .O(N__18250),
            .I(N__18241));
    InMux I__4044 (
            .O(N__18249),
            .I(N__18241));
    LocalMux I__4043 (
            .O(N__18246),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    LocalMux I__4042 (
            .O(N__18241),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    CascadeMux I__4041 (
            .O(N__18236),
            .I(N__18232));
    CascadeMux I__4040 (
            .O(N__18235),
            .I(N__18229));
    InMux I__4039 (
            .O(N__18232),
            .I(N__18226));
    InMux I__4038 (
            .O(N__18229),
            .I(N__18223));
    LocalMux I__4037 (
            .O(N__18226),
            .I(N__18220));
    LocalMux I__4036 (
            .O(N__18223),
            .I(N__18217));
    Span4Mux_h I__4035 (
            .O(N__18220),
            .I(N__18214));
    Span4Mux_h I__4034 (
            .O(N__18217),
            .I(N__18211));
    Odrv4 I__4033 (
            .O(N__18214),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    Odrv4 I__4032 (
            .O(N__18211),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    InMux I__4031 (
            .O(N__18206),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__4030 (
            .O(N__18203),
            .I(N__18200));
    LocalMux I__4029 (
            .O(N__18200),
            .I(\delay_measurement_inst.N_164 ));
    InMux I__4028 (
            .O(N__18197),
            .I(N__18179));
    InMux I__4027 (
            .O(N__18196),
            .I(N__18179));
    InMux I__4026 (
            .O(N__18195),
            .I(N__18179));
    InMux I__4025 (
            .O(N__18194),
            .I(N__18179));
    InMux I__4024 (
            .O(N__18193),
            .I(N__18179));
    InMux I__4023 (
            .O(N__18192),
            .I(N__18179));
    LocalMux I__4022 (
            .O(N__18179),
            .I(\delay_measurement_inst.N_187 ));
    InMux I__4021 (
            .O(N__18176),
            .I(N__18173));
    LocalMux I__4020 (
            .O(N__18173),
            .I(N__18170));
    Odrv4 I__4019 (
            .O(N__18170),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_7 ));
    CascadeMux I__4018 (
            .O(N__18167),
            .I(\delay_measurement_inst.N_187_cascade_ ));
    InMux I__4017 (
            .O(N__18164),
            .I(N__18161));
    LocalMux I__4016 (
            .O(N__18161),
            .I(\delay_measurement_inst.delay_tr_timer.N_177 ));
    CascadeMux I__4015 (
            .O(N__18158),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_cascade_ ));
    CascadeMux I__4014 (
            .O(N__18155),
            .I(N__18152));
    InMux I__4013 (
            .O(N__18152),
            .I(N__18136));
    InMux I__4012 (
            .O(N__18151),
            .I(N__18136));
    InMux I__4011 (
            .O(N__18150),
            .I(N__18136));
    InMux I__4010 (
            .O(N__18149),
            .I(N__18136));
    InMux I__4009 (
            .O(N__18148),
            .I(N__18136));
    InMux I__4008 (
            .O(N__18147),
            .I(N__18133));
    LocalMux I__4007 (
            .O(N__18136),
            .I(\delay_measurement_inst.N_162_1 ));
    LocalMux I__4006 (
            .O(N__18133),
            .I(\delay_measurement_inst.N_162_1 ));
    CascadeMux I__4005 (
            .O(N__18128),
            .I(N__18123));
    InMux I__4004 (
            .O(N__18127),
            .I(N__18115));
    InMux I__4003 (
            .O(N__18126),
            .I(N__18115));
    InMux I__4002 (
            .O(N__18123),
            .I(N__18115));
    InMux I__4001 (
            .O(N__18122),
            .I(N__18112));
    LocalMux I__4000 (
            .O(N__18115),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10 ));
    LocalMux I__3999 (
            .O(N__18112),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10 ));
    CascadeMux I__3998 (
            .O(N__18107),
            .I(N__18102));
    CascadeMux I__3997 (
            .O(N__18106),
            .I(N__18099));
    InMux I__3996 (
            .O(N__18105),
            .I(N__18096));
    InMux I__3995 (
            .O(N__18102),
            .I(N__18093));
    InMux I__3994 (
            .O(N__18099),
            .I(N__18090));
    LocalMux I__3993 (
            .O(N__18096),
            .I(N__18086));
    LocalMux I__3992 (
            .O(N__18093),
            .I(N__18081));
    LocalMux I__3991 (
            .O(N__18090),
            .I(N__18081));
    InMux I__3990 (
            .O(N__18089),
            .I(N__18078));
    Span4Mux_v I__3989 (
            .O(N__18086),
            .I(N__18074));
    Span4Mux_v I__3988 (
            .O(N__18081),
            .I(N__18069));
    LocalMux I__3987 (
            .O(N__18078),
            .I(N__18069));
    InMux I__3986 (
            .O(N__18077),
            .I(N__18066));
    Odrv4 I__3985 (
            .O(N__18074),
            .I(\delay_measurement_inst.delay_tr_reg3lto9 ));
    Odrv4 I__3984 (
            .O(N__18069),
            .I(\delay_measurement_inst.delay_tr_reg3lto9 ));
    LocalMux I__3983 (
            .O(N__18066),
            .I(\delay_measurement_inst.delay_tr_reg3lto9 ));
    InMux I__3982 (
            .O(N__18059),
            .I(N__18053));
    InMux I__3981 (
            .O(N__18058),
            .I(N__18050));
    InMux I__3980 (
            .O(N__18057),
            .I(N__18047));
    CascadeMux I__3979 (
            .O(N__18056),
            .I(N__18044));
    LocalMux I__3978 (
            .O(N__18053),
            .I(N__18040));
    LocalMux I__3977 (
            .O(N__18050),
            .I(N__18035));
    LocalMux I__3976 (
            .O(N__18047),
            .I(N__18035));
    InMux I__3975 (
            .O(N__18044),
            .I(N__18030));
    InMux I__3974 (
            .O(N__18043),
            .I(N__18030));
    Odrv12 I__3973 (
            .O(N__18040),
            .I(\delay_measurement_inst.delay_tr_reg3lto14 ));
    Odrv4 I__3972 (
            .O(N__18035),
            .I(\delay_measurement_inst.delay_tr_reg3lto14 ));
    LocalMux I__3971 (
            .O(N__18030),
            .I(\delay_measurement_inst.delay_tr_reg3lto14 ));
    InMux I__3970 (
            .O(N__18023),
            .I(N__18019));
    CascadeMux I__3969 (
            .O(N__18022),
            .I(N__18015));
    LocalMux I__3968 (
            .O(N__18019),
            .I(N__18012));
    InMux I__3967 (
            .O(N__18018),
            .I(N__18009));
    InMux I__3966 (
            .O(N__18015),
            .I(N__18006));
    Span4Mux_h I__3965 (
            .O(N__18012),
            .I(N__18002));
    LocalMux I__3964 (
            .O(N__18009),
            .I(N__17999));
    LocalMux I__3963 (
            .O(N__18006),
            .I(N__17996));
    InMux I__3962 (
            .O(N__18005),
            .I(N__17993));
    Odrv4 I__3961 (
            .O(N__18002),
            .I(\delay_measurement_inst.N_39 ));
    Odrv4 I__3960 (
            .O(N__17999),
            .I(\delay_measurement_inst.N_39 ));
    Odrv4 I__3959 (
            .O(N__17996),
            .I(\delay_measurement_inst.N_39 ));
    LocalMux I__3958 (
            .O(N__17993),
            .I(\delay_measurement_inst.N_39 ));
    CascadeMux I__3957 (
            .O(N__17984),
            .I(\delay_measurement_inst.delay_tr_timer.N_180_cascade_ ));
    CascadeMux I__3956 (
            .O(N__17981),
            .I(N__17978));
    InMux I__3955 (
            .O(N__17978),
            .I(N__17974));
    InMux I__3954 (
            .O(N__17977),
            .I(N__17971));
    LocalMux I__3953 (
            .O(N__17974),
            .I(N__17967));
    LocalMux I__3952 (
            .O(N__17971),
            .I(N__17964));
    InMux I__3951 (
            .O(N__17970),
            .I(N__17961));
    Span4Mux_v I__3950 (
            .O(N__17967),
            .I(N__17957));
    Span4Mux_v I__3949 (
            .O(N__17964),
            .I(N__17952));
    LocalMux I__3948 (
            .O(N__17961),
            .I(N__17952));
    InMux I__3947 (
            .O(N__17960),
            .I(N__17949));
    Odrv4 I__3946 (
            .O(N__17957),
            .I(\delay_measurement_inst.delay_tr_reg3lto6 ));
    Odrv4 I__3945 (
            .O(N__17952),
            .I(\delay_measurement_inst.delay_tr_reg3lto6 ));
    LocalMux I__3944 (
            .O(N__17949),
            .I(\delay_measurement_inst.delay_tr_reg3lto6 ));
    InMux I__3943 (
            .O(N__17942),
            .I(N__17932));
    InMux I__3942 (
            .O(N__17941),
            .I(N__17932));
    InMux I__3941 (
            .O(N__17940),
            .I(N__17927));
    InMux I__3940 (
            .O(N__17939),
            .I(N__17927));
    InMux I__3939 (
            .O(N__17938),
            .I(N__17922));
    InMux I__3938 (
            .O(N__17937),
            .I(N__17922));
    LocalMux I__3937 (
            .O(N__17932),
            .I(N__17913));
    LocalMux I__3936 (
            .O(N__17927),
            .I(N__17913));
    LocalMux I__3935 (
            .O(N__17922),
            .I(N__17913));
    InMux I__3934 (
            .O(N__17921),
            .I(N__17908));
    InMux I__3933 (
            .O(N__17920),
            .I(N__17908));
    Odrv4 I__3932 (
            .O(N__17913),
            .I(\delay_measurement_inst.delay_tr_reg3lto15 ));
    LocalMux I__3931 (
            .O(N__17908),
            .I(\delay_measurement_inst.delay_tr_reg3lto15 ));
    CascadeMux I__3930 (
            .O(N__17903),
            .I(N__17896));
    CascadeMux I__3929 (
            .O(N__17902),
            .I(N__17893));
    InMux I__3928 (
            .O(N__17901),
            .I(N__17882));
    InMux I__3927 (
            .O(N__17900),
            .I(N__17882));
    InMux I__3926 (
            .O(N__17899),
            .I(N__17882));
    InMux I__3925 (
            .O(N__17896),
            .I(N__17882));
    InMux I__3924 (
            .O(N__17893),
            .I(N__17882));
    LocalMux I__3923 (
            .O(N__17882),
            .I(\delay_measurement_inst.delay_tr_reg_5_0_a2_0_6 ));
    InMux I__3922 (
            .O(N__17879),
            .I(N__17875));
    InMux I__3921 (
            .O(N__17878),
            .I(N__17872));
    LocalMux I__3920 (
            .O(N__17875),
            .I(N__17866));
    LocalMux I__3919 (
            .O(N__17872),
            .I(N__17866));
    InMux I__3918 (
            .O(N__17871),
            .I(N__17863));
    Span4Mux_v I__3917 (
            .O(N__17866),
            .I(N__17858));
    LocalMux I__3916 (
            .O(N__17863),
            .I(N__17858));
    Odrv4 I__3915 (
            .O(N__17858),
            .I(\delay_measurement_inst.elapsed_time_tr_7 ));
    InMux I__3914 (
            .O(N__17855),
            .I(N__17852));
    LocalMux I__3913 (
            .O(N__17852),
            .I(N__17846));
    InMux I__3912 (
            .O(N__17851),
            .I(N__17843));
    CascadeMux I__3911 (
            .O(N__17850),
            .I(N__17840));
    CascadeMux I__3910 (
            .O(N__17849),
            .I(N__17837));
    Span4Mux_v I__3909 (
            .O(N__17846),
            .I(N__17834));
    LocalMux I__3908 (
            .O(N__17843),
            .I(N__17831));
    InMux I__3907 (
            .O(N__17840),
            .I(N__17828));
    InMux I__3906 (
            .O(N__17837),
            .I(N__17825));
    Span4Mux_h I__3905 (
            .O(N__17834),
            .I(N__17820));
    Span4Mux_h I__3904 (
            .O(N__17831),
            .I(N__17820));
    LocalMux I__3903 (
            .O(N__17828),
            .I(N__17817));
    LocalMux I__3902 (
            .O(N__17825),
            .I(measured_delay_tr_7));
    Odrv4 I__3901 (
            .O(N__17820),
            .I(measured_delay_tr_7));
    Odrv4 I__3900 (
            .O(N__17817),
            .I(measured_delay_tr_7));
    InMux I__3899 (
            .O(N__17810),
            .I(N__17804));
    InMux I__3898 (
            .O(N__17809),
            .I(N__17804));
    LocalMux I__3897 (
            .O(N__17804),
            .I(\delay_measurement_inst.delay_tr_timer.N_177_4 ));
    InMux I__3896 (
            .O(N__17801),
            .I(N__17798));
    LocalMux I__3895 (
            .O(N__17798),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_4 ));
    CascadeMux I__3894 (
            .O(N__17795),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3_cascade_ ));
    InMux I__3893 (
            .O(N__17792),
            .I(N__17789));
    LocalMux I__3892 (
            .O(N__17789),
            .I(N__17784));
    InMux I__3891 (
            .O(N__17788),
            .I(N__17779));
    InMux I__3890 (
            .O(N__17787),
            .I(N__17779));
    Odrv12 I__3889 (
            .O(N__17784),
            .I(\delay_measurement_inst.elapsed_time_tr_16 ));
    LocalMux I__3888 (
            .O(N__17779),
            .I(\delay_measurement_inst.elapsed_time_tr_16 ));
    InMux I__3887 (
            .O(N__17774),
            .I(N__17770));
    CascadeMux I__3886 (
            .O(N__17773),
            .I(N__17766));
    LocalMux I__3885 (
            .O(N__17770),
            .I(N__17763));
    InMux I__3884 (
            .O(N__17769),
            .I(N__17760));
    InMux I__3883 (
            .O(N__17766),
            .I(N__17757));
    Odrv12 I__3882 (
            .O(N__17763),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    LocalMux I__3881 (
            .O(N__17760),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    LocalMux I__3880 (
            .O(N__17757),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    InMux I__3879 (
            .O(N__17750),
            .I(N__17747));
    LocalMux I__3878 (
            .O(N__17747),
            .I(N__17742));
    InMux I__3877 (
            .O(N__17746),
            .I(N__17739));
    InMux I__3876 (
            .O(N__17745),
            .I(N__17736));
    Odrv12 I__3875 (
            .O(N__17742),
            .I(\delay_measurement_inst.elapsed_time_tr_18 ));
    LocalMux I__3874 (
            .O(N__17739),
            .I(\delay_measurement_inst.elapsed_time_tr_18 ));
    LocalMux I__3873 (
            .O(N__17736),
            .I(\delay_measurement_inst.elapsed_time_tr_18 ));
    InMux I__3872 (
            .O(N__17729),
            .I(N__17726));
    LocalMux I__3871 (
            .O(N__17726),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ));
    InMux I__3870 (
            .O(N__17723),
            .I(N__17720));
    LocalMux I__3869 (
            .O(N__17720),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__3868 (
            .O(N__17717),
            .I(N__17713));
    InMux I__3867 (
            .O(N__17716),
            .I(N__17710));
    LocalMux I__3866 (
            .O(N__17713),
            .I(N__17707));
    LocalMux I__3865 (
            .O(N__17710),
            .I(N__17704));
    Span4Mux_h I__3864 (
            .O(N__17707),
            .I(N__17701));
    Odrv12 I__3863 (
            .O(N__17704),
            .I(\delay_measurement_inst.elapsed_time_tr_12 ));
    Odrv4 I__3862 (
            .O(N__17701),
            .I(\delay_measurement_inst.elapsed_time_tr_12 ));
    InMux I__3861 (
            .O(N__17696),
            .I(N__17692));
    InMux I__3860 (
            .O(N__17695),
            .I(N__17689));
    LocalMux I__3859 (
            .O(N__17692),
            .I(N__17686));
    LocalMux I__3858 (
            .O(N__17689),
            .I(N__17683));
    Span4Mux_h I__3857 (
            .O(N__17686),
            .I(N__17680));
    Odrv12 I__3856 (
            .O(N__17683),
            .I(\delay_measurement_inst.elapsed_time_tr_11 ));
    Odrv4 I__3855 (
            .O(N__17680),
            .I(\delay_measurement_inst.elapsed_time_tr_11 ));
    InMux I__3854 (
            .O(N__17675),
            .I(N__17671));
    CascadeMux I__3853 (
            .O(N__17674),
            .I(N__17668));
    LocalMux I__3852 (
            .O(N__17671),
            .I(N__17665));
    InMux I__3851 (
            .O(N__17668),
            .I(N__17662));
    Span4Mux_v I__3850 (
            .O(N__17665),
            .I(N__17657));
    LocalMux I__3849 (
            .O(N__17662),
            .I(N__17657));
    Odrv4 I__3848 (
            .O(N__17657),
            .I(\delay_measurement_inst.elapsed_time_tr_13 ));
    InMux I__3847 (
            .O(N__17654),
            .I(N__17650));
    InMux I__3846 (
            .O(N__17653),
            .I(N__17647));
    LocalMux I__3845 (
            .O(N__17650),
            .I(N__17644));
    LocalMux I__3844 (
            .O(N__17647),
            .I(N__17641));
    Odrv12 I__3843 (
            .O(N__17644),
            .I(\delay_measurement_inst.elapsed_time_tr_10 ));
    Odrv4 I__3842 (
            .O(N__17641),
            .I(\delay_measurement_inst.elapsed_time_tr_10 ));
    InMux I__3841 (
            .O(N__17636),
            .I(N__17633));
    LocalMux I__3840 (
            .O(N__17633),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__3839 (
            .O(N__17630),
            .I(N__17627));
    LocalMux I__3838 (
            .O(N__17627),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    CascadeMux I__3837 (
            .O(N__17624),
            .I(N__17621));
    InMux I__3836 (
            .O(N__17621),
            .I(N__17618));
    LocalMux I__3835 (
            .O(N__17618),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__3834 (
            .O(N__17615),
            .I(N__17612));
    LocalMux I__3833 (
            .O(N__17612),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__3832 (
            .O(N__17609),
            .I(N__17606));
    LocalMux I__3831 (
            .O(N__17606),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__3830 (
            .O(N__17603),
            .I(N__17600));
    LocalMux I__3829 (
            .O(N__17600),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19 ));
    CascadeMux I__3828 (
            .O(N__17597),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19_cascade_ ));
    InMux I__3827 (
            .O(N__17594),
            .I(N__17591));
    LocalMux I__3826 (
            .O(N__17591),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19 ));
    InMux I__3825 (
            .O(N__17588),
            .I(N__17585));
    LocalMux I__3824 (
            .O(N__17585),
            .I(N__17582));
    Odrv4 I__3823 (
            .O(N__17582),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6 ));
    CascadeMux I__3822 (
            .O(N__17579),
            .I(\delay_measurement_inst.N_35_cascade_ ));
    InMux I__3821 (
            .O(N__17576),
            .I(N__17573));
    LocalMux I__3820 (
            .O(N__17573),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_7 ));
    CascadeMux I__3819 (
            .O(N__17570),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_ ));
    InMux I__3818 (
            .O(N__17567),
            .I(N__17533));
    InMux I__3817 (
            .O(N__17566),
            .I(N__17533));
    InMux I__3816 (
            .O(N__17565),
            .I(N__17533));
    InMux I__3815 (
            .O(N__17564),
            .I(N__17533));
    InMux I__3814 (
            .O(N__17563),
            .I(N__17524));
    InMux I__3813 (
            .O(N__17562),
            .I(N__17524));
    InMux I__3812 (
            .O(N__17561),
            .I(N__17515));
    InMux I__3811 (
            .O(N__17560),
            .I(N__17515));
    InMux I__3810 (
            .O(N__17559),
            .I(N__17515));
    InMux I__3809 (
            .O(N__17558),
            .I(N__17515));
    InMux I__3808 (
            .O(N__17557),
            .I(N__17506));
    InMux I__3807 (
            .O(N__17556),
            .I(N__17506));
    InMux I__3806 (
            .O(N__17555),
            .I(N__17506));
    InMux I__3805 (
            .O(N__17554),
            .I(N__17506));
    InMux I__3804 (
            .O(N__17553),
            .I(N__17497));
    InMux I__3803 (
            .O(N__17552),
            .I(N__17497));
    InMux I__3802 (
            .O(N__17551),
            .I(N__17497));
    InMux I__3801 (
            .O(N__17550),
            .I(N__17497));
    InMux I__3800 (
            .O(N__17549),
            .I(N__17488));
    InMux I__3799 (
            .O(N__17548),
            .I(N__17488));
    InMux I__3798 (
            .O(N__17547),
            .I(N__17488));
    InMux I__3797 (
            .O(N__17546),
            .I(N__17488));
    InMux I__3796 (
            .O(N__17545),
            .I(N__17479));
    InMux I__3795 (
            .O(N__17544),
            .I(N__17479));
    InMux I__3794 (
            .O(N__17543),
            .I(N__17479));
    InMux I__3793 (
            .O(N__17542),
            .I(N__17479));
    LocalMux I__3792 (
            .O(N__17533),
            .I(N__17476));
    InMux I__3791 (
            .O(N__17532),
            .I(N__17467));
    InMux I__3790 (
            .O(N__17531),
            .I(N__17467));
    InMux I__3789 (
            .O(N__17530),
            .I(N__17467));
    InMux I__3788 (
            .O(N__17529),
            .I(N__17467));
    LocalMux I__3787 (
            .O(N__17524),
            .I(N__17464));
    LocalMux I__3786 (
            .O(N__17515),
            .I(N__17459));
    LocalMux I__3785 (
            .O(N__17506),
            .I(N__17459));
    LocalMux I__3784 (
            .O(N__17497),
            .I(N__17452));
    LocalMux I__3783 (
            .O(N__17488),
            .I(N__17452));
    LocalMux I__3782 (
            .O(N__17479),
            .I(N__17452));
    Span4Mux_v I__3781 (
            .O(N__17476),
            .I(N__17441));
    LocalMux I__3780 (
            .O(N__17467),
            .I(N__17441));
    Span4Mux_v I__3779 (
            .O(N__17464),
            .I(N__17441));
    Span4Mux_v I__3778 (
            .O(N__17459),
            .I(N__17441));
    Span4Mux_v I__3777 (
            .O(N__17452),
            .I(N__17441));
    Odrv4 I__3776 (
            .O(N__17441),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    CascadeMux I__3775 (
            .O(N__17438),
            .I(N__17435));
    InMux I__3774 (
            .O(N__17435),
            .I(N__17432));
    LocalMux I__3773 (
            .O(N__17432),
            .I(N__17429));
    Span4Mux_v I__3772 (
            .O(N__17429),
            .I(N__17425));
    InMux I__3771 (
            .O(N__17428),
            .I(N__17422));
    Odrv4 I__3770 (
            .O(N__17425),
            .I(\delay_measurement_inst.elapsed_time_tr_5 ));
    LocalMux I__3769 (
            .O(N__17422),
            .I(\delay_measurement_inst.elapsed_time_tr_5 ));
    InMux I__3768 (
            .O(N__17417),
            .I(N__17414));
    LocalMux I__3767 (
            .O(N__17414),
            .I(N__17410));
    InMux I__3766 (
            .O(N__17413),
            .I(N__17407));
    Odrv12 I__3765 (
            .O(N__17410),
            .I(\delay_measurement_inst.elapsed_time_tr_4 ));
    LocalMux I__3764 (
            .O(N__17407),
            .I(\delay_measurement_inst.elapsed_time_tr_4 ));
    CascadeMux I__3763 (
            .O(N__17402),
            .I(N__17399));
    InMux I__3762 (
            .O(N__17399),
            .I(N__17396));
    LocalMux I__3761 (
            .O(N__17396),
            .I(N__17392));
    InMux I__3760 (
            .O(N__17395),
            .I(N__17389));
    Span4Mux_v I__3759 (
            .O(N__17392),
            .I(N__17383));
    LocalMux I__3758 (
            .O(N__17389),
            .I(N__17383));
    InMux I__3757 (
            .O(N__17388),
            .I(N__17380));
    Odrv4 I__3756 (
            .O(N__17383),
            .I(\delay_measurement_inst.elapsed_time_tr_3 ));
    LocalMux I__3755 (
            .O(N__17380),
            .I(\delay_measurement_inst.elapsed_time_tr_3 ));
    CascadeMux I__3754 (
            .O(N__17375),
            .I(N__17372));
    InMux I__3753 (
            .O(N__17372),
            .I(N__17368));
    CascadeMux I__3752 (
            .O(N__17371),
            .I(N__17365));
    LocalMux I__3751 (
            .O(N__17368),
            .I(N__17362));
    InMux I__3750 (
            .O(N__17365),
            .I(N__17359));
    Span4Mux_v I__3749 (
            .O(N__17362),
            .I(N__17356));
    LocalMux I__3748 (
            .O(N__17359),
            .I(N__17353));
    Odrv4 I__3747 (
            .O(N__17356),
            .I(\delay_measurement_inst.elapsed_time_tr_1 ));
    Odrv12 I__3746 (
            .O(N__17353),
            .I(\delay_measurement_inst.elapsed_time_tr_1 ));
    InMux I__3745 (
            .O(N__17348),
            .I(N__17345));
    LocalMux I__3744 (
            .O(N__17345),
            .I(N__17341));
    InMux I__3743 (
            .O(N__17344),
            .I(N__17338));
    Span4Mux_v I__3742 (
            .O(N__17341),
            .I(N__17332));
    LocalMux I__3741 (
            .O(N__17338),
            .I(N__17332));
    InMux I__3740 (
            .O(N__17337),
            .I(N__17329));
    Odrv4 I__3739 (
            .O(N__17332),
            .I(\delay_measurement_inst.elapsed_time_tr_2 ));
    LocalMux I__3738 (
            .O(N__17329),
            .I(\delay_measurement_inst.elapsed_time_tr_2 ));
    InMux I__3737 (
            .O(N__17324),
            .I(N__17321));
    LocalMux I__3736 (
            .O(N__17321),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__3735 (
            .O(N__17318),
            .I(N__17315));
    LocalMux I__3734 (
            .O(N__17315),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    CascadeMux I__3733 (
            .O(N__17312),
            .I(N__17309));
    InMux I__3732 (
            .O(N__17309),
            .I(N__17306));
    LocalMux I__3731 (
            .O(N__17306),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    InMux I__3730 (
            .O(N__17303),
            .I(N__17300));
    LocalMux I__3729 (
            .O(N__17300),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    CascadeMux I__3728 (
            .O(N__17297),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5_cascade_ ));
    InMux I__3727 (
            .O(N__17294),
            .I(bfn_9_24_0_));
    InMux I__3726 (
            .O(N__17291),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    InMux I__3725 (
            .O(N__17288),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    InMux I__3724 (
            .O(N__17285),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    InMux I__3723 (
            .O(N__17282),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__3722 (
            .O(N__17279),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    InMux I__3721 (
            .O(N__17276),
            .I(N__17273));
    LocalMux I__3720 (
            .O(N__17273),
            .I(N__17270));
    Span4Mux_s1_v I__3719 (
            .O(N__17270),
            .I(N__17267));
    Span4Mux_v I__3718 (
            .O(N__17267),
            .I(N__17261));
    InMux I__3717 (
            .O(N__17266),
            .I(N__17258));
    InMux I__3716 (
            .O(N__17265),
            .I(N__17255));
    InMux I__3715 (
            .O(N__17264),
            .I(N__17252));
    Odrv4 I__3714 (
            .O(N__17261),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    LocalMux I__3713 (
            .O(N__17258),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    LocalMux I__3712 (
            .O(N__17255),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    LocalMux I__3711 (
            .O(N__17252),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    IoInMux I__3710 (
            .O(N__17243),
            .I(N__17240));
    LocalMux I__3709 (
            .O(N__17240),
            .I(s3_phy_c));
    InMux I__3708 (
            .O(N__17237),
            .I(N__17234));
    LocalMux I__3707 (
            .O(N__17234),
            .I(N__17229));
    InMux I__3706 (
            .O(N__17233),
            .I(N__17226));
    InMux I__3705 (
            .O(N__17232),
            .I(N__17223));
    Odrv4 I__3704 (
            .O(N__17229),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__3703 (
            .O(N__17226),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__3702 (
            .O(N__17223),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    InMux I__3701 (
            .O(N__17216),
            .I(N__17213));
    LocalMux I__3700 (
            .O(N__17213),
            .I(N__17208));
    InMux I__3699 (
            .O(N__17212),
            .I(N__17205));
    InMux I__3698 (
            .O(N__17211),
            .I(N__17202));
    Odrv4 I__3697 (
            .O(N__17208),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__3696 (
            .O(N__17205),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__3695 (
            .O(N__17202),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    CEMux I__3694 (
            .O(N__17195),
            .I(N__17180));
    CEMux I__3693 (
            .O(N__17194),
            .I(N__17180));
    CEMux I__3692 (
            .O(N__17193),
            .I(N__17180));
    CEMux I__3691 (
            .O(N__17192),
            .I(N__17180));
    CEMux I__3690 (
            .O(N__17191),
            .I(N__17180));
    GlobalMux I__3689 (
            .O(N__17180),
            .I(N__17177));
    gio2CtrlBuf I__3688 (
            .O(N__17177),
            .I(\delay_measurement_inst.delay_tr_timer.N_255_i_g ));
    InMux I__3687 (
            .O(N__17174),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    InMux I__3686 (
            .O(N__17171),
            .I(bfn_9_23_0_));
    InMux I__3685 (
            .O(N__17168),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    InMux I__3684 (
            .O(N__17165),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    InMux I__3683 (
            .O(N__17162),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    InMux I__3682 (
            .O(N__17159),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    InMux I__3681 (
            .O(N__17156),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    InMux I__3680 (
            .O(N__17153),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    InMux I__3679 (
            .O(N__17150),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    InMux I__3678 (
            .O(N__17147),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    InMux I__3677 (
            .O(N__17144),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    InMux I__3676 (
            .O(N__17141),
            .I(bfn_9_22_0_));
    InMux I__3675 (
            .O(N__17138),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    InMux I__3674 (
            .O(N__17135),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    InMux I__3673 (
            .O(N__17132),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    InMux I__3672 (
            .O(N__17129),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    InMux I__3671 (
            .O(N__17126),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    InMux I__3670 (
            .O(N__17123),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    InMux I__3669 (
            .O(N__17120),
            .I(N__17117));
    LocalMux I__3668 (
            .O(N__17117),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3 ));
    CascadeMux I__3667 (
            .O(N__17114),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_9_cascade_ ));
    InMux I__3666 (
            .O(N__17111),
            .I(N__17107));
    InMux I__3665 (
            .O(N__17110),
            .I(N__17104));
    LocalMux I__3664 (
            .O(N__17107),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_0_6 ));
    LocalMux I__3663 (
            .O(N__17104),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_0_6 ));
    InMux I__3662 (
            .O(N__17099),
            .I(N__17096));
    LocalMux I__3661 (
            .O(N__17096),
            .I(N__17093));
    Span4Mux_h I__3660 (
            .O(N__17093),
            .I(N__17089));
    InMux I__3659 (
            .O(N__17092),
            .I(N__17086));
    Span4Mux_h I__3658 (
            .O(N__17089),
            .I(N__17082));
    LocalMux I__3657 (
            .O(N__17086),
            .I(N__17079));
    InMux I__3656 (
            .O(N__17085),
            .I(N__17076));
    Odrv4 I__3655 (
            .O(N__17082),
            .I(\phase_controller_inst1.stoper_tr.N_97 ));
    Odrv12 I__3654 (
            .O(N__17079),
            .I(\phase_controller_inst1.stoper_tr.N_97 ));
    LocalMux I__3653 (
            .O(N__17076),
            .I(\phase_controller_inst1.stoper_tr.N_97 ));
    InMux I__3652 (
            .O(N__17069),
            .I(N__17065));
    InMux I__3651 (
            .O(N__17068),
            .I(N__17062));
    LocalMux I__3650 (
            .O(N__17065),
            .I(N__17058));
    LocalMux I__3649 (
            .O(N__17062),
            .I(N__17055));
    InMux I__3648 (
            .O(N__17061),
            .I(N__17052));
    Span12Mux_s9_h I__3647 (
            .O(N__17058),
            .I(N__17049));
    Span4Mux_h I__3646 (
            .O(N__17055),
            .I(N__17044));
    LocalMux I__3645 (
            .O(N__17052),
            .I(N__17044));
    Odrv12 I__3644 (
            .O(N__17049),
            .I(measured_delay_tr_4));
    Odrv4 I__3643 (
            .O(N__17044),
            .I(measured_delay_tr_4));
    InMux I__3642 (
            .O(N__17039),
            .I(N__17035));
    InMux I__3641 (
            .O(N__17038),
            .I(N__17032));
    LocalMux I__3640 (
            .O(N__17035),
            .I(N__17026));
    LocalMux I__3639 (
            .O(N__17032),
            .I(N__17026));
    InMux I__3638 (
            .O(N__17031),
            .I(N__17023));
    Span4Mux_v I__3637 (
            .O(N__17026),
            .I(N__17017));
    LocalMux I__3636 (
            .O(N__17023),
            .I(N__17017));
    InMux I__3635 (
            .O(N__17022),
            .I(N__17013));
    Span4Mux_h I__3634 (
            .O(N__17017),
            .I(N__17010));
    InMux I__3633 (
            .O(N__17016),
            .I(N__17007));
    LocalMux I__3632 (
            .O(N__17013),
            .I(measured_delay_tr_14));
    Odrv4 I__3631 (
            .O(N__17010),
            .I(measured_delay_tr_14));
    LocalMux I__3630 (
            .O(N__17007),
            .I(measured_delay_tr_14));
    InMux I__3629 (
            .O(N__17000),
            .I(N__16987));
    InMux I__3628 (
            .O(N__16999),
            .I(N__16987));
    InMux I__3627 (
            .O(N__16998),
            .I(N__16987));
    InMux I__3626 (
            .O(N__16997),
            .I(N__16984));
    InMux I__3625 (
            .O(N__16996),
            .I(N__16979));
    InMux I__3624 (
            .O(N__16995),
            .I(N__16979));
    InMux I__3623 (
            .O(N__16994),
            .I(N__16976));
    LocalMux I__3622 (
            .O(N__16987),
            .I(N__16973));
    LocalMux I__3621 (
            .O(N__16984),
            .I(N__16966));
    LocalMux I__3620 (
            .O(N__16979),
            .I(N__16966));
    LocalMux I__3619 (
            .O(N__16976),
            .I(N__16966));
    Span4Mux_v I__3618 (
            .O(N__16973),
            .I(N__16960));
    Span4Mux_v I__3617 (
            .O(N__16966),
            .I(N__16957));
    InMux I__3616 (
            .O(N__16965),
            .I(N__16952));
    InMux I__3615 (
            .O(N__16964),
            .I(N__16952));
    CascadeMux I__3614 (
            .O(N__16963),
            .I(N__16949));
    Span4Mux_h I__3613 (
            .O(N__16960),
            .I(N__16942));
    Span4Mux_h I__3612 (
            .O(N__16957),
            .I(N__16942));
    LocalMux I__3611 (
            .O(N__16952),
            .I(N__16942));
    InMux I__3610 (
            .O(N__16949),
            .I(N__16939));
    Sp12to4 I__3609 (
            .O(N__16942),
            .I(N__16934));
    LocalMux I__3608 (
            .O(N__16939),
            .I(N__16934));
    Odrv12 I__3607 (
            .O(N__16934),
            .I(measured_delay_tr_15));
    InMux I__3606 (
            .O(N__16931),
            .I(N__16928));
    LocalMux I__3605 (
            .O(N__16928),
            .I(N__16924));
    InMux I__3604 (
            .O(N__16927),
            .I(N__16921));
    Span4Mux_v I__3603 (
            .O(N__16924),
            .I(N__16915));
    LocalMux I__3602 (
            .O(N__16921),
            .I(N__16915));
    InMux I__3601 (
            .O(N__16920),
            .I(N__16912));
    Span4Mux_h I__3600 (
            .O(N__16915),
            .I(N__16907));
    LocalMux I__3599 (
            .O(N__16912),
            .I(N__16907));
    Odrv4 I__3598 (
            .O(N__16907),
            .I(measured_delay_tr_5));
    InMux I__3597 (
            .O(N__16904),
            .I(N__16901));
    LocalMux I__3596 (
            .O(N__16901),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3 ));
    InMux I__3595 (
            .O(N__16898),
            .I(N__16895));
    LocalMux I__3594 (
            .O(N__16895),
            .I(N__16892));
    Span4Mux_h I__3593 (
            .O(N__16892),
            .I(N__16886));
    CascadeMux I__3592 (
            .O(N__16891),
            .I(N__16883));
    CascadeMux I__3591 (
            .O(N__16890),
            .I(N__16880));
    InMux I__3590 (
            .O(N__16889),
            .I(N__16877));
    Span4Mux_v I__3589 (
            .O(N__16886),
            .I(N__16874));
    InMux I__3588 (
            .O(N__16883),
            .I(N__16869));
    InMux I__3587 (
            .O(N__16880),
            .I(N__16869));
    LocalMux I__3586 (
            .O(N__16877),
            .I(N__16866));
    Odrv4 I__3585 (
            .O(N__16874),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    LocalMux I__3584 (
            .O(N__16869),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    Odrv4 I__3583 (
            .O(N__16866),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    IoInMux I__3582 (
            .O(N__16859),
            .I(N__16856));
    LocalMux I__3581 (
            .O(N__16856),
            .I(N__16853));
    Span4Mux_s2_v I__3580 (
            .O(N__16853),
            .I(N__16850));
    Span4Mux_h I__3579 (
            .O(N__16850),
            .I(N__16847));
    Span4Mux_v I__3578 (
            .O(N__16847),
            .I(N__16844));
    Span4Mux_v I__3577 (
            .O(N__16844),
            .I(N__16841));
    Odrv4 I__3576 (
            .O(N__16841),
            .I(s1_phy_c));
    InMux I__3575 (
            .O(N__16838),
            .I(bfn_9_21_0_));
    InMux I__3574 (
            .O(N__16835),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    InMux I__3573 (
            .O(N__16832),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    InMux I__3572 (
            .O(N__16829),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    InMux I__3571 (
            .O(N__16826),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    InMux I__3570 (
            .O(N__16823),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    InMux I__3569 (
            .O(N__16820),
            .I(N__16816));
    InMux I__3568 (
            .O(N__16819),
            .I(N__16813));
    LocalMux I__3567 (
            .O(N__16816),
            .I(N__16808));
    LocalMux I__3566 (
            .O(N__16813),
            .I(N__16808));
    Span4Mux_v I__3565 (
            .O(N__16808),
            .I(N__16804));
    InMux I__3564 (
            .O(N__16807),
            .I(N__16801));
    Span4Mux_h I__3563 (
            .O(N__16804),
            .I(N__16796));
    LocalMux I__3562 (
            .O(N__16801),
            .I(N__16796));
    Odrv4 I__3561 (
            .O(N__16796),
            .I(measured_delay_tr_6));
    InMux I__3560 (
            .O(N__16793),
            .I(N__16789));
    InMux I__3559 (
            .O(N__16792),
            .I(N__16786));
    LocalMux I__3558 (
            .O(N__16789),
            .I(N__16783));
    LocalMux I__3557 (
            .O(N__16786),
            .I(N__16779));
    Span4Mux_h I__3556 (
            .O(N__16783),
            .I(N__16775));
    InMux I__3555 (
            .O(N__16782),
            .I(N__16772));
    Span4Mux_h I__3554 (
            .O(N__16779),
            .I(N__16769));
    InMux I__3553 (
            .O(N__16778),
            .I(N__16766));
    Span4Mux_h I__3552 (
            .O(N__16775),
            .I(N__16761));
    LocalMux I__3551 (
            .O(N__16772),
            .I(N__16761));
    Odrv4 I__3550 (
            .O(N__16769),
            .I(measured_delay_tr_18));
    LocalMux I__3549 (
            .O(N__16766),
            .I(measured_delay_tr_18));
    Odrv4 I__3548 (
            .O(N__16761),
            .I(measured_delay_tr_18));
    InMux I__3547 (
            .O(N__16754),
            .I(N__16751));
    LocalMux I__3546 (
            .O(N__16751),
            .I(N__16747));
    InMux I__3545 (
            .O(N__16750),
            .I(N__16744));
    Span4Mux_h I__3544 (
            .O(N__16747),
            .I(N__16741));
    LocalMux I__3543 (
            .O(N__16744),
            .I(N__16738));
    Span4Mux_h I__3542 (
            .O(N__16741),
            .I(N__16733));
    Span4Mux_h I__3541 (
            .O(N__16738),
            .I(N__16730));
    InMux I__3540 (
            .O(N__16737),
            .I(N__16727));
    InMux I__3539 (
            .O(N__16736),
            .I(N__16724));
    Odrv4 I__3538 (
            .O(N__16733),
            .I(measured_delay_tr_17));
    Odrv4 I__3537 (
            .O(N__16730),
            .I(measured_delay_tr_17));
    LocalMux I__3536 (
            .O(N__16727),
            .I(measured_delay_tr_17));
    LocalMux I__3535 (
            .O(N__16724),
            .I(measured_delay_tr_17));
    InMux I__3534 (
            .O(N__16715),
            .I(N__16712));
    LocalMux I__3533 (
            .O(N__16712),
            .I(N__16708));
    InMux I__3532 (
            .O(N__16711),
            .I(N__16705));
    Span4Mux_v I__3531 (
            .O(N__16708),
            .I(N__16702));
    LocalMux I__3530 (
            .O(N__16705),
            .I(N__16699));
    Span4Mux_h I__3529 (
            .O(N__16702),
            .I(N__16694));
    Span4Mux_v I__3528 (
            .O(N__16699),
            .I(N__16691));
    InMux I__3527 (
            .O(N__16698),
            .I(N__16688));
    InMux I__3526 (
            .O(N__16697),
            .I(N__16685));
    Odrv4 I__3525 (
            .O(N__16694),
            .I(measured_delay_tr_16));
    Odrv4 I__3524 (
            .O(N__16691),
            .I(measured_delay_tr_16));
    LocalMux I__3523 (
            .O(N__16688),
            .I(measured_delay_tr_16));
    LocalMux I__3522 (
            .O(N__16685),
            .I(measured_delay_tr_16));
    InMux I__3521 (
            .O(N__16676),
            .I(N__16673));
    LocalMux I__3520 (
            .O(N__16673),
            .I(N__16669));
    InMux I__3519 (
            .O(N__16672),
            .I(N__16666));
    Span12Mux_v I__3518 (
            .O(N__16669),
            .I(N__16660));
    LocalMux I__3517 (
            .O(N__16666),
            .I(N__16660));
    InMux I__3516 (
            .O(N__16665),
            .I(N__16657));
    Odrv12 I__3515 (
            .O(N__16660),
            .I(measured_delay_tr_12));
    LocalMux I__3514 (
            .O(N__16657),
            .I(measured_delay_tr_12));
    InMux I__3513 (
            .O(N__16652),
            .I(N__16649));
    LocalMux I__3512 (
            .O(N__16649),
            .I(N__16646));
    Span4Mux_h I__3511 (
            .O(N__16646),
            .I(N__16642));
    InMux I__3510 (
            .O(N__16645),
            .I(N__16639));
    Span4Mux_h I__3509 (
            .O(N__16642),
            .I(N__16635));
    LocalMux I__3508 (
            .O(N__16639),
            .I(N__16632));
    InMux I__3507 (
            .O(N__16638),
            .I(N__16629));
    Odrv4 I__3506 (
            .O(N__16635),
            .I(measured_delay_tr_11));
    Odrv12 I__3505 (
            .O(N__16632),
            .I(measured_delay_tr_11));
    LocalMux I__3504 (
            .O(N__16629),
            .I(measured_delay_tr_11));
    InMux I__3503 (
            .O(N__16622),
            .I(N__16619));
    LocalMux I__3502 (
            .O(N__16619),
            .I(N__16615));
    InMux I__3501 (
            .O(N__16618),
            .I(N__16612));
    Span4Mux_h I__3500 (
            .O(N__16615),
            .I(N__16606));
    LocalMux I__3499 (
            .O(N__16612),
            .I(N__16606));
    CascadeMux I__3498 (
            .O(N__16611),
            .I(N__16603));
    Span4Mux_h I__3497 (
            .O(N__16606),
            .I(N__16600));
    InMux I__3496 (
            .O(N__16603),
            .I(N__16597));
    Odrv4 I__3495 (
            .O(N__16600),
            .I(measured_delay_tr_13));
    LocalMux I__3494 (
            .O(N__16597),
            .I(measured_delay_tr_13));
    InMux I__3493 (
            .O(N__16592),
            .I(N__16589));
    LocalMux I__3492 (
            .O(N__16589),
            .I(N__16585));
    InMux I__3491 (
            .O(N__16588),
            .I(N__16582));
    Span4Mux_h I__3490 (
            .O(N__16585),
            .I(N__16577));
    LocalMux I__3489 (
            .O(N__16582),
            .I(N__16577));
    Span4Mux_h I__3488 (
            .O(N__16577),
            .I(N__16573));
    InMux I__3487 (
            .O(N__16576),
            .I(N__16570));
    Odrv4 I__3486 (
            .O(N__16573),
            .I(measured_delay_tr_10));
    LocalMux I__3485 (
            .O(N__16570),
            .I(measured_delay_tr_10));
    CascadeMux I__3484 (
            .O(N__16565),
            .I(N__16561));
    InMux I__3483 (
            .O(N__16564),
            .I(N__16558));
    InMux I__3482 (
            .O(N__16561),
            .I(N__16555));
    LocalMux I__3481 (
            .O(N__16558),
            .I(N__16552));
    LocalMux I__3480 (
            .O(N__16555),
            .I(N__16549));
    Span4Mux_h I__3479 (
            .O(N__16552),
            .I(N__16543));
    Span4Mux_v I__3478 (
            .O(N__16549),
            .I(N__16543));
    InMux I__3477 (
            .O(N__16548),
            .I(N__16540));
    Span4Mux_h I__3476 (
            .O(N__16543),
            .I(N__16535));
    LocalMux I__3475 (
            .O(N__16540),
            .I(N__16535));
    Odrv4 I__3474 (
            .O(N__16535),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_0_6 ));
    CascadeMux I__3473 (
            .O(N__16532),
            .I(N__16528));
    InMux I__3472 (
            .O(N__16531),
            .I(N__16525));
    InMux I__3471 (
            .O(N__16528),
            .I(N__16522));
    LocalMux I__3470 (
            .O(N__16525),
            .I(N__16519));
    LocalMux I__3469 (
            .O(N__16522),
            .I(N__16516));
    Span4Mux_v I__3468 (
            .O(N__16519),
            .I(N__16510));
    Span4Mux_h I__3467 (
            .O(N__16516),
            .I(N__16510));
    InMux I__3466 (
            .O(N__16515),
            .I(N__16507));
    Span4Mux_h I__3465 (
            .O(N__16510),
            .I(N__16504));
    LocalMux I__3464 (
            .O(N__16507),
            .I(N__16501));
    Odrv4 I__3463 (
            .O(N__16504),
            .I(measured_delay_tr_9));
    Odrv4 I__3462 (
            .O(N__16501),
            .I(measured_delay_tr_9));
    CascadeMux I__3461 (
            .O(N__16496),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_0_6_cascade_ ));
    InMux I__3460 (
            .O(N__16493),
            .I(N__16490));
    LocalMux I__3459 (
            .O(N__16490),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_9 ));
    CascadeMux I__3458 (
            .O(N__16487),
            .I(N__16484));
    InMux I__3457 (
            .O(N__16484),
            .I(N__16480));
    CascadeMux I__3456 (
            .O(N__16483),
            .I(N__16477));
    LocalMux I__3455 (
            .O(N__16480),
            .I(N__16474));
    InMux I__3454 (
            .O(N__16477),
            .I(N__16471));
    Span4Mux_v I__3453 (
            .O(N__16474),
            .I(N__16466));
    LocalMux I__3452 (
            .O(N__16471),
            .I(N__16466));
    Span4Mux_h I__3451 (
            .O(N__16466),
            .I(N__16463));
    Odrv4 I__3450 (
            .O(N__16463),
            .I(measured_delay_tr_1));
    CascadeMux I__3449 (
            .O(N__16460),
            .I(N__16457));
    InMux I__3448 (
            .O(N__16457),
            .I(N__16453));
    InMux I__3447 (
            .O(N__16456),
            .I(N__16450));
    LocalMux I__3446 (
            .O(N__16453),
            .I(N__16446));
    LocalMux I__3445 (
            .O(N__16450),
            .I(N__16443));
    InMux I__3444 (
            .O(N__16449),
            .I(N__16440));
    Span4Mux_h I__3443 (
            .O(N__16446),
            .I(N__16437));
    Span4Mux_h I__3442 (
            .O(N__16443),
            .I(N__16432));
    LocalMux I__3441 (
            .O(N__16440),
            .I(N__16432));
    Span4Mux_h I__3440 (
            .O(N__16437),
            .I(N__16429));
    Span4Mux_h I__3439 (
            .O(N__16432),
            .I(N__16426));
    Odrv4 I__3438 (
            .O(N__16429),
            .I(measured_delay_tr_2));
    Odrv4 I__3437 (
            .O(N__16426),
            .I(measured_delay_tr_2));
    CascadeMux I__3436 (
            .O(N__16421),
            .I(N__16417));
    CascadeMux I__3435 (
            .O(N__16420),
            .I(N__16414));
    InMux I__3434 (
            .O(N__16417),
            .I(N__16411));
    InMux I__3433 (
            .O(N__16414),
            .I(N__16408));
    LocalMux I__3432 (
            .O(N__16411),
            .I(N__16405));
    LocalMux I__3431 (
            .O(N__16408),
            .I(N__16402));
    Span4Mux_h I__3430 (
            .O(N__16405),
            .I(N__16398));
    Span4Mux_h I__3429 (
            .O(N__16402),
            .I(N__16395));
    InMux I__3428 (
            .O(N__16401),
            .I(N__16392));
    Span4Mux_h I__3427 (
            .O(N__16398),
            .I(N__16389));
    Span4Mux_h I__3426 (
            .O(N__16395),
            .I(N__16386));
    LocalMux I__3425 (
            .O(N__16392),
            .I(N__16383));
    Odrv4 I__3424 (
            .O(N__16389),
            .I(measured_delay_tr_3));
    Odrv4 I__3423 (
            .O(N__16386),
            .I(measured_delay_tr_3));
    Odrv4 I__3422 (
            .O(N__16383),
            .I(measured_delay_tr_3));
    CascadeMux I__3421 (
            .O(N__16376),
            .I(N__16371));
    CascadeMux I__3420 (
            .O(N__16375),
            .I(N__16368));
    InMux I__3419 (
            .O(N__16374),
            .I(N__16365));
    InMux I__3418 (
            .O(N__16371),
            .I(N__16360));
    InMux I__3417 (
            .O(N__16368),
            .I(N__16360));
    LocalMux I__3416 (
            .O(N__16365),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__3415 (
            .O(N__16360),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__3414 (
            .O(N__16355),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__3413 (
            .O(N__16352),
            .I(N__16347));
    CascadeMux I__3412 (
            .O(N__16351),
            .I(N__16344));
    InMux I__3411 (
            .O(N__16350),
            .I(N__16341));
    InMux I__3410 (
            .O(N__16347),
            .I(N__16336));
    InMux I__3409 (
            .O(N__16344),
            .I(N__16336));
    LocalMux I__3408 (
            .O(N__16341),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__3407 (
            .O(N__16336),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__3406 (
            .O(N__16331),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__3405 (
            .O(N__16328),
            .I(N__16323));
    InMux I__3404 (
            .O(N__16327),
            .I(N__16320));
    InMux I__3403 (
            .O(N__16326),
            .I(N__16317));
    LocalMux I__3402 (
            .O(N__16323),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__3401 (
            .O(N__16320),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__3400 (
            .O(N__16317),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__3399 (
            .O(N__16310),
            .I(bfn_9_16_0_));
    InMux I__3398 (
            .O(N__16307),
            .I(N__16302));
    InMux I__3397 (
            .O(N__16306),
            .I(N__16299));
    InMux I__3396 (
            .O(N__16305),
            .I(N__16296));
    LocalMux I__3395 (
            .O(N__16302),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__3394 (
            .O(N__16299),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__3393 (
            .O(N__16296),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    InMux I__3392 (
            .O(N__16289),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__3391 (
            .O(N__16286),
            .I(N__16282));
    InMux I__3390 (
            .O(N__16285),
            .I(N__16279));
    LocalMux I__3389 (
            .O(N__16282),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    LocalMux I__3388 (
            .O(N__16279),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    CascadeMux I__3387 (
            .O(N__16274),
            .I(N__16269));
    CascadeMux I__3386 (
            .O(N__16273),
            .I(N__16266));
    InMux I__3385 (
            .O(N__16272),
            .I(N__16263));
    InMux I__3384 (
            .O(N__16269),
            .I(N__16258));
    InMux I__3383 (
            .O(N__16266),
            .I(N__16258));
    LocalMux I__3382 (
            .O(N__16263),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    LocalMux I__3381 (
            .O(N__16258),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    InMux I__3380 (
            .O(N__16253),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__3379 (
            .O(N__16250),
            .I(N__16246));
    InMux I__3378 (
            .O(N__16249),
            .I(N__16243));
    LocalMux I__3377 (
            .O(N__16246),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    LocalMux I__3376 (
            .O(N__16243),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CascadeMux I__3375 (
            .O(N__16238),
            .I(N__16233));
    CascadeMux I__3374 (
            .O(N__16237),
            .I(N__16230));
    InMux I__3373 (
            .O(N__16236),
            .I(N__16227));
    InMux I__3372 (
            .O(N__16233),
            .I(N__16222));
    InMux I__3371 (
            .O(N__16230),
            .I(N__16222));
    LocalMux I__3370 (
            .O(N__16227),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    LocalMux I__3369 (
            .O(N__16222),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__3368 (
            .O(N__16217),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__3367 (
            .O(N__16214),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    CascadeMux I__3366 (
            .O(N__16211),
            .I(N__16206));
    CascadeMux I__3365 (
            .O(N__16210),
            .I(N__16203));
    InMux I__3364 (
            .O(N__16209),
            .I(N__16200));
    InMux I__3363 (
            .O(N__16206),
            .I(N__16195));
    InMux I__3362 (
            .O(N__16203),
            .I(N__16195));
    LocalMux I__3361 (
            .O(N__16200),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__3360 (
            .O(N__16195),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__3359 (
            .O(N__16190),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__3358 (
            .O(N__16187),
            .I(N__16182));
    CascadeMux I__3357 (
            .O(N__16186),
            .I(N__16179));
    InMux I__3356 (
            .O(N__16185),
            .I(N__16176));
    InMux I__3355 (
            .O(N__16182),
            .I(N__16171));
    InMux I__3354 (
            .O(N__16179),
            .I(N__16171));
    LocalMux I__3353 (
            .O(N__16176),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__3352 (
            .O(N__16171),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__3351 (
            .O(N__16166),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__3350 (
            .O(N__16163),
            .I(N__16158));
    InMux I__3349 (
            .O(N__16162),
            .I(N__16155));
    InMux I__3348 (
            .O(N__16161),
            .I(N__16152));
    LocalMux I__3347 (
            .O(N__16158),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__3346 (
            .O(N__16155),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__3345 (
            .O(N__16152),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__3344 (
            .O(N__16145),
            .I(bfn_9_15_0_));
    InMux I__3343 (
            .O(N__16142),
            .I(N__16137));
    InMux I__3342 (
            .O(N__16141),
            .I(N__16134));
    InMux I__3341 (
            .O(N__16140),
            .I(N__16131));
    LocalMux I__3340 (
            .O(N__16137),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__3339 (
            .O(N__16134),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__3338 (
            .O(N__16131),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__3337 (
            .O(N__16124),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__3336 (
            .O(N__16121),
            .I(N__16116));
    CascadeMux I__3335 (
            .O(N__16120),
            .I(N__16113));
    InMux I__3334 (
            .O(N__16119),
            .I(N__16110));
    InMux I__3333 (
            .O(N__16116),
            .I(N__16105));
    InMux I__3332 (
            .O(N__16113),
            .I(N__16105));
    LocalMux I__3331 (
            .O(N__16110),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    LocalMux I__3330 (
            .O(N__16105),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__3329 (
            .O(N__16100),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__3328 (
            .O(N__16097),
            .I(N__16092));
    CascadeMux I__3327 (
            .O(N__16096),
            .I(N__16089));
    InMux I__3326 (
            .O(N__16095),
            .I(N__16086));
    InMux I__3325 (
            .O(N__16092),
            .I(N__16081));
    InMux I__3324 (
            .O(N__16089),
            .I(N__16081));
    LocalMux I__3323 (
            .O(N__16086),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    LocalMux I__3322 (
            .O(N__16081),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__3321 (
            .O(N__16076),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__3320 (
            .O(N__16073),
            .I(N__16068));
    InMux I__3319 (
            .O(N__16072),
            .I(N__16063));
    InMux I__3318 (
            .O(N__16071),
            .I(N__16063));
    LocalMux I__3317 (
            .O(N__16068),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    LocalMux I__3316 (
            .O(N__16063),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__3315 (
            .O(N__16058),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__3314 (
            .O(N__16055),
            .I(N__16050));
    InMux I__3313 (
            .O(N__16054),
            .I(N__16045));
    InMux I__3312 (
            .O(N__16053),
            .I(N__16045));
    LocalMux I__3311 (
            .O(N__16050),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__3310 (
            .O(N__16045),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__3309 (
            .O(N__16040),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__3308 (
            .O(N__16037),
            .I(N__16032));
    InMux I__3307 (
            .O(N__16036),
            .I(N__16027));
    InMux I__3306 (
            .O(N__16035),
            .I(N__16027));
    LocalMux I__3305 (
            .O(N__16032),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__3304 (
            .O(N__16027),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__3303 (
            .O(N__16022),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__3302 (
            .O(N__16019),
            .I(N__16014));
    CascadeMux I__3301 (
            .O(N__16018),
            .I(N__16011));
    InMux I__3300 (
            .O(N__16017),
            .I(N__16008));
    InMux I__3299 (
            .O(N__16014),
            .I(N__16003));
    InMux I__3298 (
            .O(N__16011),
            .I(N__16003));
    LocalMux I__3297 (
            .O(N__16008),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__3296 (
            .O(N__16003),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__3295 (
            .O(N__15998),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__3294 (
            .O(N__15995),
            .I(N__15990));
    CascadeMux I__3293 (
            .O(N__15994),
            .I(N__15987));
    InMux I__3292 (
            .O(N__15993),
            .I(N__15984));
    InMux I__3291 (
            .O(N__15990),
            .I(N__15979));
    InMux I__3290 (
            .O(N__15987),
            .I(N__15979));
    LocalMux I__3289 (
            .O(N__15984),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__3288 (
            .O(N__15979),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__3287 (
            .O(N__15974),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__3286 (
            .O(N__15971),
            .I(N__15966));
    InMux I__3285 (
            .O(N__15970),
            .I(N__15963));
    InMux I__3284 (
            .O(N__15969),
            .I(N__15960));
    LocalMux I__3283 (
            .O(N__15966),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__3282 (
            .O(N__15963),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__3281 (
            .O(N__15960),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__3280 (
            .O(N__15953),
            .I(bfn_9_14_0_));
    InMux I__3279 (
            .O(N__15950),
            .I(N__15945));
    InMux I__3278 (
            .O(N__15949),
            .I(N__15942));
    InMux I__3277 (
            .O(N__15948),
            .I(N__15939));
    LocalMux I__3276 (
            .O(N__15945),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__3275 (
            .O(N__15942),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__3274 (
            .O(N__15939),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__3273 (
            .O(N__15932),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__3272 (
            .O(N__15929),
            .I(N__15924));
    CascadeMux I__3271 (
            .O(N__15928),
            .I(N__15921));
    InMux I__3270 (
            .O(N__15927),
            .I(N__15918));
    InMux I__3269 (
            .O(N__15924),
            .I(N__15913));
    InMux I__3268 (
            .O(N__15921),
            .I(N__15913));
    LocalMux I__3267 (
            .O(N__15918),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    LocalMux I__3266 (
            .O(N__15913),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__3265 (
            .O(N__15908),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__3264 (
            .O(N__15905),
            .I(N__15900));
    CascadeMux I__3263 (
            .O(N__15904),
            .I(N__15897));
    InMux I__3262 (
            .O(N__15903),
            .I(N__15894));
    InMux I__3261 (
            .O(N__15900),
            .I(N__15889));
    InMux I__3260 (
            .O(N__15897),
            .I(N__15889));
    LocalMux I__3259 (
            .O(N__15894),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    LocalMux I__3258 (
            .O(N__15889),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__3257 (
            .O(N__15884),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__3256 (
            .O(N__15881),
            .I(N__15876));
    InMux I__3255 (
            .O(N__15880),
            .I(N__15871));
    InMux I__3254 (
            .O(N__15879),
            .I(N__15871));
    LocalMux I__3253 (
            .O(N__15876),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    LocalMux I__3252 (
            .O(N__15871),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__3251 (
            .O(N__15866),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__3250 (
            .O(N__15863),
            .I(N__15858));
    InMux I__3249 (
            .O(N__15862),
            .I(N__15853));
    InMux I__3248 (
            .O(N__15861),
            .I(N__15853));
    LocalMux I__3247 (
            .O(N__15858),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__3246 (
            .O(N__15853),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__3245 (
            .O(N__15848),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__3244 (
            .O(N__15845),
            .I(N__15836));
    InMux I__3243 (
            .O(N__15844),
            .I(N__15836));
    InMux I__3242 (
            .O(N__15843),
            .I(N__15836));
    LocalMux I__3241 (
            .O(N__15836),
            .I(\delay_measurement_inst.N_243 ));
    InMux I__3240 (
            .O(N__15833),
            .I(N__15816));
    InMux I__3239 (
            .O(N__15832),
            .I(N__15816));
    InMux I__3238 (
            .O(N__15831),
            .I(N__15816));
    InMux I__3237 (
            .O(N__15830),
            .I(N__15816));
    InMux I__3236 (
            .O(N__15829),
            .I(N__15816));
    InMux I__3235 (
            .O(N__15828),
            .I(N__15813));
    InMux I__3234 (
            .O(N__15827),
            .I(N__15810));
    LocalMux I__3233 (
            .O(N__15816),
            .I(\delay_measurement_inst.N_247 ));
    LocalMux I__3232 (
            .O(N__15813),
            .I(\delay_measurement_inst.N_247 ));
    LocalMux I__3231 (
            .O(N__15810),
            .I(\delay_measurement_inst.N_247 ));
    InMux I__3230 (
            .O(N__15803),
            .I(N__15791));
    InMux I__3229 (
            .O(N__15802),
            .I(N__15791));
    InMux I__3228 (
            .O(N__15801),
            .I(N__15791));
    InMux I__3227 (
            .O(N__15800),
            .I(N__15786));
    InMux I__3226 (
            .O(N__15799),
            .I(N__15786));
    InMux I__3225 (
            .O(N__15798),
            .I(N__15783));
    LocalMux I__3224 (
            .O(N__15791),
            .I(\delay_measurement_inst.N_216_1 ));
    LocalMux I__3223 (
            .O(N__15786),
            .I(\delay_measurement_inst.N_216_1 ));
    LocalMux I__3222 (
            .O(N__15783),
            .I(\delay_measurement_inst.N_216_1 ));
    InMux I__3221 (
            .O(N__15776),
            .I(N__15773));
    LocalMux I__3220 (
            .O(N__15773),
            .I(N__15768));
    InMux I__3219 (
            .O(N__15772),
            .I(N__15765));
    CascadeMux I__3218 (
            .O(N__15771),
            .I(N__15762));
    Span4Mux_v I__3217 (
            .O(N__15768),
            .I(N__15759));
    LocalMux I__3216 (
            .O(N__15765),
            .I(N__15756));
    InMux I__3215 (
            .O(N__15762),
            .I(N__15753));
    Span4Mux_v I__3214 (
            .O(N__15759),
            .I(N__15746));
    Span4Mux_v I__3213 (
            .O(N__15756),
            .I(N__15746));
    LocalMux I__3212 (
            .O(N__15753),
            .I(N__15746));
    Span4Mux_h I__3211 (
            .O(N__15746),
            .I(N__15743));
    Odrv4 I__3210 (
            .O(N__15743),
            .I(measured_delay_hc_13));
    CEMux I__3209 (
            .O(N__15740),
            .I(N__15736));
    CEMux I__3208 (
            .O(N__15739),
            .I(N__15733));
    LocalMux I__3207 (
            .O(N__15736),
            .I(N__15729));
    LocalMux I__3206 (
            .O(N__15733),
            .I(N__15726));
    CEMux I__3205 (
            .O(N__15732),
            .I(N__15723));
    Span4Mux_v I__3204 (
            .O(N__15729),
            .I(N__15720));
    Span4Mux_h I__3203 (
            .O(N__15726),
            .I(N__15717));
    LocalMux I__3202 (
            .O(N__15723),
            .I(N__15714));
    Odrv4 I__3201 (
            .O(N__15720),
            .I(\delay_measurement_inst.un3_elapsed_time_hc_0_i_0 ));
    Odrv4 I__3200 (
            .O(N__15717),
            .I(\delay_measurement_inst.un3_elapsed_time_hc_0_i_0 ));
    Odrv4 I__3199 (
            .O(N__15714),
            .I(\delay_measurement_inst.un3_elapsed_time_hc_0_i_0 ));
    CascadeMux I__3198 (
            .O(N__15707),
            .I(N__15703));
    InMux I__3197 (
            .O(N__15706),
            .I(N__15700));
    InMux I__3196 (
            .O(N__15703),
            .I(N__15696));
    LocalMux I__3195 (
            .O(N__15700),
            .I(N__15692));
    InMux I__3194 (
            .O(N__15699),
            .I(N__15689));
    LocalMux I__3193 (
            .O(N__15696),
            .I(N__15686));
    InMux I__3192 (
            .O(N__15695),
            .I(N__15683));
    Span4Mux_h I__3191 (
            .O(N__15692),
            .I(N__15678));
    LocalMux I__3190 (
            .O(N__15689),
            .I(N__15678));
    Odrv4 I__3189 (
            .O(N__15686),
            .I(\phase_controller_slave.stateZ0Z_1 ));
    LocalMux I__3188 (
            .O(N__15683),
            .I(\phase_controller_slave.stateZ0Z_1 ));
    Odrv4 I__3187 (
            .O(N__15678),
            .I(\phase_controller_slave.stateZ0Z_1 ));
    IoInMux I__3186 (
            .O(N__15671),
            .I(N__15668));
    LocalMux I__3185 (
            .O(N__15668),
            .I(N__15665));
    Odrv12 I__3184 (
            .O(N__15665),
            .I(s4_phy_c));
    InMux I__3183 (
            .O(N__15662),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__3182 (
            .O(N__15659),
            .I(N__15654));
    CascadeMux I__3181 (
            .O(N__15658),
            .I(N__15651));
    InMux I__3180 (
            .O(N__15657),
            .I(N__15648));
    InMux I__3179 (
            .O(N__15654),
            .I(N__15643));
    InMux I__3178 (
            .O(N__15651),
            .I(N__15643));
    LocalMux I__3177 (
            .O(N__15648),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    LocalMux I__3176 (
            .O(N__15643),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__3175 (
            .O(N__15638),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__3174 (
            .O(N__15635),
            .I(N__15630));
    CascadeMux I__3173 (
            .O(N__15634),
            .I(N__15627));
    InMux I__3172 (
            .O(N__15633),
            .I(N__15624));
    InMux I__3171 (
            .O(N__15630),
            .I(N__15619));
    InMux I__3170 (
            .O(N__15627),
            .I(N__15619));
    LocalMux I__3169 (
            .O(N__15624),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    LocalMux I__3168 (
            .O(N__15619),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__3167 (
            .O(N__15614),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__3166 (
            .O(N__15611),
            .I(N__15606));
    InMux I__3165 (
            .O(N__15610),
            .I(N__15601));
    InMux I__3164 (
            .O(N__15609),
            .I(N__15601));
    LocalMux I__3163 (
            .O(N__15606),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    LocalMux I__3162 (
            .O(N__15601),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__3161 (
            .O(N__15596),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__3160 (
            .O(N__15593),
            .I(\delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_3_cascade_ ));
    InMux I__3159 (
            .O(N__15590),
            .I(N__15584));
    InMux I__3158 (
            .O(N__15589),
            .I(N__15584));
    LocalMux I__3157 (
            .O(N__15584),
            .I(\delay_measurement_inst.delay_hc_timer.N_232_4 ));
    InMux I__3156 (
            .O(N__15581),
            .I(N__15578));
    LocalMux I__3155 (
            .O(N__15578),
            .I(\delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_2 ));
    CascadeMux I__3154 (
            .O(N__15575),
            .I(\delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_6_cascade_ ));
    InMux I__3153 (
            .O(N__15572),
            .I(N__15569));
    LocalMux I__3152 (
            .O(N__15569),
            .I(\delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_0_7 ));
    InMux I__3151 (
            .O(N__15566),
            .I(N__15563));
    LocalMux I__3150 (
            .O(N__15563),
            .I(\delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_7 ));
    InMux I__3149 (
            .O(N__15560),
            .I(N__15554));
    InMux I__3148 (
            .O(N__15559),
            .I(N__15554));
    LocalMux I__3147 (
            .O(N__15554),
            .I(\delay_measurement_inst.un3_elapsed_time_hc_0_i ));
    CascadeMux I__3146 (
            .O(N__15551),
            .I(\delay_measurement_inst.un3_elapsed_time_hc_0_i_cascade_ ));
    InMux I__3145 (
            .O(N__15548),
            .I(N__15545));
    LocalMux I__3144 (
            .O(N__15545),
            .I(\delay_measurement_inst.N_219 ));
    CascadeMux I__3143 (
            .O(N__15542),
            .I(\delay_measurement_inst.delay_hc_timer.N_237_cascade_ ));
    CascadeMux I__3142 (
            .O(N__15539),
            .I(N__15534));
    InMux I__3141 (
            .O(N__15538),
            .I(N__15524));
    InMux I__3140 (
            .O(N__15537),
            .I(N__15524));
    InMux I__3139 (
            .O(N__15534),
            .I(N__15517));
    InMux I__3138 (
            .O(N__15533),
            .I(N__15517));
    InMux I__3137 (
            .O(N__15532),
            .I(N__15517));
    InMux I__3136 (
            .O(N__15531),
            .I(N__15512));
    InMux I__3135 (
            .O(N__15530),
            .I(N__15512));
    InMux I__3134 (
            .O(N__15529),
            .I(N__15509));
    LocalMux I__3133 (
            .O(N__15524),
            .I(\delay_measurement_inst.N_209 ));
    LocalMux I__3132 (
            .O(N__15517),
            .I(\delay_measurement_inst.N_209 ));
    LocalMux I__3131 (
            .O(N__15512),
            .I(\delay_measurement_inst.N_209 ));
    LocalMux I__3130 (
            .O(N__15509),
            .I(\delay_measurement_inst.N_209 ));
    InMux I__3129 (
            .O(N__15500),
            .I(N__15495));
    InMux I__3128 (
            .O(N__15499),
            .I(N__15492));
    InMux I__3127 (
            .O(N__15498),
            .I(N__15489));
    LocalMux I__3126 (
            .O(N__15495),
            .I(\delay_measurement_inst.N_207 ));
    LocalMux I__3125 (
            .O(N__15492),
            .I(\delay_measurement_inst.N_207 ));
    LocalMux I__3124 (
            .O(N__15489),
            .I(\delay_measurement_inst.N_207 ));
    CascadeMux I__3123 (
            .O(N__15482),
            .I(\delay_measurement_inst.N_207_cascade_ ));
    CascadeMux I__3122 (
            .O(N__15479),
            .I(N__15475));
    CascadeMux I__3121 (
            .O(N__15478),
            .I(N__15472));
    InMux I__3120 (
            .O(N__15475),
            .I(N__15463));
    InMux I__3119 (
            .O(N__15472),
            .I(N__15460));
    InMux I__3118 (
            .O(N__15471),
            .I(N__15440));
    InMux I__3117 (
            .O(N__15470),
            .I(N__15440));
    InMux I__3116 (
            .O(N__15469),
            .I(N__15440));
    InMux I__3115 (
            .O(N__15468),
            .I(N__15440));
    InMux I__3114 (
            .O(N__15467),
            .I(N__15440));
    InMux I__3113 (
            .O(N__15466),
            .I(N__15437));
    LocalMux I__3112 (
            .O(N__15463),
            .I(N__15429));
    LocalMux I__3111 (
            .O(N__15460),
            .I(N__15426));
    InMux I__3110 (
            .O(N__15459),
            .I(N__15421));
    InMux I__3109 (
            .O(N__15458),
            .I(N__15421));
    InMux I__3108 (
            .O(N__15457),
            .I(N__15405));
    InMux I__3107 (
            .O(N__15456),
            .I(N__15405));
    InMux I__3106 (
            .O(N__15455),
            .I(N__15405));
    InMux I__3105 (
            .O(N__15454),
            .I(N__15405));
    InMux I__3104 (
            .O(N__15453),
            .I(N__15405));
    InMux I__3103 (
            .O(N__15452),
            .I(N__15405));
    InMux I__3102 (
            .O(N__15451),
            .I(N__15405));
    LocalMux I__3101 (
            .O(N__15440),
            .I(N__15402));
    LocalMux I__3100 (
            .O(N__15437),
            .I(N__15399));
    InMux I__3099 (
            .O(N__15436),
            .I(N__15395));
    InMux I__3098 (
            .O(N__15435),
            .I(N__15392));
    InMux I__3097 (
            .O(N__15434),
            .I(N__15385));
    InMux I__3096 (
            .O(N__15433),
            .I(N__15385));
    InMux I__3095 (
            .O(N__15432),
            .I(N__15385));
    Span4Mux_h I__3094 (
            .O(N__15429),
            .I(N__15382));
    Sp12to4 I__3093 (
            .O(N__15426),
            .I(N__15377));
    LocalMux I__3092 (
            .O(N__15421),
            .I(N__15377));
    InMux I__3091 (
            .O(N__15420),
            .I(N__15374));
    LocalMux I__3090 (
            .O(N__15405),
            .I(N__15367));
    Span4Mux_h I__3089 (
            .O(N__15402),
            .I(N__15367));
    Span4Mux_h I__3088 (
            .O(N__15399),
            .I(N__15367));
    InMux I__3087 (
            .O(N__15398),
            .I(N__15364));
    LocalMux I__3086 (
            .O(N__15395),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__3085 (
            .O(N__15392),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__3084 (
            .O(N__15385),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__3083 (
            .O(N__15382),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv12 I__3082 (
            .O(N__15377),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__3081 (
            .O(N__15374),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__3080 (
            .O(N__15367),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__3079 (
            .O(N__15364),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    CascadeMux I__3078 (
            .O(N__15347),
            .I(N__15338));
    CascadeMux I__3077 (
            .O(N__15346),
            .I(N__15331));
    CascadeMux I__3076 (
            .O(N__15345),
            .I(N__15327));
    CascadeMux I__3075 (
            .O(N__15344),
            .I(N__15324));
    CascadeMux I__3074 (
            .O(N__15343),
            .I(N__15321));
    CascadeMux I__3073 (
            .O(N__15342),
            .I(N__15313));
    CascadeMux I__3072 (
            .O(N__15341),
            .I(N__15310));
    InMux I__3071 (
            .O(N__15338),
            .I(N__15307));
    CascadeMux I__3070 (
            .O(N__15337),
            .I(N__15300));
    CascadeMux I__3069 (
            .O(N__15336),
            .I(N__15297));
    CascadeMux I__3068 (
            .O(N__15335),
            .I(N__15294));
    CascadeMux I__3067 (
            .O(N__15334),
            .I(N__15291));
    InMux I__3066 (
            .O(N__15331),
            .I(N__15286));
    InMux I__3065 (
            .O(N__15330),
            .I(N__15286));
    InMux I__3064 (
            .O(N__15327),
            .I(N__15282));
    InMux I__3063 (
            .O(N__15324),
            .I(N__15275));
    InMux I__3062 (
            .O(N__15321),
            .I(N__15275));
    InMux I__3061 (
            .O(N__15320),
            .I(N__15275));
    InMux I__3060 (
            .O(N__15319),
            .I(N__15262));
    InMux I__3059 (
            .O(N__15318),
            .I(N__15262));
    InMux I__3058 (
            .O(N__15317),
            .I(N__15262));
    InMux I__3057 (
            .O(N__15316),
            .I(N__15262));
    InMux I__3056 (
            .O(N__15313),
            .I(N__15262));
    InMux I__3055 (
            .O(N__15310),
            .I(N__15262));
    LocalMux I__3054 (
            .O(N__15307),
            .I(N__15259));
    InMux I__3053 (
            .O(N__15306),
            .I(N__15242));
    InMux I__3052 (
            .O(N__15305),
            .I(N__15242));
    InMux I__3051 (
            .O(N__15304),
            .I(N__15242));
    InMux I__3050 (
            .O(N__15303),
            .I(N__15242));
    InMux I__3049 (
            .O(N__15300),
            .I(N__15242));
    InMux I__3048 (
            .O(N__15297),
            .I(N__15242));
    InMux I__3047 (
            .O(N__15294),
            .I(N__15242));
    InMux I__3046 (
            .O(N__15291),
            .I(N__15242));
    LocalMux I__3045 (
            .O(N__15286),
            .I(N__15239));
    InMux I__3044 (
            .O(N__15285),
            .I(N__15236));
    LocalMux I__3043 (
            .O(N__15282),
            .I(N__15230));
    LocalMux I__3042 (
            .O(N__15275),
            .I(N__15230));
    LocalMux I__3041 (
            .O(N__15262),
            .I(N__15227));
    Span4Mux_v I__3040 (
            .O(N__15259),
            .I(N__15222));
    LocalMux I__3039 (
            .O(N__15242),
            .I(N__15222));
    Span4Mux_h I__3038 (
            .O(N__15239),
            .I(N__15218));
    LocalMux I__3037 (
            .O(N__15236),
            .I(N__15215));
    InMux I__3036 (
            .O(N__15235),
            .I(N__15212));
    Span4Mux_v I__3035 (
            .O(N__15230),
            .I(N__15209));
    Span4Mux_v I__3034 (
            .O(N__15227),
            .I(N__15204));
    Span4Mux_h I__3033 (
            .O(N__15222),
            .I(N__15204));
    InMux I__3032 (
            .O(N__15221),
            .I(N__15201));
    Span4Mux_v I__3031 (
            .O(N__15218),
            .I(N__15196));
    Span4Mux_h I__3030 (
            .O(N__15215),
            .I(N__15196));
    LocalMux I__3029 (
            .O(N__15212),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    Odrv4 I__3028 (
            .O(N__15209),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    Odrv4 I__3027 (
            .O(N__15204),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    LocalMux I__3026 (
            .O(N__15201),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    Odrv4 I__3025 (
            .O(N__15196),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    InMux I__3024 (
            .O(N__15185),
            .I(N__15181));
    InMux I__3023 (
            .O(N__15184),
            .I(N__15178));
    LocalMux I__3022 (
            .O(N__15181),
            .I(N__15172));
    LocalMux I__3021 (
            .O(N__15178),
            .I(N__15172));
    InMux I__3020 (
            .O(N__15177),
            .I(N__15169));
    Span4Mux_h I__3019 (
            .O(N__15172),
            .I(N__15164));
    LocalMux I__3018 (
            .O(N__15169),
            .I(N__15161));
    InMux I__3017 (
            .O(N__15168),
            .I(N__15156));
    InMux I__3016 (
            .O(N__15167),
            .I(N__15156));
    Odrv4 I__3015 (
            .O(N__15164),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__3014 (
            .O(N__15161),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__3013 (
            .O(N__15156),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__3012 (
            .O(N__15149),
            .I(N__15137));
    InMux I__3011 (
            .O(N__15148),
            .I(N__15124));
    InMux I__3010 (
            .O(N__15147),
            .I(N__15124));
    InMux I__3009 (
            .O(N__15146),
            .I(N__15111));
    InMux I__3008 (
            .O(N__15145),
            .I(N__15111));
    InMux I__3007 (
            .O(N__15144),
            .I(N__15111));
    InMux I__3006 (
            .O(N__15143),
            .I(N__15111));
    InMux I__3005 (
            .O(N__15142),
            .I(N__15111));
    InMux I__3004 (
            .O(N__15141),
            .I(N__15111));
    InMux I__3003 (
            .O(N__15140),
            .I(N__15108));
    InMux I__3002 (
            .O(N__15137),
            .I(N__15100));
    InMux I__3001 (
            .O(N__15136),
            .I(N__15083));
    InMux I__3000 (
            .O(N__15135),
            .I(N__15083));
    InMux I__2999 (
            .O(N__15134),
            .I(N__15083));
    InMux I__2998 (
            .O(N__15133),
            .I(N__15083));
    InMux I__2997 (
            .O(N__15132),
            .I(N__15083));
    InMux I__2996 (
            .O(N__15131),
            .I(N__15083));
    InMux I__2995 (
            .O(N__15130),
            .I(N__15083));
    InMux I__2994 (
            .O(N__15129),
            .I(N__15083));
    LocalMux I__2993 (
            .O(N__15124),
            .I(N__15078));
    LocalMux I__2992 (
            .O(N__15111),
            .I(N__15078));
    LocalMux I__2991 (
            .O(N__15108),
            .I(N__15075));
    InMux I__2990 (
            .O(N__15107),
            .I(N__15071));
    InMux I__2989 (
            .O(N__15106),
            .I(N__15068));
    InMux I__2988 (
            .O(N__15105),
            .I(N__15063));
    InMux I__2987 (
            .O(N__15104),
            .I(N__15063));
    InMux I__2986 (
            .O(N__15103),
            .I(N__15060));
    LocalMux I__2985 (
            .O(N__15100),
            .I(N__15051));
    LocalMux I__2984 (
            .O(N__15083),
            .I(N__15051));
    Span4Mux_h I__2983 (
            .O(N__15078),
            .I(N__15051));
    Span4Mux_h I__2982 (
            .O(N__15075),
            .I(N__15051));
    InMux I__2981 (
            .O(N__15074),
            .I(N__15048));
    LocalMux I__2980 (
            .O(N__15071),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__2979 (
            .O(N__15068),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__2978 (
            .O(N__15063),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__2977 (
            .O(N__15060),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__2976 (
            .O(N__15051),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__2975 (
            .O(N__15048),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    CascadeMux I__2974 (
            .O(N__15035),
            .I(N__15031));
    CascadeMux I__2973 (
            .O(N__15034),
            .I(N__15028));
    InMux I__2972 (
            .O(N__15031),
            .I(N__15025));
    InMux I__2971 (
            .O(N__15028),
            .I(N__15022));
    LocalMux I__2970 (
            .O(N__15025),
            .I(\delay_measurement_inst.elapsed_time_hc_1 ));
    LocalMux I__2969 (
            .O(N__15022),
            .I(\delay_measurement_inst.elapsed_time_hc_1 ));
    CascadeMux I__2968 (
            .O(N__15017),
            .I(N__15014));
    InMux I__2967 (
            .O(N__15014),
            .I(N__15011));
    LocalMux I__2966 (
            .O(N__15011),
            .I(\delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_0_4 ));
    InMux I__2965 (
            .O(N__15008),
            .I(N__15005));
    LocalMux I__2964 (
            .O(N__15005),
            .I(\delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_0_3 ));
    InMux I__2963 (
            .O(N__15002),
            .I(N__14997));
    InMux I__2962 (
            .O(N__15001),
            .I(N__14992));
    InMux I__2961 (
            .O(N__15000),
            .I(N__14992));
    LocalMux I__2960 (
            .O(N__14997),
            .I(\delay_measurement_inst.elapsed_time_hc_2 ));
    LocalMux I__2959 (
            .O(N__14992),
            .I(\delay_measurement_inst.elapsed_time_hc_2 ));
    InMux I__2958 (
            .O(N__14987),
            .I(N__14984));
    LocalMux I__2957 (
            .O(N__14984),
            .I(N__14980));
    InMux I__2956 (
            .O(N__14983),
            .I(N__14977));
    Span4Mux_h I__2955 (
            .O(N__14980),
            .I(N__14974));
    LocalMux I__2954 (
            .O(N__14977),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__2953 (
            .O(N__14974),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__2952 (
            .O(N__14969),
            .I(N__14966));
    LocalMux I__2951 (
            .O(N__14966),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16 ));
    InMux I__2950 (
            .O(N__14963),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ));
    InMux I__2949 (
            .O(N__14960),
            .I(N__14956));
    InMux I__2948 (
            .O(N__14959),
            .I(N__14953));
    LocalMux I__2947 (
            .O(N__14956),
            .I(N__14950));
    LocalMux I__2946 (
            .O(N__14953),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__2945 (
            .O(N__14950),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__2944 (
            .O(N__14945),
            .I(N__14942));
    LocalMux I__2943 (
            .O(N__14942),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17 ));
    InMux I__2942 (
            .O(N__14939),
            .I(bfn_8_19_0_));
    InMux I__2941 (
            .O(N__14936),
            .I(N__14932));
    InMux I__2940 (
            .O(N__14935),
            .I(N__14929));
    LocalMux I__2939 (
            .O(N__14932),
            .I(N__14926));
    LocalMux I__2938 (
            .O(N__14929),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__2937 (
            .O(N__14926),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__2936 (
            .O(N__14921),
            .I(N__14918));
    LocalMux I__2935 (
            .O(N__14918),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18 ));
    InMux I__2934 (
            .O(N__14915),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ));
    InMux I__2933 (
            .O(N__14912),
            .I(N__14908));
    InMux I__2932 (
            .O(N__14911),
            .I(N__14905));
    LocalMux I__2931 (
            .O(N__14908),
            .I(N__14902));
    LocalMux I__2930 (
            .O(N__14905),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__2929 (
            .O(N__14902),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__2928 (
            .O(N__14897),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17 ));
    InMux I__2927 (
            .O(N__14894),
            .I(N__14891));
    LocalMux I__2926 (
            .O(N__14891),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19 ));
    InMux I__2925 (
            .O(N__14888),
            .I(N__14884));
    InMux I__2924 (
            .O(N__14887),
            .I(N__14881));
    LocalMux I__2923 (
            .O(N__14884),
            .I(N__14876));
    LocalMux I__2922 (
            .O(N__14881),
            .I(N__14873));
    InMux I__2921 (
            .O(N__14880),
            .I(N__14868));
    InMux I__2920 (
            .O(N__14879),
            .I(N__14868));
    Span4Mux_h I__2919 (
            .O(N__14876),
            .I(N__14865));
    Span4Mux_h I__2918 (
            .O(N__14873),
            .I(N__14862));
    LocalMux I__2917 (
            .O(N__14868),
            .I(N__14859));
    Odrv4 I__2916 (
            .O(N__14865),
            .I(\phase_controller_inst1.stoper_tr.N_55 ));
    Odrv4 I__2915 (
            .O(N__14862),
            .I(\phase_controller_inst1.stoper_tr.N_55 ));
    Odrv12 I__2914 (
            .O(N__14859),
            .I(\phase_controller_inst1.stoper_tr.N_55 ));
    InMux I__2913 (
            .O(N__14852),
            .I(N__14849));
    LocalMux I__2912 (
            .O(N__14849),
            .I(N__14843));
    InMux I__2911 (
            .O(N__14848),
            .I(N__14836));
    InMux I__2910 (
            .O(N__14847),
            .I(N__14836));
    InMux I__2909 (
            .O(N__14846),
            .I(N__14836));
    Span4Mux_v I__2908 (
            .O(N__14843),
            .I(N__14831));
    LocalMux I__2907 (
            .O(N__14836),
            .I(N__14831));
    Odrv4 I__2906 (
            .O(N__14831),
            .I(\phase_controller_slave.stoper_tr.time_passed11 ));
    InMux I__2905 (
            .O(N__14828),
            .I(N__14816));
    InMux I__2904 (
            .O(N__14827),
            .I(N__14816));
    InMux I__2903 (
            .O(N__14826),
            .I(N__14816));
    InMux I__2902 (
            .O(N__14825),
            .I(N__14807));
    InMux I__2901 (
            .O(N__14824),
            .I(N__14807));
    InMux I__2900 (
            .O(N__14823),
            .I(N__14807));
    LocalMux I__2899 (
            .O(N__14816),
            .I(N__14804));
    CascadeMux I__2898 (
            .O(N__14815),
            .I(N__14801));
    CascadeMux I__2897 (
            .O(N__14814),
            .I(N__14795));
    LocalMux I__2896 (
            .O(N__14807),
            .I(N__14791));
    Span4Mux_v I__2895 (
            .O(N__14804),
            .I(N__14788));
    InMux I__2894 (
            .O(N__14801),
            .I(N__14775));
    InMux I__2893 (
            .O(N__14800),
            .I(N__14775));
    InMux I__2892 (
            .O(N__14799),
            .I(N__14775));
    InMux I__2891 (
            .O(N__14798),
            .I(N__14775));
    InMux I__2890 (
            .O(N__14795),
            .I(N__14775));
    InMux I__2889 (
            .O(N__14794),
            .I(N__14775));
    Span4Mux_v I__2888 (
            .O(N__14791),
            .I(N__14772));
    Span4Mux_h I__2887 (
            .O(N__14788),
            .I(N__14769));
    LocalMux I__2886 (
            .O(N__14775),
            .I(N__14766));
    Odrv4 I__2885 (
            .O(N__14772),
            .I(\phase_controller_inst1.stoper_tr.N_50 ));
    Odrv4 I__2884 (
            .O(N__14769),
            .I(\phase_controller_inst1.stoper_tr.N_50 ));
    Odrv12 I__2883 (
            .O(N__14766),
            .I(\phase_controller_inst1.stoper_tr.N_50 ));
    InMux I__2882 (
            .O(N__14759),
            .I(N__14751));
    InMux I__2881 (
            .O(N__14758),
            .I(N__14751));
    InMux I__2880 (
            .O(N__14757),
            .I(N__14746));
    InMux I__2879 (
            .O(N__14756),
            .I(N__14746));
    LocalMux I__2878 (
            .O(N__14751),
            .I(N__14742));
    LocalMux I__2877 (
            .O(N__14746),
            .I(N__14739));
    InMux I__2876 (
            .O(N__14745),
            .I(N__14736));
    Span4Mux_v I__2875 (
            .O(N__14742),
            .I(N__14729));
    Span4Mux_v I__2874 (
            .O(N__14739),
            .I(N__14729));
    LocalMux I__2873 (
            .O(N__14736),
            .I(N__14729));
    Odrv4 I__2872 (
            .O(N__14729),
            .I(\phase_controller_inst1.stoper_tr.N_32 ));
    CascadeMux I__2871 (
            .O(N__14726),
            .I(\phase_controller_inst1.stoper_tr.N_32_cascade_ ));
    InMux I__2870 (
            .O(N__14723),
            .I(N__14709));
    InMux I__2869 (
            .O(N__14722),
            .I(N__14709));
    InMux I__2868 (
            .O(N__14721),
            .I(N__14709));
    InMux I__2867 (
            .O(N__14720),
            .I(N__14698));
    InMux I__2866 (
            .O(N__14719),
            .I(N__14698));
    InMux I__2865 (
            .O(N__14718),
            .I(N__14698));
    InMux I__2864 (
            .O(N__14717),
            .I(N__14698));
    InMux I__2863 (
            .O(N__14716),
            .I(N__14698));
    LocalMux I__2862 (
            .O(N__14709),
            .I(N__14687));
    LocalMux I__2861 (
            .O(N__14698),
            .I(N__14684));
    InMux I__2860 (
            .O(N__14697),
            .I(N__14667));
    InMux I__2859 (
            .O(N__14696),
            .I(N__14667));
    InMux I__2858 (
            .O(N__14695),
            .I(N__14667));
    InMux I__2857 (
            .O(N__14694),
            .I(N__14667));
    InMux I__2856 (
            .O(N__14693),
            .I(N__14667));
    InMux I__2855 (
            .O(N__14692),
            .I(N__14667));
    InMux I__2854 (
            .O(N__14691),
            .I(N__14667));
    InMux I__2853 (
            .O(N__14690),
            .I(N__14667));
    Span4Mux_h I__2852 (
            .O(N__14687),
            .I(N__14664));
    Span4Mux_h I__2851 (
            .O(N__14684),
            .I(N__14661));
    LocalMux I__2850 (
            .O(N__14667),
            .I(N__14658));
    Odrv4 I__2849 (
            .O(N__14664),
            .I(\phase_controller_inst1.stoper_tr.N_33 ));
    Odrv4 I__2848 (
            .O(N__14661),
            .I(\phase_controller_inst1.stoper_tr.N_33 ));
    Odrv12 I__2847 (
            .O(N__14658),
            .I(\phase_controller_inst1.stoper_tr.N_33 ));
    InMux I__2846 (
            .O(N__14651),
            .I(N__14647));
    InMux I__2845 (
            .O(N__14650),
            .I(N__14644));
    LocalMux I__2844 (
            .O(N__14647),
            .I(N__14641));
    LocalMux I__2843 (
            .O(N__14644),
            .I(N__14636));
    Span4Mux_h I__2842 (
            .O(N__14641),
            .I(N__14636));
    Odrv4 I__2841 (
            .O(N__14636),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ));
    CascadeMux I__2840 (
            .O(N__14633),
            .I(N__14630));
    InMux I__2839 (
            .O(N__14630),
            .I(N__14627));
    LocalMux I__2838 (
            .O(N__14627),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8 ));
    InMux I__2837 (
            .O(N__14624),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ));
    InMux I__2836 (
            .O(N__14621),
            .I(N__14617));
    InMux I__2835 (
            .O(N__14620),
            .I(N__14614));
    LocalMux I__2834 (
            .O(N__14617),
            .I(N__14611));
    LocalMux I__2833 (
            .O(N__14614),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__2832 (
            .O(N__14611),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__2831 (
            .O(N__14606),
            .I(N__14603));
    LocalMux I__2830 (
            .O(N__14603),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9 ));
    InMux I__2829 (
            .O(N__14600),
            .I(bfn_8_18_0_));
    InMux I__2828 (
            .O(N__14597),
            .I(N__14593));
    InMux I__2827 (
            .O(N__14596),
            .I(N__14590));
    LocalMux I__2826 (
            .O(N__14593),
            .I(N__14587));
    LocalMux I__2825 (
            .O(N__14590),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv4 I__2824 (
            .O(N__14587),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ));
    CascadeMux I__2823 (
            .O(N__14582),
            .I(N__14579));
    InMux I__2822 (
            .O(N__14579),
            .I(N__14576));
    LocalMux I__2821 (
            .O(N__14576),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10 ));
    InMux I__2820 (
            .O(N__14573),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ));
    InMux I__2819 (
            .O(N__14570),
            .I(N__14566));
    InMux I__2818 (
            .O(N__14569),
            .I(N__14563));
    LocalMux I__2817 (
            .O(N__14566),
            .I(N__14560));
    LocalMux I__2816 (
            .O(N__14563),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv4 I__2815 (
            .O(N__14560),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__2814 (
            .O(N__14555),
            .I(N__14552));
    LocalMux I__2813 (
            .O(N__14552),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11 ));
    InMux I__2812 (
            .O(N__14549),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ));
    InMux I__2811 (
            .O(N__14546),
            .I(N__14543));
    LocalMux I__2810 (
            .O(N__14543),
            .I(N__14539));
    InMux I__2809 (
            .O(N__14542),
            .I(N__14536));
    Span4Mux_h I__2808 (
            .O(N__14539),
            .I(N__14533));
    LocalMux I__2807 (
            .O(N__14536),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__2806 (
            .O(N__14533),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ));
    CascadeMux I__2805 (
            .O(N__14528),
            .I(N__14525));
    InMux I__2804 (
            .O(N__14525),
            .I(N__14522));
    LocalMux I__2803 (
            .O(N__14522),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12 ));
    InMux I__2802 (
            .O(N__14519),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ));
    InMux I__2801 (
            .O(N__14516),
            .I(N__14512));
    InMux I__2800 (
            .O(N__14515),
            .I(N__14509));
    LocalMux I__2799 (
            .O(N__14512),
            .I(N__14506));
    LocalMux I__2798 (
            .O(N__14509),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__2797 (
            .O(N__14506),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__2796 (
            .O(N__14501),
            .I(N__14498));
    LocalMux I__2795 (
            .O(N__14498),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13 ));
    InMux I__2794 (
            .O(N__14495),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ));
    InMux I__2793 (
            .O(N__14492),
            .I(N__14488));
    InMux I__2792 (
            .O(N__14491),
            .I(N__14485));
    LocalMux I__2791 (
            .O(N__14488),
            .I(N__14482));
    LocalMux I__2790 (
            .O(N__14485),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__2789 (
            .O(N__14482),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ));
    CascadeMux I__2788 (
            .O(N__14477),
            .I(N__14474));
    InMux I__2787 (
            .O(N__14474),
            .I(N__14471));
    LocalMux I__2786 (
            .O(N__14471),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14 ));
    InMux I__2785 (
            .O(N__14468),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ));
    InMux I__2784 (
            .O(N__14465),
            .I(N__14461));
    InMux I__2783 (
            .O(N__14464),
            .I(N__14458));
    LocalMux I__2782 (
            .O(N__14461),
            .I(N__14455));
    LocalMux I__2781 (
            .O(N__14458),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv4 I__2780 (
            .O(N__14455),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__2779 (
            .O(N__14450),
            .I(N__14447));
    LocalMux I__2778 (
            .O(N__14447),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15 ));
    InMux I__2777 (
            .O(N__14444),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ));
    InMux I__2776 (
            .O(N__14441),
            .I(N__14437));
    InMux I__2775 (
            .O(N__14440),
            .I(N__14434));
    LocalMux I__2774 (
            .O(N__14437),
            .I(N__14430));
    LocalMux I__2773 (
            .O(N__14434),
            .I(N__14427));
    InMux I__2772 (
            .O(N__14433),
            .I(N__14424));
    Odrv4 I__2771 (
            .O(N__14430),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv12 I__2770 (
            .O(N__14427),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__2769 (
            .O(N__14424),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ));
    CascadeMux I__2768 (
            .O(N__14417),
            .I(N__14414));
    InMux I__2767 (
            .O(N__14414),
            .I(N__14411));
    LocalMux I__2766 (
            .O(N__14411),
            .I(N__14408));
    Span4Mux_h I__2765 (
            .O(N__14408),
            .I(N__14405));
    Odrv4 I__2764 (
            .O(N__14405),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ));
    InMux I__2763 (
            .O(N__14402),
            .I(N__14399));
    LocalMux I__2762 (
            .O(N__14399),
            .I(N__14395));
    InMux I__2761 (
            .O(N__14398),
            .I(N__14392));
    Odrv12 I__2760 (
            .O(N__14395),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__2759 (
            .O(N__14392),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__2758 (
            .O(N__14387),
            .I(N__14384));
    LocalMux I__2757 (
            .O(N__14384),
            .I(N__14381));
    Span4Mux_h I__2756 (
            .O(N__14381),
            .I(N__14378));
    Odrv4 I__2755 (
            .O(N__14378),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2 ));
    InMux I__2754 (
            .O(N__14375),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ));
    InMux I__2753 (
            .O(N__14372),
            .I(N__14369));
    LocalMux I__2752 (
            .O(N__14369),
            .I(N__14365));
    InMux I__2751 (
            .O(N__14368),
            .I(N__14362));
    Odrv12 I__2750 (
            .O(N__14365),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__2749 (
            .O(N__14362),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ));
    CascadeMux I__2748 (
            .O(N__14357),
            .I(N__14354));
    InMux I__2747 (
            .O(N__14354),
            .I(N__14351));
    LocalMux I__2746 (
            .O(N__14351),
            .I(N__14348));
    Span4Mux_h I__2745 (
            .O(N__14348),
            .I(N__14345));
    Odrv4 I__2744 (
            .O(N__14345),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6 ));
    CascadeMux I__2743 (
            .O(N__14342),
            .I(N__14339));
    InMux I__2742 (
            .O(N__14339),
            .I(N__14336));
    LocalMux I__2741 (
            .O(N__14336),
            .I(N__14333));
    Odrv12 I__2740 (
            .O(N__14333),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3 ));
    InMux I__2739 (
            .O(N__14330),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ));
    CascadeMux I__2738 (
            .O(N__14327),
            .I(N__14324));
    InMux I__2737 (
            .O(N__14324),
            .I(N__14321));
    LocalMux I__2736 (
            .O(N__14321),
            .I(N__14317));
    InMux I__2735 (
            .O(N__14320),
            .I(N__14314));
    Odrv12 I__2734 (
            .O(N__14317),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__2733 (
            .O(N__14314),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__2732 (
            .O(N__14309),
            .I(N__14306));
    LocalMux I__2731 (
            .O(N__14306),
            .I(N__14303));
    Span4Mux_h I__2730 (
            .O(N__14303),
            .I(N__14300));
    Odrv4 I__2729 (
            .O(N__14300),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4 ));
    InMux I__2728 (
            .O(N__14297),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ));
    CascadeMux I__2727 (
            .O(N__14294),
            .I(N__14291));
    InMux I__2726 (
            .O(N__14291),
            .I(N__14288));
    LocalMux I__2725 (
            .O(N__14288),
            .I(N__14284));
    InMux I__2724 (
            .O(N__14287),
            .I(N__14281));
    Odrv12 I__2723 (
            .O(N__14284),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__2722 (
            .O(N__14281),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ));
    CascadeMux I__2721 (
            .O(N__14276),
            .I(N__14273));
    InMux I__2720 (
            .O(N__14273),
            .I(N__14270));
    LocalMux I__2719 (
            .O(N__14270),
            .I(N__14267));
    Span4Mux_h I__2718 (
            .O(N__14267),
            .I(N__14264));
    Odrv4 I__2717 (
            .O(N__14264),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5 ));
    InMux I__2716 (
            .O(N__14261),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ));
    InMux I__2715 (
            .O(N__14258),
            .I(N__14255));
    LocalMux I__2714 (
            .O(N__14255),
            .I(N__14251));
    InMux I__2713 (
            .O(N__14254),
            .I(N__14248));
    Odrv12 I__2712 (
            .O(N__14251),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__2711 (
            .O(N__14248),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ));
    CascadeMux I__2710 (
            .O(N__14243),
            .I(N__14240));
    InMux I__2709 (
            .O(N__14240),
            .I(N__14237));
    LocalMux I__2708 (
            .O(N__14237),
            .I(N__14234));
    Span4Mux_h I__2707 (
            .O(N__14234),
            .I(N__14231));
    Odrv4 I__2706 (
            .O(N__14231),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6 ));
    InMux I__2705 (
            .O(N__14228),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ));
    InMux I__2704 (
            .O(N__14225),
            .I(N__14221));
    InMux I__2703 (
            .O(N__14224),
            .I(N__14218));
    LocalMux I__2702 (
            .O(N__14221),
            .I(N__14215));
    LocalMux I__2701 (
            .O(N__14218),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv4 I__2700 (
            .O(N__14215),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__2699 (
            .O(N__14210),
            .I(N__14207));
    LocalMux I__2698 (
            .O(N__14207),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7 ));
    InMux I__2697 (
            .O(N__14204),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ));
    InMux I__2696 (
            .O(N__14201),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    InMux I__2695 (
            .O(N__14198),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    InMux I__2694 (
            .O(N__14195),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    InMux I__2693 (
            .O(N__14192),
            .I(bfn_8_16_0_));
    InMux I__2692 (
            .O(N__14189),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    InMux I__2691 (
            .O(N__14186),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    InMux I__2690 (
            .O(N__14183),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__2689 (
            .O(N__14180),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__2688 (
            .O(N__14177),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    CEMux I__2687 (
            .O(N__14174),
            .I(N__14162));
    CEMux I__2686 (
            .O(N__14173),
            .I(N__14162));
    CEMux I__2685 (
            .O(N__14172),
            .I(N__14162));
    CEMux I__2684 (
            .O(N__14171),
            .I(N__14162));
    GlobalMux I__2683 (
            .O(N__14162),
            .I(N__14159));
    gio2CtrlBuf I__2682 (
            .O(N__14159),
            .I(\delay_measurement_inst.delay_tr_timer.N_256_i_g ));
    InMux I__2681 (
            .O(N__14156),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    InMux I__2680 (
            .O(N__14153),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    InMux I__2679 (
            .O(N__14150),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    InMux I__2678 (
            .O(N__14147),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    InMux I__2677 (
            .O(N__14144),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    InMux I__2676 (
            .O(N__14141),
            .I(bfn_8_15_0_));
    InMux I__2675 (
            .O(N__14138),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    InMux I__2674 (
            .O(N__14135),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    InMux I__2673 (
            .O(N__14132),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    InMux I__2672 (
            .O(N__14129),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    InMux I__2671 (
            .O(N__14126),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    InMux I__2670 (
            .O(N__14123),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    InMux I__2669 (
            .O(N__14120),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    InMux I__2668 (
            .O(N__14117),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    InMux I__2667 (
            .O(N__14114),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    InMux I__2666 (
            .O(N__14111),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    InMux I__2665 (
            .O(N__14108),
            .I(bfn_8_14_0_));
    InMux I__2664 (
            .O(N__14105),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    InMux I__2663 (
            .O(N__14102),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    InMux I__2662 (
            .O(N__14099),
            .I(N__14096));
    LocalMux I__2661 (
            .O(N__14096),
            .I(N__14092));
    InMux I__2660 (
            .O(N__14095),
            .I(N__14089));
    Span4Mux_h I__2659 (
            .O(N__14092),
            .I(N__14085));
    LocalMux I__2658 (
            .O(N__14089),
            .I(N__14082));
    InMux I__2657 (
            .O(N__14088),
            .I(N__14079));
    Span4Mux_v I__2656 (
            .O(N__14085),
            .I(N__14076));
    Span4Mux_v I__2655 (
            .O(N__14082),
            .I(N__14071));
    LocalMux I__2654 (
            .O(N__14079),
            .I(N__14071));
    Odrv4 I__2653 (
            .O(N__14076),
            .I(measured_delay_hc_6));
    Odrv4 I__2652 (
            .O(N__14071),
            .I(measured_delay_hc_6));
    InMux I__2651 (
            .O(N__14066),
            .I(N__14063));
    LocalMux I__2650 (
            .O(N__14063),
            .I(N__14058));
    InMux I__2649 (
            .O(N__14062),
            .I(N__14055));
    InMux I__2648 (
            .O(N__14061),
            .I(N__14051));
    Span4Mux_v I__2647 (
            .O(N__14058),
            .I(N__14048));
    LocalMux I__2646 (
            .O(N__14055),
            .I(N__14045));
    InMux I__2645 (
            .O(N__14054),
            .I(N__14042));
    LocalMux I__2644 (
            .O(N__14051),
            .I(N__14039));
    Span4Mux_v I__2643 (
            .O(N__14048),
            .I(N__14032));
    Span4Mux_v I__2642 (
            .O(N__14045),
            .I(N__14032));
    LocalMux I__2641 (
            .O(N__14042),
            .I(N__14032));
    Span4Mux_h I__2640 (
            .O(N__14039),
            .I(N__14029));
    Odrv4 I__2639 (
            .O(N__14032),
            .I(measured_delay_hc_17));
    Odrv4 I__2638 (
            .O(N__14029),
            .I(measured_delay_hc_17));
    InMux I__2637 (
            .O(N__14024),
            .I(N__14021));
    LocalMux I__2636 (
            .O(N__14021),
            .I(N__14016));
    InMux I__2635 (
            .O(N__14020),
            .I(N__14012));
    InMux I__2634 (
            .O(N__14019),
            .I(N__14009));
    Span4Mux_h I__2633 (
            .O(N__14016),
            .I(N__14006));
    InMux I__2632 (
            .O(N__14015),
            .I(N__14003));
    LocalMux I__2631 (
            .O(N__14012),
            .I(N__14000));
    LocalMux I__2630 (
            .O(N__14009),
            .I(N__13997));
    Span4Mux_v I__2629 (
            .O(N__14006),
            .I(N__13994));
    LocalMux I__2628 (
            .O(N__14003),
            .I(N__13991));
    Span4Mux_h I__2627 (
            .O(N__14000),
            .I(N__13986));
    Span4Mux_h I__2626 (
            .O(N__13997),
            .I(N__13986));
    Odrv4 I__2625 (
            .O(N__13994),
            .I(measured_delay_hc_16));
    Odrv4 I__2624 (
            .O(N__13991),
            .I(measured_delay_hc_16));
    Odrv4 I__2623 (
            .O(N__13986),
            .I(measured_delay_hc_16));
    InMux I__2622 (
            .O(N__13979),
            .I(N__13976));
    LocalMux I__2621 (
            .O(N__13976),
            .I(N__13970));
    InMux I__2620 (
            .O(N__13975),
            .I(N__13967));
    InMux I__2619 (
            .O(N__13974),
            .I(N__13961));
    InMux I__2618 (
            .O(N__13973),
            .I(N__13961));
    Span4Mux_v I__2617 (
            .O(N__13970),
            .I(N__13958));
    LocalMux I__2616 (
            .O(N__13967),
            .I(N__13955));
    InMux I__2615 (
            .O(N__13966),
            .I(N__13952));
    LocalMux I__2614 (
            .O(N__13961),
            .I(N__13949));
    Span4Mux_v I__2613 (
            .O(N__13958),
            .I(N__13942));
    Span4Mux_v I__2612 (
            .O(N__13955),
            .I(N__13942));
    LocalMux I__2611 (
            .O(N__13952),
            .I(N__13942));
    Span4Mux_h I__2610 (
            .O(N__13949),
            .I(N__13939));
    Odrv4 I__2609 (
            .O(N__13942),
            .I(measured_delay_hc_14));
    Odrv4 I__2608 (
            .O(N__13939),
            .I(measured_delay_hc_14));
    InMux I__2607 (
            .O(N__13934),
            .I(N__13930));
    InMux I__2606 (
            .O(N__13933),
            .I(N__13927));
    LocalMux I__2605 (
            .O(N__13930),
            .I(N__13923));
    LocalMux I__2604 (
            .O(N__13927),
            .I(N__13919));
    InMux I__2603 (
            .O(N__13926),
            .I(N__13916));
    Span4Mux_h I__2602 (
            .O(N__13923),
            .I(N__13913));
    InMux I__2601 (
            .O(N__13922),
            .I(N__13910));
    Span4Mux_h I__2600 (
            .O(N__13919),
            .I(N__13907));
    LocalMux I__2599 (
            .O(N__13916),
            .I(N__13904));
    Span4Mux_v I__2598 (
            .O(N__13913),
            .I(N__13901));
    LocalMux I__2597 (
            .O(N__13910),
            .I(N__13898));
    Span4Mux_v I__2596 (
            .O(N__13907),
            .I(N__13893));
    Span4Mux_h I__2595 (
            .O(N__13904),
            .I(N__13893));
    Span4Mux_v I__2594 (
            .O(N__13901),
            .I(N__13888));
    Span4Mux_h I__2593 (
            .O(N__13898),
            .I(N__13888));
    Odrv4 I__2592 (
            .O(N__13893),
            .I(measured_delay_hc_18));
    Odrv4 I__2591 (
            .O(N__13888),
            .I(measured_delay_hc_18));
    InMux I__2590 (
            .O(N__13883),
            .I(N__13878));
    InMux I__2589 (
            .O(N__13882),
            .I(N__13875));
    InMux I__2588 (
            .O(N__13881),
            .I(N__13872));
    LocalMux I__2587 (
            .O(N__13878),
            .I(N__13868));
    LocalMux I__2586 (
            .O(N__13875),
            .I(N__13863));
    LocalMux I__2585 (
            .O(N__13872),
            .I(N__13863));
    InMux I__2584 (
            .O(N__13871),
            .I(N__13860));
    Span12Mux_v I__2583 (
            .O(N__13868),
            .I(N__13857));
    Span4Mux_v I__2582 (
            .O(N__13863),
            .I(N__13854));
    LocalMux I__2581 (
            .O(N__13860),
            .I(measured_delay_hc_7));
    Odrv12 I__2580 (
            .O(N__13857),
            .I(measured_delay_hc_7));
    Odrv4 I__2579 (
            .O(N__13854),
            .I(measured_delay_hc_7));
    InMux I__2578 (
            .O(N__13847),
            .I(N__13843));
    InMux I__2577 (
            .O(N__13846),
            .I(N__13839));
    LocalMux I__2576 (
            .O(N__13843),
            .I(N__13835));
    InMux I__2575 (
            .O(N__13842),
            .I(N__13832));
    LocalMux I__2574 (
            .O(N__13839),
            .I(N__13829));
    InMux I__2573 (
            .O(N__13838),
            .I(N__13826));
    Span12Mux_s7_h I__2572 (
            .O(N__13835),
            .I(N__13823));
    LocalMux I__2571 (
            .O(N__13832),
            .I(N__13820));
    Span4Mux_h I__2570 (
            .O(N__13829),
            .I(N__13817));
    LocalMux I__2569 (
            .O(N__13826),
            .I(measured_delay_hc_8));
    Odrv12 I__2568 (
            .O(N__13823),
            .I(measured_delay_hc_8));
    Odrv4 I__2567 (
            .O(N__13820),
            .I(measured_delay_hc_8));
    Odrv4 I__2566 (
            .O(N__13817),
            .I(measured_delay_hc_8));
    InMux I__2565 (
            .O(N__13808),
            .I(bfn_8_13_0_));
    InMux I__2564 (
            .O(N__13805),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    InMux I__2563 (
            .O(N__13802),
            .I(N__13799));
    LocalMux I__2562 (
            .O(N__13799),
            .I(N__13795));
    InMux I__2561 (
            .O(N__13798),
            .I(N__13792));
    Span4Mux_v I__2560 (
            .O(N__13795),
            .I(N__13788));
    LocalMux I__2559 (
            .O(N__13792),
            .I(N__13785));
    InMux I__2558 (
            .O(N__13791),
            .I(N__13782));
    Span4Mux_v I__2557 (
            .O(N__13788),
            .I(N__13775));
    Span4Mux_v I__2556 (
            .O(N__13785),
            .I(N__13775));
    LocalMux I__2555 (
            .O(N__13782),
            .I(N__13775));
    Odrv4 I__2554 (
            .O(N__13775),
            .I(measured_delay_hc_11));
    InMux I__2553 (
            .O(N__13772),
            .I(N__13769));
    LocalMux I__2552 (
            .O(N__13769),
            .I(N__13765));
    InMux I__2551 (
            .O(N__13768),
            .I(N__13762));
    Span4Mux_v I__2550 (
            .O(N__13765),
            .I(N__13758));
    LocalMux I__2549 (
            .O(N__13762),
            .I(N__13755));
    InMux I__2548 (
            .O(N__13761),
            .I(N__13752));
    Span4Mux_v I__2547 (
            .O(N__13758),
            .I(N__13745));
    Span4Mux_v I__2546 (
            .O(N__13755),
            .I(N__13745));
    LocalMux I__2545 (
            .O(N__13752),
            .I(N__13745));
    Odrv4 I__2544 (
            .O(N__13745),
            .I(measured_delay_hc_12));
    CascadeMux I__2543 (
            .O(N__13742),
            .I(N__13738));
    CascadeMux I__2542 (
            .O(N__13741),
            .I(N__13735));
    InMux I__2541 (
            .O(N__13738),
            .I(N__13732));
    InMux I__2540 (
            .O(N__13735),
            .I(N__13729));
    LocalMux I__2539 (
            .O(N__13732),
            .I(N__13726));
    LocalMux I__2538 (
            .O(N__13729),
            .I(N__13722));
    Span4Mux_v I__2537 (
            .O(N__13726),
            .I(N__13719));
    InMux I__2536 (
            .O(N__13725),
            .I(N__13716));
    Span4Mux_h I__2535 (
            .O(N__13722),
            .I(N__13713));
    Span4Mux_v I__2534 (
            .O(N__13719),
            .I(N__13708));
    LocalMux I__2533 (
            .O(N__13716),
            .I(N__13708));
    Odrv4 I__2532 (
            .O(N__13713),
            .I(measured_delay_hc_3));
    Odrv4 I__2531 (
            .O(N__13708),
            .I(measured_delay_hc_3));
    InMux I__2530 (
            .O(N__13703),
            .I(N__13700));
    LocalMux I__2529 (
            .O(N__13700),
            .I(N__13696));
    InMux I__2528 (
            .O(N__13699),
            .I(N__13693));
    Span4Mux_v I__2527 (
            .O(N__13696),
            .I(N__13689));
    LocalMux I__2526 (
            .O(N__13693),
            .I(N__13686));
    InMux I__2525 (
            .O(N__13692),
            .I(N__13683));
    Span4Mux_v I__2524 (
            .O(N__13689),
            .I(N__13676));
    Span4Mux_v I__2523 (
            .O(N__13686),
            .I(N__13676));
    LocalMux I__2522 (
            .O(N__13683),
            .I(N__13676));
    Odrv4 I__2521 (
            .O(N__13676),
            .I(measured_delay_hc_4));
    CascadeMux I__2520 (
            .O(N__13673),
            .I(N__13666));
    InMux I__2519 (
            .O(N__13672),
            .I(N__13655));
    InMux I__2518 (
            .O(N__13671),
            .I(N__13655));
    InMux I__2517 (
            .O(N__13670),
            .I(N__13655));
    InMux I__2516 (
            .O(N__13669),
            .I(N__13655));
    InMux I__2515 (
            .O(N__13666),
            .I(N__13655));
    LocalMux I__2514 (
            .O(N__13655),
            .I(\delay_measurement_inst.delay_hc_reg_3_0_a2_0_6 ));
    CascadeMux I__2513 (
            .O(N__13652),
            .I(N__13649));
    InMux I__2512 (
            .O(N__13649),
            .I(N__13645));
    CascadeMux I__2511 (
            .O(N__13648),
            .I(N__13642));
    LocalMux I__2510 (
            .O(N__13645),
            .I(N__13639));
    InMux I__2509 (
            .O(N__13642),
            .I(N__13636));
    Span4Mux_h I__2508 (
            .O(N__13639),
            .I(N__13633));
    LocalMux I__2507 (
            .O(N__13636),
            .I(N__13630));
    Span4Mux_v I__2506 (
            .O(N__13633),
            .I(N__13627));
    Span4Mux_h I__2505 (
            .O(N__13630),
            .I(N__13624));
    Odrv4 I__2504 (
            .O(N__13627),
            .I(measured_delay_hc_1));
    Odrv4 I__2503 (
            .O(N__13624),
            .I(measured_delay_hc_1));
    InMux I__2502 (
            .O(N__13619),
            .I(N__13615));
    InMux I__2501 (
            .O(N__13618),
            .I(N__13612));
    LocalMux I__2500 (
            .O(N__13615),
            .I(N__13608));
    LocalMux I__2499 (
            .O(N__13612),
            .I(N__13605));
    InMux I__2498 (
            .O(N__13611),
            .I(N__13602));
    Span12Mux_v I__2497 (
            .O(N__13608),
            .I(N__13599));
    Span4Mux_v I__2496 (
            .O(N__13605),
            .I(N__13594));
    LocalMux I__2495 (
            .O(N__13602),
            .I(N__13594));
    Odrv12 I__2494 (
            .O(N__13599),
            .I(measured_delay_hc_10));
    Odrv4 I__2493 (
            .O(N__13594),
            .I(measured_delay_hc_10));
    InMux I__2492 (
            .O(N__13589),
            .I(N__13586));
    LocalMux I__2491 (
            .O(N__13586),
            .I(N__13581));
    InMux I__2490 (
            .O(N__13585),
            .I(N__13578));
    InMux I__2489 (
            .O(N__13584),
            .I(N__13575));
    Span4Mux_v I__2488 (
            .O(N__13581),
            .I(N__13572));
    LocalMux I__2487 (
            .O(N__13578),
            .I(N__13569));
    LocalMux I__2486 (
            .O(N__13575),
            .I(N__13566));
    Span4Mux_v I__2485 (
            .O(N__13572),
            .I(N__13559));
    Span4Mux_v I__2484 (
            .O(N__13569),
            .I(N__13559));
    Span4Mux_v I__2483 (
            .O(N__13566),
            .I(N__13559));
    Odrv4 I__2482 (
            .O(N__13559),
            .I(measured_delay_hc_9));
    InMux I__2481 (
            .O(N__13556),
            .I(N__13543));
    InMux I__2480 (
            .O(N__13555),
            .I(N__13543));
    InMux I__2479 (
            .O(N__13554),
            .I(N__13543));
    CascadeMux I__2478 (
            .O(N__13553),
            .I(N__13537));
    InMux I__2477 (
            .O(N__13552),
            .I(N__13530));
    InMux I__2476 (
            .O(N__13551),
            .I(N__13530));
    InMux I__2475 (
            .O(N__13550),
            .I(N__13530));
    LocalMux I__2474 (
            .O(N__13543),
            .I(N__13527));
    InMux I__2473 (
            .O(N__13542),
            .I(N__13522));
    InMux I__2472 (
            .O(N__13541),
            .I(N__13522));
    InMux I__2471 (
            .O(N__13540),
            .I(N__13517));
    InMux I__2470 (
            .O(N__13537),
            .I(N__13517));
    LocalMux I__2469 (
            .O(N__13530),
            .I(N__13514));
    Span4Mux_v I__2468 (
            .O(N__13527),
            .I(N__13507));
    LocalMux I__2467 (
            .O(N__13522),
            .I(N__13507));
    LocalMux I__2466 (
            .O(N__13517),
            .I(N__13507));
    Span4Mux_v I__2465 (
            .O(N__13514),
            .I(N__13502));
    Span4Mux_v I__2464 (
            .O(N__13507),
            .I(N__13502));
    Odrv4 I__2463 (
            .O(N__13502),
            .I(measured_delay_hc_15));
    CascadeMux I__2462 (
            .O(N__13499),
            .I(N__13495));
    InMux I__2461 (
            .O(N__13498),
            .I(N__13492));
    InMux I__2460 (
            .O(N__13495),
            .I(N__13487));
    LocalMux I__2459 (
            .O(N__13492),
            .I(N__13484));
    InMux I__2458 (
            .O(N__13491),
            .I(N__13481));
    CascadeMux I__2457 (
            .O(N__13490),
            .I(N__13478));
    LocalMux I__2456 (
            .O(N__13487),
            .I(N__13475));
    Span4Mux_v I__2455 (
            .O(N__13484),
            .I(N__13472));
    LocalMux I__2454 (
            .O(N__13481),
            .I(N__13469));
    InMux I__2453 (
            .O(N__13478),
            .I(N__13466));
    Span4Mux_h I__2452 (
            .O(N__13475),
            .I(N__13463));
    Span4Mux_v I__2451 (
            .O(N__13472),
            .I(N__13458));
    Span4Mux_v I__2450 (
            .O(N__13469),
            .I(N__13458));
    LocalMux I__2449 (
            .O(N__13466),
            .I(N__13455));
    Span4Mux_h I__2448 (
            .O(N__13463),
            .I(N__13452));
    Odrv4 I__2447 (
            .O(N__13458),
            .I(measured_delay_hc_19));
    Odrv12 I__2446 (
            .O(N__13455),
            .I(measured_delay_hc_19));
    Odrv4 I__2445 (
            .O(N__13452),
            .I(measured_delay_hc_19));
    CascadeMux I__2444 (
            .O(N__13445),
            .I(N__13442));
    InMux I__2443 (
            .O(N__13442),
            .I(N__13439));
    LocalMux I__2442 (
            .O(N__13439),
            .I(N__13436));
    Span4Mux_h I__2441 (
            .O(N__13436),
            .I(N__13433));
    Odrv4 I__2440 (
            .O(N__13433),
            .I(\phase_controller_slave.stoper_tr.time_passed_1_sqmuxa ));
    InMux I__2439 (
            .O(N__13430),
            .I(N__13427));
    LocalMux I__2438 (
            .O(N__13427),
            .I(N__13424));
    Odrv12 I__2437 (
            .O(N__13424),
            .I(il_min_comp2_D1));
    CascadeMux I__2436 (
            .O(N__13421),
            .I(N__13418));
    InMux I__2435 (
            .O(N__13418),
            .I(N__13413));
    InMux I__2434 (
            .O(N__13417),
            .I(N__13410));
    InMux I__2433 (
            .O(N__13416),
            .I(N__13407));
    LocalMux I__2432 (
            .O(N__13413),
            .I(N__13404));
    LocalMux I__2431 (
            .O(N__13410),
            .I(N__13401));
    LocalMux I__2430 (
            .O(N__13407),
            .I(N__13398));
    Span4Mux_v I__2429 (
            .O(N__13404),
            .I(N__13395));
    Span4Mux_h I__2428 (
            .O(N__13401),
            .I(N__13392));
    Span4Mux_h I__2427 (
            .O(N__13398),
            .I(N__13389));
    Odrv4 I__2426 (
            .O(N__13395),
            .I(il_min_comp2_D2));
    Odrv4 I__2425 (
            .O(N__13392),
            .I(il_min_comp2_D2));
    Odrv4 I__2424 (
            .O(N__13389),
            .I(il_min_comp2_D2));
    InMux I__2423 (
            .O(N__13382),
            .I(N__13379));
    LocalMux I__2422 (
            .O(N__13379),
            .I(N__13374));
    InMux I__2421 (
            .O(N__13378),
            .I(N__13371));
    InMux I__2420 (
            .O(N__13377),
            .I(N__13368));
    Span4Mux_h I__2419 (
            .O(N__13374),
            .I(N__13365));
    LocalMux I__2418 (
            .O(N__13371),
            .I(N__13362));
    LocalMux I__2417 (
            .O(N__13368),
            .I(N__13359));
    Span4Mux_v I__2416 (
            .O(N__13365),
            .I(N__13356));
    Span4Mux_h I__2415 (
            .O(N__13362),
            .I(N__13353));
    Span4Mux_h I__2414 (
            .O(N__13359),
            .I(N__13350));
    Odrv4 I__2413 (
            .O(N__13356),
            .I(measured_delay_hc_5));
    Odrv4 I__2412 (
            .O(N__13353),
            .I(measured_delay_hc_5));
    Odrv4 I__2411 (
            .O(N__13350),
            .I(measured_delay_hc_5));
    InMux I__2410 (
            .O(N__13343),
            .I(N__13340));
    LocalMux I__2409 (
            .O(N__13340),
            .I(N__13336));
    InMux I__2408 (
            .O(N__13339),
            .I(N__13333));
    Span4Mux_h I__2407 (
            .O(N__13336),
            .I(N__13329));
    LocalMux I__2406 (
            .O(N__13333),
            .I(N__13326));
    InMux I__2405 (
            .O(N__13332),
            .I(N__13323));
    Span4Mux_v I__2404 (
            .O(N__13329),
            .I(N__13320));
    Span4Mux_h I__2403 (
            .O(N__13326),
            .I(N__13317));
    LocalMux I__2402 (
            .O(N__13323),
            .I(N__13314));
    Odrv4 I__2401 (
            .O(N__13320),
            .I(measured_delay_hc_2));
    Odrv4 I__2400 (
            .O(N__13317),
            .I(measured_delay_hc_2));
    Odrv12 I__2399 (
            .O(N__13314),
            .I(measured_delay_hc_2));
    CascadeMux I__2398 (
            .O(N__13307),
            .I(N__13303));
    InMux I__2397 (
            .O(N__13306),
            .I(N__13297));
    InMux I__2396 (
            .O(N__13303),
            .I(N__13297));
    InMux I__2395 (
            .O(N__13302),
            .I(N__13294));
    LocalMux I__2394 (
            .O(N__13297),
            .I(\phase_controller_slave.stateZ0Z_2 ));
    LocalMux I__2393 (
            .O(N__13294),
            .I(\phase_controller_slave.stateZ0Z_2 ));
    InMux I__2392 (
            .O(N__13289),
            .I(N__13283));
    InMux I__2391 (
            .O(N__13288),
            .I(N__13283));
    LocalMux I__2390 (
            .O(N__13283),
            .I(N__13278));
    InMux I__2389 (
            .O(N__13282),
            .I(N__13275));
    InMux I__2388 (
            .O(N__13281),
            .I(N__13272));
    Span4Mux_h I__2387 (
            .O(N__13278),
            .I(N__13267));
    LocalMux I__2386 (
            .O(N__13275),
            .I(N__13267));
    LocalMux I__2385 (
            .O(N__13272),
            .I(\phase_controller_slave.hc_time_passed ));
    Odrv4 I__2384 (
            .O(N__13267),
            .I(\phase_controller_slave.hc_time_passed ));
    CascadeMux I__2383 (
            .O(N__13262),
            .I(N__13259));
    InMux I__2382 (
            .O(N__13259),
            .I(N__13256));
    LocalMux I__2381 (
            .O(N__13256),
            .I(N__13253));
    Odrv4 I__2380 (
            .O(N__13253),
            .I(\phase_controller_slave.start_timer_hc_RNOZ0Z_0 ));
    InMux I__2379 (
            .O(N__13250),
            .I(N__13247));
    LocalMux I__2378 (
            .O(N__13247),
            .I(N__13244));
    Span4Mux_v I__2377 (
            .O(N__13244),
            .I(N__13241));
    Span4Mux_v I__2376 (
            .O(N__13241),
            .I(N__13238));
    Odrv4 I__2375 (
            .O(N__13238),
            .I(il_max_comp1_c));
    InMux I__2374 (
            .O(N__13235),
            .I(N__13232));
    LocalMux I__2373 (
            .O(N__13232),
            .I(N__13229));
    Span12Mux_v I__2372 (
            .O(N__13229),
            .I(N__13226));
    Odrv12 I__2371 (
            .O(N__13226),
            .I(il_min_comp2_c));
    InMux I__2370 (
            .O(N__13223),
            .I(N__13220));
    LocalMux I__2369 (
            .O(N__13220),
            .I(il_max_comp1_D1));
    InMux I__2368 (
            .O(N__13217),
            .I(N__13213));
    InMux I__2367 (
            .O(N__13216),
            .I(N__13210));
    LocalMux I__2366 (
            .O(N__13213),
            .I(N__13205));
    LocalMux I__2365 (
            .O(N__13210),
            .I(N__13205));
    Span4Mux_h I__2364 (
            .O(N__13205),
            .I(N__13201));
    InMux I__2363 (
            .O(N__13204),
            .I(N__13198));
    Odrv4 I__2362 (
            .O(N__13201),
            .I(il_max_comp1_D2));
    LocalMux I__2361 (
            .O(N__13198),
            .I(il_max_comp1_D2));
    InMux I__2360 (
            .O(N__13193),
            .I(N__13190));
    LocalMux I__2359 (
            .O(N__13190),
            .I(N__13187));
    Odrv12 I__2358 (
            .O(N__13187),
            .I(\phase_controller_inst1.start_timer_hc_0_sqmuxa ));
    InMux I__2357 (
            .O(N__13184),
            .I(N__13181));
    LocalMux I__2356 (
            .O(N__13181),
            .I(N__13178));
    Span4Mux_v I__2355 (
            .O(N__13178),
            .I(N__13175));
    Sp12to4 I__2354 (
            .O(N__13175),
            .I(N__13172));
    Span12Mux_h I__2353 (
            .O(N__13172),
            .I(N__13169));
    Odrv12 I__2352 (
            .O(N__13169),
            .I(il_min_comp1_c));
    InMux I__2351 (
            .O(N__13166),
            .I(N__13163));
    LocalMux I__2350 (
            .O(N__13163),
            .I(il_min_comp1_D1));
    InMux I__2349 (
            .O(N__13160),
            .I(N__13154));
    InMux I__2348 (
            .O(N__13159),
            .I(N__13154));
    LocalMux I__2347 (
            .O(N__13154),
            .I(N__13151));
    Span4Mux_h I__2346 (
            .O(N__13151),
            .I(N__13147));
    InMux I__2345 (
            .O(N__13150),
            .I(N__13144));
    Odrv4 I__2344 (
            .O(N__13147),
            .I(il_min_comp1_D2));
    LocalMux I__2343 (
            .O(N__13144),
            .I(il_min_comp1_D2));
    InMux I__2342 (
            .O(N__13139),
            .I(N__13133));
    InMux I__2341 (
            .O(N__13138),
            .I(N__13133));
    LocalMux I__2340 (
            .O(N__13133),
            .I(N__13130));
    Odrv4 I__2339 (
            .O(N__13130),
            .I(\phase_controller_inst1.T01_0_sqmuxa ));
    InMux I__2338 (
            .O(N__13127),
            .I(N__13122));
    InMux I__2337 (
            .O(N__13126),
            .I(N__13119));
    InMux I__2336 (
            .O(N__13125),
            .I(N__13116));
    LocalMux I__2335 (
            .O(N__13122),
            .I(N__13113));
    LocalMux I__2334 (
            .O(N__13119),
            .I(\phase_controller_slave.tr_time_passed ));
    LocalMux I__2333 (
            .O(N__13116),
            .I(\phase_controller_slave.tr_time_passed ));
    Odrv4 I__2332 (
            .O(N__13113),
            .I(\phase_controller_slave.tr_time_passed ));
    InMux I__2331 (
            .O(N__13106),
            .I(N__13102));
    InMux I__2330 (
            .O(N__13105),
            .I(N__13099));
    LocalMux I__2329 (
            .O(N__13102),
            .I(\phase_controller_slave.stateZ0Z_0 ));
    LocalMux I__2328 (
            .O(N__13099),
            .I(\phase_controller_slave.stateZ0Z_0 ));
    InMux I__2327 (
            .O(N__13094),
            .I(N__13088));
    InMux I__2326 (
            .O(N__13093),
            .I(N__13088));
    LocalMux I__2325 (
            .O(N__13088),
            .I(\phase_controller_slave.state_RNIVDE2Z0Z_0 ));
    InMux I__2324 (
            .O(N__13085),
            .I(N__13078));
    InMux I__2323 (
            .O(N__13084),
            .I(N__13078));
    CascadeMux I__2322 (
            .O(N__13083),
            .I(N__13075));
    LocalMux I__2321 (
            .O(N__13078),
            .I(N__13072));
    InMux I__2320 (
            .O(N__13075),
            .I(N__13068));
    Span4Mux_s3_v I__2319 (
            .O(N__13072),
            .I(N__13065));
    InMux I__2318 (
            .O(N__13071),
            .I(N__13062));
    LocalMux I__2317 (
            .O(N__13068),
            .I(N__13059));
    Span4Mux_h I__2316 (
            .O(N__13065),
            .I(N__13052));
    LocalMux I__2315 (
            .O(N__13062),
            .I(N__13052));
    Span4Mux_v I__2314 (
            .O(N__13059),
            .I(N__13049));
    InMux I__2313 (
            .O(N__13058),
            .I(N__13046));
    InMux I__2312 (
            .O(N__13057),
            .I(N__13043));
    Sp12to4 I__2311 (
            .O(N__13052),
            .I(N__13040));
    Span4Mux_v I__2310 (
            .O(N__13049),
            .I(N__13035));
    LocalMux I__2309 (
            .O(N__13046),
            .I(N__13035));
    LocalMux I__2308 (
            .O(N__13043),
            .I(N__13032));
    Span12Mux_v I__2307 (
            .O(N__13040),
            .I(N__13025));
    Sp12to4 I__2306 (
            .O(N__13035),
            .I(N__13025));
    Sp12to4 I__2305 (
            .O(N__13032),
            .I(N__13025));
    Span12Mux_v I__2304 (
            .O(N__13025),
            .I(N__13022));
    Span12Mux_h I__2303 (
            .O(N__13022),
            .I(N__13019));
    Odrv12 I__2302 (
            .O(N__13019),
            .I(start_stop_c));
    CascadeMux I__2301 (
            .O(N__13016),
            .I(N__13011));
    InMux I__2300 (
            .O(N__13015),
            .I(N__13008));
    InMux I__2299 (
            .O(N__13014),
            .I(N__13005));
    InMux I__2298 (
            .O(N__13011),
            .I(N__13002));
    LocalMux I__2297 (
            .O(N__13008),
            .I(N__12997));
    LocalMux I__2296 (
            .O(N__13005),
            .I(N__12997));
    LocalMux I__2295 (
            .O(N__13002),
            .I(shift_flag_start));
    Odrv12 I__2294 (
            .O(N__12997),
            .I(shift_flag_start));
    InMux I__2293 (
            .O(N__12992),
            .I(N__12989));
    LocalMux I__2292 (
            .O(N__12989),
            .I(N__12986));
    Span12Mux_v I__2291 (
            .O(N__12986),
            .I(N__12983));
    Span12Mux_v I__2290 (
            .O(N__12983),
            .I(N__12980));
    Odrv12 I__2289 (
            .O(N__12980),
            .I(il_max_comp2_c));
    InMux I__2288 (
            .O(N__12977),
            .I(N__12974));
    LocalMux I__2287 (
            .O(N__12974),
            .I(il_max_comp2_D1));
    InMux I__2286 (
            .O(N__12971),
            .I(N__12968));
    LocalMux I__2285 (
            .O(N__12968),
            .I(N__12965));
    Odrv4 I__2284 (
            .O(N__12965),
            .I(\phase_controller_slave.state_RNO_0Z0Z_3 ));
    InMux I__2283 (
            .O(N__12962),
            .I(N__12955));
    InMux I__2282 (
            .O(N__12961),
            .I(N__12955));
    InMux I__2281 (
            .O(N__12960),
            .I(N__12952));
    LocalMux I__2280 (
            .O(N__12955),
            .I(il_max_comp2_D2));
    LocalMux I__2279 (
            .O(N__12952),
            .I(il_max_comp2_D2));
    InMux I__2278 (
            .O(N__12947),
            .I(N__12944));
    LocalMux I__2277 (
            .O(N__12944),
            .I(\phase_controller_slave.start_timer_hc_0_sqmuxa ));
    CascadeMux I__2276 (
            .O(N__12941),
            .I(N__12937));
    InMux I__2275 (
            .O(N__12940),
            .I(N__12931));
    InMux I__2274 (
            .O(N__12937),
            .I(N__12931));
    CascadeMux I__2273 (
            .O(N__12936),
            .I(N__12928));
    LocalMux I__2272 (
            .O(N__12931),
            .I(N__12924));
    InMux I__2271 (
            .O(N__12928),
            .I(N__12919));
    InMux I__2270 (
            .O(N__12927),
            .I(N__12919));
    Odrv4 I__2269 (
            .O(N__12924),
            .I(\phase_controller_slave.stateZ0Z_4 ));
    LocalMux I__2268 (
            .O(N__12919),
            .I(\phase_controller_slave.stateZ0Z_4 ));
    CascadeMux I__2267 (
            .O(N__12914),
            .I(N__12899));
    CascadeMux I__2266 (
            .O(N__12913),
            .I(N__12896));
    CascadeMux I__2265 (
            .O(N__12912),
            .I(N__12893));
    CascadeMux I__2264 (
            .O(N__12911),
            .I(N__12889));
    CascadeMux I__2263 (
            .O(N__12910),
            .I(N__12885));
    CascadeMux I__2262 (
            .O(N__12909),
            .I(N__12882));
    CascadeMux I__2261 (
            .O(N__12908),
            .I(N__12875));
    CascadeMux I__2260 (
            .O(N__12907),
            .I(N__12872));
    CascadeMux I__2259 (
            .O(N__12906),
            .I(N__12869));
    CascadeMux I__2258 (
            .O(N__12905),
            .I(N__12866));
    CascadeMux I__2257 (
            .O(N__12904),
            .I(N__12863));
    CascadeMux I__2256 (
            .O(N__12903),
            .I(N__12858));
    CascadeMux I__2255 (
            .O(N__12902),
            .I(N__12855));
    InMux I__2254 (
            .O(N__12899),
            .I(N__12844));
    InMux I__2253 (
            .O(N__12896),
            .I(N__12844));
    InMux I__2252 (
            .O(N__12893),
            .I(N__12844));
    InMux I__2251 (
            .O(N__12892),
            .I(N__12844));
    InMux I__2250 (
            .O(N__12889),
            .I(N__12835));
    InMux I__2249 (
            .O(N__12888),
            .I(N__12835));
    InMux I__2248 (
            .O(N__12885),
            .I(N__12835));
    InMux I__2247 (
            .O(N__12882),
            .I(N__12835));
    InMux I__2246 (
            .O(N__12881),
            .I(N__12818));
    InMux I__2245 (
            .O(N__12880),
            .I(N__12818));
    InMux I__2244 (
            .O(N__12879),
            .I(N__12818));
    InMux I__2243 (
            .O(N__12878),
            .I(N__12818));
    InMux I__2242 (
            .O(N__12875),
            .I(N__12818));
    InMux I__2241 (
            .O(N__12872),
            .I(N__12818));
    InMux I__2240 (
            .O(N__12869),
            .I(N__12818));
    InMux I__2239 (
            .O(N__12866),
            .I(N__12818));
    InMux I__2238 (
            .O(N__12863),
            .I(N__12813));
    InMux I__2237 (
            .O(N__12862),
            .I(N__12813));
    InMux I__2236 (
            .O(N__12861),
            .I(N__12810));
    InMux I__2235 (
            .O(N__12858),
            .I(N__12803));
    InMux I__2234 (
            .O(N__12855),
            .I(N__12803));
    InMux I__2233 (
            .O(N__12854),
            .I(N__12803));
    InMux I__2232 (
            .O(N__12853),
            .I(N__12800));
    LocalMux I__2231 (
            .O(N__12844),
            .I(N__12794));
    LocalMux I__2230 (
            .O(N__12835),
            .I(N__12794));
    LocalMux I__2229 (
            .O(N__12818),
            .I(N__12791));
    LocalMux I__2228 (
            .O(N__12813),
            .I(N__12786));
    LocalMux I__2227 (
            .O(N__12810),
            .I(N__12786));
    LocalMux I__2226 (
            .O(N__12803),
            .I(N__12783));
    LocalMux I__2225 (
            .O(N__12800),
            .I(N__12780));
    InMux I__2224 (
            .O(N__12799),
            .I(N__12777));
    Span4Mux_h I__2223 (
            .O(N__12794),
            .I(N__12774));
    Span4Mux_h I__2222 (
            .O(N__12791),
            .I(N__12769));
    Span4Mux_h I__2221 (
            .O(N__12786),
            .I(N__12769));
    Span4Mux_h I__2220 (
            .O(N__12783),
            .I(N__12764));
    Span4Mux_h I__2219 (
            .O(N__12780),
            .I(N__12764));
    LocalMux I__2218 (
            .O(N__12777),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    Odrv4 I__2217 (
            .O(N__12774),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    Odrv4 I__2216 (
            .O(N__12769),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    Odrv4 I__2215 (
            .O(N__12764),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    InMux I__2214 (
            .O(N__12755),
            .I(N__12752));
    LocalMux I__2213 (
            .O(N__12752),
            .I(N__12749));
    Odrv4 I__2212 (
            .O(N__12749),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_14 ));
    InMux I__2211 (
            .O(N__12746),
            .I(N__12743));
    LocalMux I__2210 (
            .O(N__12743),
            .I(N__12740));
    Odrv4 I__2209 (
            .O(N__12740),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_15 ));
    InMux I__2208 (
            .O(N__12737),
            .I(N__12728));
    InMux I__2207 (
            .O(N__12736),
            .I(N__12728));
    InMux I__2206 (
            .O(N__12735),
            .I(N__12728));
    LocalMux I__2205 (
            .O(N__12728),
            .I(N__12718));
    InMux I__2204 (
            .O(N__12727),
            .I(N__12707));
    InMux I__2203 (
            .O(N__12726),
            .I(N__12707));
    InMux I__2202 (
            .O(N__12725),
            .I(N__12707));
    InMux I__2201 (
            .O(N__12724),
            .I(N__12707));
    InMux I__2200 (
            .O(N__12723),
            .I(N__12707));
    InMux I__2199 (
            .O(N__12722),
            .I(N__12702));
    InMux I__2198 (
            .O(N__12721),
            .I(N__12702));
    Odrv4 I__2197 (
            .O(N__12718),
            .I(\phase_controller_inst1.stoper_tr.N_38 ));
    LocalMux I__2196 (
            .O(N__12707),
            .I(\phase_controller_inst1.stoper_tr.N_38 ));
    LocalMux I__2195 (
            .O(N__12702),
            .I(\phase_controller_inst1.stoper_tr.N_38 ));
    InMux I__2194 (
            .O(N__12695),
            .I(N__12692));
    LocalMux I__2193 (
            .O(N__12692),
            .I(N__12689));
    Odrv4 I__2192 (
            .O(N__12689),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_13 ));
    InMux I__2191 (
            .O(N__12686),
            .I(N__12683));
    LocalMux I__2190 (
            .O(N__12683),
            .I(N__12680));
    Odrv4 I__2189 (
            .O(N__12680),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_18 ));
    InMux I__2188 (
            .O(N__12677),
            .I(N__12674));
    LocalMux I__2187 (
            .O(N__12674),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_17 ));
    CEMux I__2186 (
            .O(N__12671),
            .I(N__12668));
    LocalMux I__2185 (
            .O(N__12668),
            .I(N__12663));
    CEMux I__2184 (
            .O(N__12667),
            .I(N__12660));
    CEMux I__2183 (
            .O(N__12666),
            .I(N__12657));
    Span4Mux_v I__2182 (
            .O(N__12663),
            .I(N__12652));
    LocalMux I__2181 (
            .O(N__12660),
            .I(N__12652));
    LocalMux I__2180 (
            .O(N__12657),
            .I(N__12649));
    Span4Mux_v I__2179 (
            .O(N__12652),
            .I(N__12646));
    Span4Mux_h I__2178 (
            .O(N__12649),
            .I(N__12641));
    Span4Mux_v I__2177 (
            .O(N__12646),
            .I(N__12641));
    Odrv4 I__2176 (
            .O(N__12641),
            .I(\phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ));
    InMux I__2175 (
            .O(N__12638),
            .I(N__12635));
    LocalMux I__2174 (
            .O(N__12635),
            .I(\phase_controller_slave.start_timer_tr_0_sqmuxa ));
    CascadeMux I__2173 (
            .O(N__12632),
            .I(N__12629));
    InMux I__2172 (
            .O(N__12629),
            .I(N__12626));
    LocalMux I__2171 (
            .O(N__12626),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_19 ));
    InMux I__2170 (
            .O(N__12623),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19 ));
    CascadeMux I__2169 (
            .O(N__12620),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_ ));
    InMux I__2168 (
            .O(N__12617),
            .I(N__12614));
    LocalMux I__2167 (
            .O(N__12614),
            .I(N__12611));
    Odrv4 I__2166 (
            .O(N__12611),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0 ));
    InMux I__2165 (
            .O(N__12608),
            .I(N__12605));
    LocalMux I__2164 (
            .O(N__12605),
            .I(N__12602));
    Odrv4 I__2163 (
            .O(N__12602),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_16 ));
    InMux I__2162 (
            .O(N__12599),
            .I(N__12596));
    LocalMux I__2161 (
            .O(N__12596),
            .I(N__12593));
    Odrv4 I__2160 (
            .O(N__12593),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_10 ));
    InMux I__2159 (
            .O(N__12590),
            .I(N__12587));
    LocalMux I__2158 (
            .O(N__12587),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_19 ));
    InMux I__2157 (
            .O(N__12584),
            .I(N__12581));
    LocalMux I__2156 (
            .O(N__12581),
            .I(N__12578));
    Odrv4 I__2155 (
            .O(N__12578),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_11 ));
    CascadeMux I__2154 (
            .O(N__12575),
            .I(N__12572));
    InMux I__2153 (
            .O(N__12572),
            .I(N__12569));
    LocalMux I__2152 (
            .O(N__12569),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_11 ));
    InMux I__2151 (
            .O(N__12566),
            .I(N__12563));
    LocalMux I__2150 (
            .O(N__12563),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_12 ));
    CascadeMux I__2149 (
            .O(N__12560),
            .I(N__12557));
    InMux I__2148 (
            .O(N__12557),
            .I(N__12554));
    LocalMux I__2147 (
            .O(N__12554),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_12 ));
    CascadeMux I__2146 (
            .O(N__12551),
            .I(N__12548));
    InMux I__2145 (
            .O(N__12548),
            .I(N__12545));
    LocalMux I__2144 (
            .O(N__12545),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_13 ));
    CascadeMux I__2143 (
            .O(N__12542),
            .I(N__12539));
    InMux I__2142 (
            .O(N__12539),
            .I(N__12536));
    LocalMux I__2141 (
            .O(N__12536),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_14 ));
    CascadeMux I__2140 (
            .O(N__12533),
            .I(N__12530));
    InMux I__2139 (
            .O(N__12530),
            .I(N__12527));
    LocalMux I__2138 (
            .O(N__12527),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_15 ));
    CascadeMux I__2137 (
            .O(N__12524),
            .I(N__12521));
    InMux I__2136 (
            .O(N__12521),
            .I(N__12518));
    LocalMux I__2135 (
            .O(N__12518),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_16 ));
    CascadeMux I__2134 (
            .O(N__12515),
            .I(N__12512));
    InMux I__2133 (
            .O(N__12512),
            .I(N__12509));
    LocalMux I__2132 (
            .O(N__12509),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_17 ));
    CascadeMux I__2131 (
            .O(N__12506),
            .I(N__12503));
    InMux I__2130 (
            .O(N__12503),
            .I(N__12500));
    LocalMux I__2129 (
            .O(N__12500),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_18 ));
    InMux I__2128 (
            .O(N__12497),
            .I(N__12494));
    LocalMux I__2127 (
            .O(N__12494),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__2126 (
            .O(N__12491),
            .I(N__12488));
    InMux I__2125 (
            .O(N__12488),
            .I(N__12485));
    LocalMux I__2124 (
            .O(N__12485),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_3 ));
    InMux I__2123 (
            .O(N__12482),
            .I(N__12479));
    LocalMux I__2122 (
            .O(N__12479),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_4 ));
    CascadeMux I__2121 (
            .O(N__12476),
            .I(N__12473));
    InMux I__2120 (
            .O(N__12473),
            .I(N__12470));
    LocalMux I__2119 (
            .O(N__12470),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_4 ));
    InMux I__2118 (
            .O(N__12467),
            .I(N__12464));
    LocalMux I__2117 (
            .O(N__12464),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_5 ));
    CascadeMux I__2116 (
            .O(N__12461),
            .I(N__12458));
    InMux I__2115 (
            .O(N__12458),
            .I(N__12455));
    LocalMux I__2114 (
            .O(N__12455),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_5 ));
    InMux I__2113 (
            .O(N__12452),
            .I(N__12449));
    LocalMux I__2112 (
            .O(N__12449),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__2111 (
            .O(N__12446),
            .I(N__12443));
    InMux I__2110 (
            .O(N__12443),
            .I(N__12440));
    LocalMux I__2109 (
            .O(N__12440),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_6 ));
    InMux I__2108 (
            .O(N__12437),
            .I(N__12434));
    LocalMux I__2107 (
            .O(N__12434),
            .I(N__12431));
    Odrv4 I__2106 (
            .O(N__12431),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_7 ));
    CascadeMux I__2105 (
            .O(N__12428),
            .I(N__12425));
    InMux I__2104 (
            .O(N__12425),
            .I(N__12422));
    LocalMux I__2103 (
            .O(N__12422),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_7 ));
    InMux I__2102 (
            .O(N__12419),
            .I(N__12416));
    LocalMux I__2101 (
            .O(N__12416),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__2100 (
            .O(N__12413),
            .I(N__12410));
    InMux I__2099 (
            .O(N__12410),
            .I(N__12407));
    LocalMux I__2098 (
            .O(N__12407),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_8 ));
    InMux I__2097 (
            .O(N__12404),
            .I(N__12401));
    LocalMux I__2096 (
            .O(N__12401),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_9 ));
    CascadeMux I__2095 (
            .O(N__12398),
            .I(N__12395));
    InMux I__2094 (
            .O(N__12395),
            .I(N__12392));
    LocalMux I__2093 (
            .O(N__12392),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_9 ));
    CascadeMux I__2092 (
            .O(N__12389),
            .I(N__12386));
    InMux I__2091 (
            .O(N__12386),
            .I(N__12383));
    LocalMux I__2090 (
            .O(N__12383),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_10 ));
    InMux I__2089 (
            .O(N__12380),
            .I(N__12375));
    InMux I__2088 (
            .O(N__12379),
            .I(N__12372));
    InMux I__2087 (
            .O(N__12378),
            .I(N__12369));
    LocalMux I__2086 (
            .O(N__12375),
            .I(N__12364));
    LocalMux I__2085 (
            .O(N__12372),
            .I(N__12364));
    LocalMux I__2084 (
            .O(N__12369),
            .I(\phase_controller_inst1.tr_time_passed ));
    Odrv4 I__2083 (
            .O(N__12364),
            .I(\phase_controller_inst1.tr_time_passed ));
    InMux I__2082 (
            .O(N__12359),
            .I(N__12355));
    InMux I__2081 (
            .O(N__12358),
            .I(N__12352));
    LocalMux I__2080 (
            .O(N__12355),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    LocalMux I__2079 (
            .O(N__12352),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    InMux I__2078 (
            .O(N__12347),
            .I(N__12341));
    InMux I__2077 (
            .O(N__12346),
            .I(N__12341));
    LocalMux I__2076 (
            .O(N__12341),
            .I(N__12336));
    InMux I__2075 (
            .O(N__12340),
            .I(N__12333));
    InMux I__2074 (
            .O(N__12339),
            .I(N__12330));
    Odrv4 I__2073 (
            .O(N__12336),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__2072 (
            .O(N__12333),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__2071 (
            .O(N__12330),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    InMux I__2070 (
            .O(N__12323),
            .I(N__12318));
    InMux I__2069 (
            .O(N__12322),
            .I(N__12315));
    InMux I__2068 (
            .O(N__12321),
            .I(N__12311));
    LocalMux I__2067 (
            .O(N__12318),
            .I(N__12308));
    LocalMux I__2066 (
            .O(N__12315),
            .I(N__12305));
    InMux I__2065 (
            .O(N__12314),
            .I(N__12302));
    LocalMux I__2064 (
            .O(N__12311),
            .I(N__12295));
    Span4Mux_v I__2063 (
            .O(N__12308),
            .I(N__12295));
    Span4Mux_h I__2062 (
            .O(N__12305),
            .I(N__12295));
    LocalMux I__2061 (
            .O(N__12302),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv4 I__2060 (
            .O(N__12295),
            .I(\phase_controller_inst1.hc_time_passed ));
    CascadeMux I__2059 (
            .O(N__12290),
            .I(N__12287));
    InMux I__2058 (
            .O(N__12287),
            .I(N__12281));
    InMux I__2057 (
            .O(N__12286),
            .I(N__12278));
    InMux I__2056 (
            .O(N__12285),
            .I(N__12272));
    InMux I__2055 (
            .O(N__12284),
            .I(N__12272));
    LocalMux I__2054 (
            .O(N__12281),
            .I(N__12267));
    LocalMux I__2053 (
            .O(N__12278),
            .I(N__12267));
    InMux I__2052 (
            .O(N__12277),
            .I(N__12264));
    LocalMux I__2051 (
            .O(N__12272),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    Odrv4 I__2050 (
            .O(N__12267),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    LocalMux I__2049 (
            .O(N__12264),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    InMux I__2048 (
            .O(N__12257),
            .I(N__12253));
    InMux I__2047 (
            .O(N__12256),
            .I(N__12250));
    LocalMux I__2046 (
            .O(N__12253),
            .I(\phase_controller_inst1.N_107 ));
    LocalMux I__2045 (
            .O(N__12250),
            .I(\phase_controller_inst1.N_107 ));
    CascadeMux I__2044 (
            .O(N__12245),
            .I(N__12238));
    CascadeMux I__2043 (
            .O(N__12244),
            .I(N__12235));
    CascadeMux I__2042 (
            .O(N__12243),
            .I(N__12232));
    CascadeMux I__2041 (
            .O(N__12242),
            .I(N__12217));
    CascadeMux I__2040 (
            .O(N__12241),
            .I(N__12214));
    InMux I__2039 (
            .O(N__12238),
            .I(N__12199));
    InMux I__2038 (
            .O(N__12235),
            .I(N__12199));
    InMux I__2037 (
            .O(N__12232),
            .I(N__12199));
    InMux I__2036 (
            .O(N__12231),
            .I(N__12199));
    InMux I__2035 (
            .O(N__12230),
            .I(N__12199));
    InMux I__2034 (
            .O(N__12229),
            .I(N__12199));
    InMux I__2033 (
            .O(N__12228),
            .I(N__12199));
    CascadeMux I__2032 (
            .O(N__12227),
            .I(N__12196));
    CascadeMux I__2031 (
            .O(N__12226),
            .I(N__12193));
    CascadeMux I__2030 (
            .O(N__12225),
            .I(N__12190));
    CascadeMux I__2029 (
            .O(N__12224),
            .I(N__12187));
    CascadeMux I__2028 (
            .O(N__12223),
            .I(N__12180));
    CascadeMux I__2027 (
            .O(N__12222),
            .I(N__12177));
    CascadeMux I__2026 (
            .O(N__12221),
            .I(N__12174));
    CascadeMux I__2025 (
            .O(N__12220),
            .I(N__12171));
    InMux I__2024 (
            .O(N__12217),
            .I(N__12164));
    InMux I__2023 (
            .O(N__12214),
            .I(N__12164));
    LocalMux I__2022 (
            .O(N__12199),
            .I(N__12161));
    InMux I__2021 (
            .O(N__12196),
            .I(N__12144));
    InMux I__2020 (
            .O(N__12193),
            .I(N__12144));
    InMux I__2019 (
            .O(N__12190),
            .I(N__12144));
    InMux I__2018 (
            .O(N__12187),
            .I(N__12144));
    InMux I__2017 (
            .O(N__12186),
            .I(N__12144));
    InMux I__2016 (
            .O(N__12185),
            .I(N__12144));
    InMux I__2015 (
            .O(N__12184),
            .I(N__12144));
    InMux I__2014 (
            .O(N__12183),
            .I(N__12144));
    InMux I__2013 (
            .O(N__12180),
            .I(N__12137));
    InMux I__2012 (
            .O(N__12177),
            .I(N__12137));
    InMux I__2011 (
            .O(N__12174),
            .I(N__12137));
    InMux I__2010 (
            .O(N__12171),
            .I(N__12134));
    InMux I__2009 (
            .O(N__12170),
            .I(N__12131));
    InMux I__2008 (
            .O(N__12169),
            .I(N__12128));
    LocalMux I__2007 (
            .O(N__12164),
            .I(N__12124));
    Sp12to4 I__2006 (
            .O(N__12161),
            .I(N__12115));
    LocalMux I__2005 (
            .O(N__12144),
            .I(N__12115));
    LocalMux I__2004 (
            .O(N__12137),
            .I(N__12115));
    LocalMux I__2003 (
            .O(N__12134),
            .I(N__12115));
    LocalMux I__2002 (
            .O(N__12131),
            .I(N__12110));
    LocalMux I__2001 (
            .O(N__12128),
            .I(N__12110));
    InMux I__2000 (
            .O(N__12127),
            .I(N__12107));
    Span4Mux_h I__1999 (
            .O(N__12124),
            .I(N__12104));
    Span12Mux_v I__1998 (
            .O(N__12115),
            .I(N__12101));
    Span4Mux_h I__1997 (
            .O(N__12110),
            .I(N__12098));
    LocalMux I__1996 (
            .O(N__12107),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__1995 (
            .O(N__12104),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv12 I__1994 (
            .O(N__12101),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__1993 (
            .O(N__12098),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    InMux I__1992 (
            .O(N__12089),
            .I(N__12086));
    LocalMux I__1991 (
            .O(N__12086),
            .I(N__12083));
    Odrv4 I__1990 (
            .O(N__12083),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__1989 (
            .O(N__12080),
            .I(N__12077));
    InMux I__1988 (
            .O(N__12077),
            .I(N__12074));
    LocalMux I__1987 (
            .O(N__12074),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_1 ));
    InMux I__1986 (
            .O(N__12071),
            .I(N__12068));
    LocalMux I__1985 (
            .O(N__12068),
            .I(N__12065));
    Span4Mux_h I__1984 (
            .O(N__12065),
            .I(N__12062));
    Odrv4 I__1983 (
            .O(N__12062),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_2 ));
    CascadeMux I__1982 (
            .O(N__12059),
            .I(N__12056));
    InMux I__1981 (
            .O(N__12056),
            .I(N__12053));
    LocalMux I__1980 (
            .O(N__12053),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_2 ));
    InMux I__1979 (
            .O(N__12050),
            .I(N__12047));
    LocalMux I__1978 (
            .O(N__12047),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_18 ));
    CEMux I__1977 (
            .O(N__12044),
            .I(N__12039));
    CEMux I__1976 (
            .O(N__12043),
            .I(N__12036));
    CEMux I__1975 (
            .O(N__12042),
            .I(N__12032));
    LocalMux I__1974 (
            .O(N__12039),
            .I(N__12027));
    LocalMux I__1973 (
            .O(N__12036),
            .I(N__12027));
    CEMux I__1972 (
            .O(N__12035),
            .I(N__12024));
    LocalMux I__1971 (
            .O(N__12032),
            .I(N__12021));
    Span4Mux_v I__1970 (
            .O(N__12027),
            .I(N__12016));
    LocalMux I__1969 (
            .O(N__12024),
            .I(N__12016));
    Span4Mux_h I__1968 (
            .O(N__12021),
            .I(N__12013));
    Span4Mux_v I__1967 (
            .O(N__12016),
            .I(N__12010));
    Span4Mux_s3_h I__1966 (
            .O(N__12013),
            .I(N__12007));
    Span4Mux_s0_v I__1965 (
            .O(N__12010),
            .I(N__12004));
    Odrv4 I__1964 (
            .O(N__12007),
            .I(\phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__1963 (
            .O(N__12004),
            .I(\phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ));
    InMux I__1962 (
            .O(N__11999),
            .I(N__11996));
    LocalMux I__1961 (
            .O(N__11996),
            .I(N__11993));
    Span4Mux_h I__1960 (
            .O(N__11993),
            .I(N__11988));
    InMux I__1959 (
            .O(N__11992),
            .I(N__11985));
    InMux I__1958 (
            .O(N__11991),
            .I(N__11982));
    Odrv4 I__1957 (
            .O(N__11988),
            .I(\phase_controller_slave.stoper_hc.time_passed11 ));
    LocalMux I__1956 (
            .O(N__11985),
            .I(\phase_controller_slave.stoper_hc.time_passed11 ));
    LocalMux I__1955 (
            .O(N__11982),
            .I(\phase_controller_slave.stoper_hc.time_passed11 ));
    CascadeMux I__1954 (
            .O(N__11975),
            .I(N__11972));
    InMux I__1953 (
            .O(N__11972),
            .I(N__11969));
    LocalMux I__1952 (
            .O(N__11969),
            .I(\phase_controller_slave.stoper_hc.time_passed_1_sqmuxa ));
    InMux I__1951 (
            .O(N__11966),
            .I(N__11959));
    InMux I__1950 (
            .O(N__11965),
            .I(N__11954));
    InMux I__1949 (
            .O(N__11964),
            .I(N__11954));
    InMux I__1948 (
            .O(N__11963),
            .I(N__11949));
    InMux I__1947 (
            .O(N__11962),
            .I(N__11949));
    LocalMux I__1946 (
            .O(N__11959),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__1945 (
            .O(N__11954),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__1944 (
            .O(N__11949),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__1943 (
            .O(N__11942),
            .I(N__11929));
    CascadeMux I__1942 (
            .O(N__11941),
            .I(N__11925));
    CascadeMux I__1941 (
            .O(N__11940),
            .I(N__11922));
    CascadeMux I__1940 (
            .O(N__11939),
            .I(N__11919));
    CascadeMux I__1939 (
            .O(N__11938),
            .I(N__11916));
    CascadeMux I__1938 (
            .O(N__11937),
            .I(N__11908));
    CascadeMux I__1937 (
            .O(N__11936),
            .I(N__11905));
    CascadeMux I__1936 (
            .O(N__11935),
            .I(N__11898));
    CascadeMux I__1935 (
            .O(N__11934),
            .I(N__11895));
    CascadeMux I__1934 (
            .O(N__11933),
            .I(N__11892));
    CascadeMux I__1933 (
            .O(N__11932),
            .I(N__11889));
    InMux I__1932 (
            .O(N__11929),
            .I(N__11883));
    InMux I__1931 (
            .O(N__11928),
            .I(N__11883));
    InMux I__1930 (
            .O(N__11925),
            .I(N__11866));
    InMux I__1929 (
            .O(N__11922),
            .I(N__11866));
    InMux I__1928 (
            .O(N__11919),
            .I(N__11866));
    InMux I__1927 (
            .O(N__11916),
            .I(N__11866));
    InMux I__1926 (
            .O(N__11915),
            .I(N__11866));
    InMux I__1925 (
            .O(N__11914),
            .I(N__11866));
    InMux I__1924 (
            .O(N__11913),
            .I(N__11866));
    InMux I__1923 (
            .O(N__11912),
            .I(N__11861));
    InMux I__1922 (
            .O(N__11911),
            .I(N__11861));
    InMux I__1921 (
            .O(N__11908),
            .I(N__11856));
    InMux I__1920 (
            .O(N__11905),
            .I(N__11856));
    InMux I__1919 (
            .O(N__11904),
            .I(N__11839));
    InMux I__1918 (
            .O(N__11903),
            .I(N__11839));
    InMux I__1917 (
            .O(N__11902),
            .I(N__11839));
    InMux I__1916 (
            .O(N__11901),
            .I(N__11839));
    InMux I__1915 (
            .O(N__11898),
            .I(N__11839));
    InMux I__1914 (
            .O(N__11895),
            .I(N__11839));
    InMux I__1913 (
            .O(N__11892),
            .I(N__11839));
    InMux I__1912 (
            .O(N__11889),
            .I(N__11839));
    CascadeMux I__1911 (
            .O(N__11888),
            .I(N__11836));
    LocalMux I__1910 (
            .O(N__11883),
            .I(N__11833));
    InMux I__1909 (
            .O(N__11882),
            .I(N__11828));
    InMux I__1908 (
            .O(N__11881),
            .I(N__11828));
    LocalMux I__1907 (
            .O(N__11866),
            .I(N__11825));
    LocalMux I__1906 (
            .O(N__11861),
            .I(N__11820));
    LocalMux I__1905 (
            .O(N__11856),
            .I(N__11820));
    LocalMux I__1904 (
            .O(N__11839),
            .I(N__11817));
    InMux I__1903 (
            .O(N__11836),
            .I(N__11814));
    Span4Mux_v I__1902 (
            .O(N__11833),
            .I(N__11809));
    LocalMux I__1901 (
            .O(N__11828),
            .I(N__11809));
    Span4Mux_h I__1900 (
            .O(N__11825),
            .I(N__11806));
    Span4Mux_h I__1899 (
            .O(N__11820),
            .I(N__11803));
    Span4Mux_h I__1898 (
            .O(N__11817),
            .I(N__11800));
    LocalMux I__1897 (
            .O(N__11814),
            .I(N__11795));
    Span4Mux_v I__1896 (
            .O(N__11809),
            .I(N__11795));
    Odrv4 I__1895 (
            .O(N__11806),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__1894 (
            .O(N__11803),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__1893 (
            .O(N__11800),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__1892 (
            .O(N__11795),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    InMux I__1891 (
            .O(N__11786),
            .I(N__11783));
    LocalMux I__1890 (
            .O(N__11783),
            .I(N__11780));
    Odrv4 I__1889 (
            .O(N__11780),
            .I(\phase_controller_inst1.N_110 ));
    InMux I__1888 (
            .O(N__11777),
            .I(N__11774));
    LocalMux I__1887 (
            .O(N__11774),
            .I(\phase_controller_inst1.N_112 ));
    InMux I__1886 (
            .O(N__11771),
            .I(N__11768));
    LocalMux I__1885 (
            .O(N__11768),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_13 ));
    InMux I__1884 (
            .O(N__11765),
            .I(N__11762));
    LocalMux I__1883 (
            .O(N__11762),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_10 ));
    InMux I__1882 (
            .O(N__11759),
            .I(N__11756));
    LocalMux I__1881 (
            .O(N__11756),
            .I(N__11753));
    Odrv4 I__1880 (
            .O(N__11753),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_12 ));
    InMux I__1879 (
            .O(N__11750),
            .I(N__11746));
    InMux I__1878 (
            .O(N__11749),
            .I(N__11743));
    LocalMux I__1877 (
            .O(N__11746),
            .I(N__11739));
    LocalMux I__1876 (
            .O(N__11743),
            .I(N__11736));
    InMux I__1875 (
            .O(N__11742),
            .I(N__11733));
    Odrv12 I__1874 (
            .O(N__11739),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_0Z0Z_6 ));
    Odrv4 I__1873 (
            .O(N__11736),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_0Z0Z_6 ));
    LocalMux I__1872 (
            .O(N__11733),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_0Z0Z_6 ));
    InMux I__1871 (
            .O(N__11726),
            .I(N__11723));
    LocalMux I__1870 (
            .O(N__11723),
            .I(N__11720));
    Span12Mux_s5_v I__1869 (
            .O(N__11720),
            .I(N__11717));
    Odrv12 I__1868 (
            .O(N__11717),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_9 ));
    CascadeMux I__1867 (
            .O(N__11714),
            .I(N__11709));
    CascadeMux I__1866 (
            .O(N__11713),
            .I(N__11703));
    InMux I__1865 (
            .O(N__11712),
            .I(N__11696));
    InMux I__1864 (
            .O(N__11709),
            .I(N__11687));
    InMux I__1863 (
            .O(N__11708),
            .I(N__11687));
    InMux I__1862 (
            .O(N__11707),
            .I(N__11687));
    InMux I__1861 (
            .O(N__11706),
            .I(N__11687));
    InMux I__1860 (
            .O(N__11703),
            .I(N__11676));
    InMux I__1859 (
            .O(N__11702),
            .I(N__11676));
    InMux I__1858 (
            .O(N__11701),
            .I(N__11676));
    InMux I__1857 (
            .O(N__11700),
            .I(N__11676));
    InMux I__1856 (
            .O(N__11699),
            .I(N__11676));
    LocalMux I__1855 (
            .O(N__11696),
            .I(N__11671));
    LocalMux I__1854 (
            .O(N__11687),
            .I(N__11671));
    LocalMux I__1853 (
            .O(N__11676),
            .I(N__11668));
    Odrv12 I__1852 (
            .O(N__11671),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2Z0Z_9 ));
    Odrv4 I__1851 (
            .O(N__11668),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2Z0Z_9 ));
    InMux I__1850 (
            .O(N__11663),
            .I(N__11660));
    LocalMux I__1849 (
            .O(N__11660),
            .I(N__11657));
    Span4Mux_v I__1848 (
            .O(N__11657),
            .I(N__11654));
    Odrv4 I__1847 (
            .O(N__11654),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_11 ));
    InMux I__1846 (
            .O(N__11651),
            .I(N__11645));
    InMux I__1845 (
            .O(N__11650),
            .I(N__11645));
    LocalMux I__1844 (
            .O(N__11645),
            .I(N__11640));
    InMux I__1843 (
            .O(N__11644),
            .I(N__11635));
    InMux I__1842 (
            .O(N__11643),
            .I(N__11635));
    Sp12to4 I__1841 (
            .O(N__11640),
            .I(N__11631));
    LocalMux I__1840 (
            .O(N__11635),
            .I(N__11628));
    InMux I__1839 (
            .O(N__11634),
            .I(N__11625));
    Odrv12 I__1838 (
            .O(N__11631),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_i_o2Z0Z_15 ));
    Odrv12 I__1837 (
            .O(N__11628),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_i_o2Z0Z_15 ));
    LocalMux I__1836 (
            .O(N__11625),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_i_o2Z0Z_15 ));
    InMux I__1835 (
            .O(N__11618),
            .I(N__11615));
    LocalMux I__1834 (
            .O(N__11615),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_14 ));
    InMux I__1833 (
            .O(N__11612),
            .I(N__11609));
    LocalMux I__1832 (
            .O(N__11609),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_16 ));
    InMux I__1831 (
            .O(N__11606),
            .I(N__11603));
    LocalMux I__1830 (
            .O(N__11603),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_19 ));
    InMux I__1829 (
            .O(N__11600),
            .I(N__11597));
    LocalMux I__1828 (
            .O(N__11597),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_17 ));
    InMux I__1827 (
            .O(N__11594),
            .I(N__11591));
    LocalMux I__1826 (
            .O(N__11591),
            .I(N__11588));
    Span4Mux_h I__1825 (
            .O(N__11588),
            .I(N__11585));
    Odrv4 I__1824 (
            .O(N__11585),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_5 ));
    InMux I__1823 (
            .O(N__11582),
            .I(N__11579));
    LocalMux I__1822 (
            .O(N__11579),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_1 ));
    InMux I__1821 (
            .O(N__11576),
            .I(N__11573));
    LocalMux I__1820 (
            .O(N__11573),
            .I(N__11570));
    Span4Mux_h I__1819 (
            .O(N__11570),
            .I(N__11567));
    Odrv4 I__1818 (
            .O(N__11567),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_7 ));
    InMux I__1817 (
            .O(N__11564),
            .I(N__11561));
    LocalMux I__1816 (
            .O(N__11561),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_6 ));
    InMux I__1815 (
            .O(N__11558),
            .I(N__11550));
    InMux I__1814 (
            .O(N__11557),
            .I(N__11550));
    InMux I__1813 (
            .O(N__11556),
            .I(N__11545));
    InMux I__1812 (
            .O(N__11555),
            .I(N__11545));
    LocalMux I__1811 (
            .O(N__11550),
            .I(N__11542));
    LocalMux I__1810 (
            .O(N__11545),
            .I(N__11539));
    Odrv12 I__1809 (
            .O(N__11542),
            .I(\phase_controller_inst1.stoper_hc.N_122 ));
    Odrv4 I__1808 (
            .O(N__11539),
            .I(\phase_controller_inst1.stoper_hc.N_122 ));
    CascadeMux I__1807 (
            .O(N__11534),
            .I(N__11531));
    InMux I__1806 (
            .O(N__11531),
            .I(N__11528));
    LocalMux I__1805 (
            .O(N__11528),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_2 ));
    InMux I__1804 (
            .O(N__11525),
            .I(N__11522));
    LocalMux I__1803 (
            .O(N__11522),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_4 ));
    InMux I__1802 (
            .O(N__11519),
            .I(N__11501));
    InMux I__1801 (
            .O(N__11518),
            .I(N__11501));
    InMux I__1800 (
            .O(N__11517),
            .I(N__11501));
    InMux I__1799 (
            .O(N__11516),
            .I(N__11501));
    InMux I__1798 (
            .O(N__11515),
            .I(N__11501));
    InMux I__1797 (
            .O(N__11514),
            .I(N__11501));
    LocalMux I__1796 (
            .O(N__11501),
            .I(N__11498));
    Span4Mux_v I__1795 (
            .O(N__11498),
            .I(N__11495));
    Span4Mux_v I__1794 (
            .O(N__11495),
            .I(N__11486));
    InMux I__1793 (
            .O(N__11494),
            .I(N__11473));
    InMux I__1792 (
            .O(N__11493),
            .I(N__11473));
    InMux I__1791 (
            .O(N__11492),
            .I(N__11473));
    InMux I__1790 (
            .O(N__11491),
            .I(N__11473));
    InMux I__1789 (
            .O(N__11490),
            .I(N__11473));
    InMux I__1788 (
            .O(N__11489),
            .I(N__11473));
    Odrv4 I__1787 (
            .O(N__11486),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a3_0Z0Z_6 ));
    LocalMux I__1786 (
            .O(N__11473),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a3_0Z0Z_6 ));
    InMux I__1785 (
            .O(N__11468),
            .I(N__11464));
    InMux I__1784 (
            .O(N__11467),
            .I(N__11461));
    LocalMux I__1783 (
            .O(N__11464),
            .I(N__11458));
    LocalMux I__1782 (
            .O(N__11461),
            .I(N__11455));
    Odrv12 I__1781 (
            .O(N__11458),
            .I(\phase_controller_inst1.stoper_hc.N_144 ));
    Odrv4 I__1780 (
            .O(N__11455),
            .I(\phase_controller_inst1.stoper_hc.N_144 ));
    InMux I__1779 (
            .O(N__11450),
            .I(N__11447));
    LocalMux I__1778 (
            .O(N__11447),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_3 ));
    CascadeMux I__1777 (
            .O(N__11444),
            .I(N__11435));
    InMux I__1776 (
            .O(N__11443),
            .I(N__11429));
    InMux I__1775 (
            .O(N__11442),
            .I(N__11429));
    InMux I__1774 (
            .O(N__11441),
            .I(N__11416));
    InMux I__1773 (
            .O(N__11440),
            .I(N__11416));
    InMux I__1772 (
            .O(N__11439),
            .I(N__11416));
    InMux I__1771 (
            .O(N__11438),
            .I(N__11416));
    InMux I__1770 (
            .O(N__11435),
            .I(N__11416));
    InMux I__1769 (
            .O(N__11434),
            .I(N__11416));
    LocalMux I__1768 (
            .O(N__11429),
            .I(N__11409));
    LocalMux I__1767 (
            .O(N__11416),
            .I(N__11409));
    CascadeMux I__1766 (
            .O(N__11415),
            .I(N__11405));
    CascadeMux I__1765 (
            .O(N__11414),
            .I(N__11398));
    Span4Mux_v I__1764 (
            .O(N__11409),
            .I(N__11394));
    InMux I__1763 (
            .O(N__11408),
            .I(N__11377));
    InMux I__1762 (
            .O(N__11405),
            .I(N__11377));
    InMux I__1761 (
            .O(N__11404),
            .I(N__11377));
    InMux I__1760 (
            .O(N__11403),
            .I(N__11377));
    InMux I__1759 (
            .O(N__11402),
            .I(N__11377));
    InMux I__1758 (
            .O(N__11401),
            .I(N__11377));
    InMux I__1757 (
            .O(N__11398),
            .I(N__11377));
    InMux I__1756 (
            .O(N__11397),
            .I(N__11377));
    Span4Mux_v I__1755 (
            .O(N__11394),
            .I(N__11372));
    LocalMux I__1754 (
            .O(N__11377),
            .I(N__11372));
    Odrv4 I__1753 (
            .O(N__11372),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2Z0Z_6 ));
    InMux I__1752 (
            .O(N__11369),
            .I(N__11366));
    LocalMux I__1751 (
            .O(N__11366),
            .I(N__11363));
    Odrv4 I__1750 (
            .O(N__11363),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_8 ));
    InMux I__1749 (
            .O(N__11360),
            .I(N__11357));
    LocalMux I__1748 (
            .O(N__11357),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_15 ));
    InMux I__1747 (
            .O(N__11354),
            .I(N__11351));
    LocalMux I__1746 (
            .O(N__11351),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_4Z0Z_3 ));
    CascadeMux I__1745 (
            .O(N__11348),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_3Z0Z_3_cascade_ ));
    CascadeMux I__1744 (
            .O(N__11345),
            .I(\phase_controller_inst1.stoper_hc.N_144_cascade_ ));
    CascadeMux I__1743 (
            .O(N__11342),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_0Z0Z_6_cascade_ ));
    InMux I__1742 (
            .O(N__11339),
            .I(N__11336));
    LocalMux I__1741 (
            .O(N__11336),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2Z0Z_9 ));
    CascadeMux I__1740 (
            .O(N__11333),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2Z0Z_9_cascade_ ));
    CascadeMux I__1739 (
            .O(N__11330),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_i_o2Z0Z_15_cascade_ ));
    InMux I__1738 (
            .O(N__11327),
            .I(N__11324));
    LocalMux I__1737 (
            .O(N__11324),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_1Z0Z_6 ));
    CascadeMux I__1736 (
            .O(N__11321),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_ ));
    InMux I__1735 (
            .O(N__11318),
            .I(N__11315));
    LocalMux I__1734 (
            .O(N__11315),
            .I(N__11312));
    Odrv4 I__1733 (
            .O(N__11312),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ));
    InMux I__1732 (
            .O(N__11309),
            .I(N__11306));
    LocalMux I__1731 (
            .O(N__11306),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ));
    InMux I__1730 (
            .O(N__11303),
            .I(N__11300));
    LocalMux I__1729 (
            .O(N__11300),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ));
    InMux I__1728 (
            .O(N__11297),
            .I(N__11294));
    LocalMux I__1727 (
            .O(N__11294),
            .I(N__11291));
    Odrv4 I__1726 (
            .O(N__11291),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ));
    InMux I__1725 (
            .O(N__11288),
            .I(N__11285));
    LocalMux I__1724 (
            .O(N__11285),
            .I(N__11282));
    Odrv4 I__1723 (
            .O(N__11282),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ));
    InMux I__1722 (
            .O(N__11279),
            .I(N__11276));
    LocalMux I__1721 (
            .O(N__11276),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ));
    CEMux I__1720 (
            .O(N__11273),
            .I(N__11270));
    LocalMux I__1719 (
            .O(N__11270),
            .I(N__11266));
    CEMux I__1718 (
            .O(N__11269),
            .I(N__11263));
    Span4Mux_v I__1717 (
            .O(N__11266),
            .I(N__11259));
    LocalMux I__1716 (
            .O(N__11263),
            .I(N__11256));
    CEMux I__1715 (
            .O(N__11262),
            .I(N__11253));
    Span4Mux_h I__1714 (
            .O(N__11259),
            .I(N__11250));
    Span4Mux_h I__1713 (
            .O(N__11256),
            .I(N__11247));
    LocalMux I__1712 (
            .O(N__11253),
            .I(N__11244));
    Odrv4 I__1711 (
            .O(N__11250),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__1710 (
            .O(N__11247),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv12 I__1709 (
            .O(N__11244),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    InMux I__1708 (
            .O(N__11237),
            .I(N__11234));
    LocalMux I__1707 (
            .O(N__11234),
            .I(N__11231));
    Odrv4 I__1706 (
            .O(N__11231),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ));
    InMux I__1705 (
            .O(N__11228),
            .I(N__11225));
    LocalMux I__1704 (
            .O(N__11225),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ));
    InMux I__1703 (
            .O(N__11222),
            .I(N__11219));
    LocalMux I__1702 (
            .O(N__11219),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ));
    InMux I__1701 (
            .O(N__11216),
            .I(N__11213));
    LocalMux I__1700 (
            .O(N__11213),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ));
    InMux I__1699 (
            .O(N__11210),
            .I(N__11207));
    LocalMux I__1698 (
            .O(N__11207),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ));
    InMux I__1697 (
            .O(N__11204),
            .I(N__11201));
    LocalMux I__1696 (
            .O(N__11201),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ));
    InMux I__1695 (
            .O(N__11198),
            .I(N__11195));
    LocalMux I__1694 (
            .O(N__11195),
            .I(N__11192));
    Odrv4 I__1693 (
            .O(N__11192),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ));
    InMux I__1692 (
            .O(N__11189),
            .I(N__11186));
    LocalMux I__1691 (
            .O(N__11186),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ));
    InMux I__1690 (
            .O(N__11183),
            .I(N__11180));
    LocalMux I__1689 (
            .O(N__11180),
            .I(N__11177));
    Odrv4 I__1688 (
            .O(N__11177),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ));
    InMux I__1687 (
            .O(N__11174),
            .I(N__11171));
    LocalMux I__1686 (
            .O(N__11171),
            .I(N__11168));
    Odrv4 I__1685 (
            .O(N__11168),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ));
    InMux I__1684 (
            .O(N__11165),
            .I(N__11162));
    LocalMux I__1683 (
            .O(N__11162),
            .I(N__11159));
    Odrv4 I__1682 (
            .O(N__11159),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ));
    InMux I__1681 (
            .O(N__11156),
            .I(N__11153));
    LocalMux I__1680 (
            .O(N__11153),
            .I(N__11150));
    Odrv4 I__1679 (
            .O(N__11150),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ));
    CEMux I__1678 (
            .O(N__11147),
            .I(N__11142));
    CEMux I__1677 (
            .O(N__11146),
            .I(N__11139));
    CEMux I__1676 (
            .O(N__11145),
            .I(N__11136));
    LocalMux I__1675 (
            .O(N__11142),
            .I(N__11133));
    LocalMux I__1674 (
            .O(N__11139),
            .I(N__11130));
    LocalMux I__1673 (
            .O(N__11136),
            .I(N__11127));
    Span4Mux_v I__1672 (
            .O(N__11133),
            .I(N__11120));
    Span4Mux_v I__1671 (
            .O(N__11130),
            .I(N__11120));
    Span4Mux_h I__1670 (
            .O(N__11127),
            .I(N__11120));
    Odrv4 I__1669 (
            .O(N__11120),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    InMux I__1668 (
            .O(N__11117),
            .I(N__11110));
    InMux I__1667 (
            .O(N__11116),
            .I(N__11110));
    InMux I__1666 (
            .O(N__11115),
            .I(N__11107));
    LocalMux I__1665 (
            .O(N__11110),
            .I(N__11104));
    LocalMux I__1664 (
            .O(N__11107),
            .I(N__11101));
    Span4Mux_v I__1663 (
            .O(N__11104),
            .I(N__11098));
    Odrv4 I__1662 (
            .O(N__11101),
            .I(\phase_controller_inst1.stoper_tr.time_passed11 ));
    Odrv4 I__1661 (
            .O(N__11098),
            .I(\phase_controller_inst1.stoper_tr.time_passed11 ));
    CascadeMux I__1660 (
            .O(N__11093),
            .I(N__11090));
    InMux I__1659 (
            .O(N__11090),
            .I(N__11087));
    LocalMux I__1658 (
            .O(N__11087),
            .I(N__11084));
    Odrv4 I__1657 (
            .O(N__11084),
            .I(\phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa ));
    InMux I__1656 (
            .O(N__11081),
            .I(N__11077));
    InMux I__1655 (
            .O(N__11080),
            .I(N__11072));
    LocalMux I__1654 (
            .O(N__11077),
            .I(N__11068));
    InMux I__1653 (
            .O(N__11076),
            .I(N__11063));
    InMux I__1652 (
            .O(N__11075),
            .I(N__11063));
    LocalMux I__1651 (
            .O(N__11072),
            .I(N__11060));
    InMux I__1650 (
            .O(N__11071),
            .I(N__11057));
    Span4Mux_h I__1649 (
            .O(N__11068),
            .I(N__11050));
    LocalMux I__1648 (
            .O(N__11063),
            .I(N__11050));
    Span4Mux_s3_h I__1647 (
            .O(N__11060),
            .I(N__11050));
    LocalMux I__1646 (
            .O(N__11057),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__1645 (
            .O(N__11050),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    InMux I__1644 (
            .O(N__11045),
            .I(N__11038));
    InMux I__1643 (
            .O(N__11044),
            .I(N__11033));
    InMux I__1642 (
            .O(N__11043),
            .I(N__11033));
    InMux I__1641 (
            .O(N__11042),
            .I(N__11028));
    InMux I__1640 (
            .O(N__11041),
            .I(N__11028));
    LocalMux I__1639 (
            .O(N__11038),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__1638 (
            .O(N__11033),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__1637 (
            .O(N__11028),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__1636 (
            .O(N__11021),
            .I(N__11018));
    InMux I__1635 (
            .O(N__11018),
            .I(N__11015));
    LocalMux I__1634 (
            .O(N__11015),
            .I(N__11012));
    Odrv4 I__1633 (
            .O(N__11012),
            .I(\phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ));
    InMux I__1632 (
            .O(N__11009),
            .I(N__11006));
    LocalMux I__1631 (
            .O(N__11006),
            .I(N__11001));
    InMux I__1630 (
            .O(N__11005),
            .I(N__10998));
    InMux I__1629 (
            .O(N__11004),
            .I(N__10995));
    Odrv4 I__1628 (
            .O(N__11001),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    LocalMux I__1627 (
            .O(N__10998),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    LocalMux I__1626 (
            .O(N__10995),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    InMux I__1625 (
            .O(N__10988),
            .I(N__10985));
    LocalMux I__1624 (
            .O(N__10985),
            .I(N__10982));
    Odrv4 I__1623 (
            .O(N__10982),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ));
    InMux I__1622 (
            .O(N__10979),
            .I(N__10976));
    LocalMux I__1621 (
            .O(N__10976),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ));
    InMux I__1620 (
            .O(N__10973),
            .I(N__10970));
    LocalMux I__1619 (
            .O(N__10970),
            .I(N__10967));
    Odrv4 I__1618 (
            .O(N__10967),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    InMux I__1617 (
            .O(N__10964),
            .I(N__10961));
    LocalMux I__1616 (
            .O(N__10961),
            .I(N__10958));
    Odrv4 I__1615 (
            .O(N__10958),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ));
    InMux I__1614 (
            .O(N__10955),
            .I(N__10952));
    LocalMux I__1613 (
            .O(N__10952),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ));
    InMux I__1612 (
            .O(N__10949),
            .I(N__10946));
    LocalMux I__1611 (
            .O(N__10946),
            .I(N__10943));
    Odrv4 I__1610 (
            .O(N__10943),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ));
    InMux I__1609 (
            .O(N__10940),
            .I(N__10937));
    LocalMux I__1608 (
            .O(N__10937),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    InMux I__1607 (
            .O(N__10934),
            .I(N__10931));
    LocalMux I__1606 (
            .O(N__10931),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ));
    InMux I__1605 (
            .O(N__10928),
            .I(N__10925));
    LocalMux I__1604 (
            .O(N__10925),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    InMux I__1603 (
            .O(N__10922),
            .I(N__10919));
    LocalMux I__1602 (
            .O(N__10919),
            .I(N__10916));
    Odrv4 I__1601 (
            .O(N__10916),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ));
    InMux I__1600 (
            .O(N__10913),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19 ));
    CascadeMux I__1599 (
            .O(N__10910),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_ ));
    CascadeMux I__1598 (
            .O(N__10907),
            .I(N__10904));
    InMux I__1597 (
            .O(N__10904),
            .I(N__10901));
    LocalMux I__1596 (
            .O(N__10901),
            .I(N__10898));
    Span4Mux_s3_h I__1595 (
            .O(N__10898),
            .I(N__10895));
    Odrv4 I__1594 (
            .O(N__10895),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ));
    CascadeMux I__1593 (
            .O(N__10892),
            .I(N__10876));
    InMux I__1592 (
            .O(N__10891),
            .I(N__10853));
    InMux I__1591 (
            .O(N__10890),
            .I(N__10853));
    InMux I__1590 (
            .O(N__10889),
            .I(N__10853));
    InMux I__1589 (
            .O(N__10888),
            .I(N__10853));
    InMux I__1588 (
            .O(N__10887),
            .I(N__10853));
    InMux I__1587 (
            .O(N__10886),
            .I(N__10853));
    InMux I__1586 (
            .O(N__10885),
            .I(N__10853));
    InMux I__1585 (
            .O(N__10884),
            .I(N__10853));
    InMux I__1584 (
            .O(N__10883),
            .I(N__10846));
    InMux I__1583 (
            .O(N__10882),
            .I(N__10846));
    InMux I__1582 (
            .O(N__10881),
            .I(N__10846));
    CascadeMux I__1581 (
            .O(N__10880),
            .I(N__10843));
    InMux I__1580 (
            .O(N__10879),
            .I(N__10825));
    InMux I__1579 (
            .O(N__10876),
            .I(N__10825));
    InMux I__1578 (
            .O(N__10875),
            .I(N__10825));
    InMux I__1577 (
            .O(N__10874),
            .I(N__10825));
    InMux I__1576 (
            .O(N__10873),
            .I(N__10825));
    InMux I__1575 (
            .O(N__10872),
            .I(N__10825));
    InMux I__1574 (
            .O(N__10871),
            .I(N__10825));
    InMux I__1573 (
            .O(N__10870),
            .I(N__10825));
    LocalMux I__1572 (
            .O(N__10853),
            .I(N__10822));
    LocalMux I__1571 (
            .O(N__10846),
            .I(N__10819));
    InMux I__1570 (
            .O(N__10843),
            .I(N__10811));
    InMux I__1569 (
            .O(N__10842),
            .I(N__10811));
    LocalMux I__1568 (
            .O(N__10825),
            .I(N__10806));
    Span4Mux_h I__1567 (
            .O(N__10822),
            .I(N__10806));
    Span4Mux_v I__1566 (
            .O(N__10819),
            .I(N__10803));
    InMux I__1565 (
            .O(N__10818),
            .I(N__10800));
    InMux I__1564 (
            .O(N__10817),
            .I(N__10797));
    InMux I__1563 (
            .O(N__10816),
            .I(N__10794));
    LocalMux I__1562 (
            .O(N__10811),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__1561 (
            .O(N__10806),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__1560 (
            .O(N__10803),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    LocalMux I__1559 (
            .O(N__10800),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    LocalMux I__1558 (
            .O(N__10797),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    LocalMux I__1557 (
            .O(N__10794),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    InMux I__1556 (
            .O(N__10781),
            .I(N__10746));
    InMux I__1555 (
            .O(N__10780),
            .I(N__10746));
    InMux I__1554 (
            .O(N__10779),
            .I(N__10746));
    InMux I__1553 (
            .O(N__10778),
            .I(N__10746));
    InMux I__1552 (
            .O(N__10777),
            .I(N__10746));
    InMux I__1551 (
            .O(N__10776),
            .I(N__10746));
    InMux I__1550 (
            .O(N__10775),
            .I(N__10746));
    InMux I__1549 (
            .O(N__10774),
            .I(N__10746));
    InMux I__1548 (
            .O(N__10773),
            .I(N__10729));
    InMux I__1547 (
            .O(N__10772),
            .I(N__10729));
    InMux I__1546 (
            .O(N__10771),
            .I(N__10729));
    InMux I__1545 (
            .O(N__10770),
            .I(N__10729));
    InMux I__1544 (
            .O(N__10769),
            .I(N__10729));
    InMux I__1543 (
            .O(N__10768),
            .I(N__10729));
    InMux I__1542 (
            .O(N__10767),
            .I(N__10729));
    InMux I__1541 (
            .O(N__10766),
            .I(N__10729));
    InMux I__1540 (
            .O(N__10765),
            .I(N__10722));
    InMux I__1539 (
            .O(N__10764),
            .I(N__10722));
    InMux I__1538 (
            .O(N__10763),
            .I(N__10722));
    LocalMux I__1537 (
            .O(N__10746),
            .I(N__10715));
    LocalMux I__1536 (
            .O(N__10729),
            .I(N__10715));
    LocalMux I__1535 (
            .O(N__10722),
            .I(N__10712));
    InMux I__1534 (
            .O(N__10721),
            .I(N__10704));
    InMux I__1533 (
            .O(N__10720),
            .I(N__10704));
    Span4Mux_v I__1532 (
            .O(N__10715),
            .I(N__10699));
    Span4Mux_v I__1531 (
            .O(N__10712),
            .I(N__10699));
    InMux I__1530 (
            .O(N__10711),
            .I(N__10696));
    InMux I__1529 (
            .O(N__10710),
            .I(N__10693));
    InMux I__1528 (
            .O(N__10709),
            .I(N__10690));
    LocalMux I__1527 (
            .O(N__10704),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__1526 (
            .O(N__10699),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    LocalMux I__1525 (
            .O(N__10696),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    LocalMux I__1524 (
            .O(N__10693),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    LocalMux I__1523 (
            .O(N__10690),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    InMux I__1522 (
            .O(N__10679),
            .I(N__10676));
    LocalMux I__1521 (
            .O(N__10676),
            .I(N__10673));
    Glb2LocalMux I__1520 (
            .O(N__10673),
            .I(N__10670));
    GlobalMux I__1519 (
            .O(N__10670),
            .I(clk_12mhz));
    IoInMux I__1518 (
            .O(N__10667),
            .I(N__10664));
    LocalMux I__1517 (
            .O(N__10664),
            .I(N__10661));
    Span4Mux_s0_v I__1516 (
            .O(N__10661),
            .I(N__10658));
    Span4Mux_h I__1515 (
            .O(N__10658),
            .I(N__10655));
    Odrv4 I__1514 (
            .O(N__10655),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__1513 (
            .O(N__10652),
            .I(N__10649));
    LocalMux I__1512 (
            .O(N__10649),
            .I(N__10646));
    Odrv4 I__1511 (
            .O(N__10646),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ));
    InMux I__1510 (
            .O(N__10643),
            .I(N__10640));
    LocalMux I__1509 (
            .O(N__10640),
            .I(N__10637));
    Odrv4 I__1508 (
            .O(N__10637),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ));
    InMux I__1507 (
            .O(N__10634),
            .I(N__10631));
    LocalMux I__1506 (
            .O(N__10631),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ));
    InMux I__1505 (
            .O(N__10628),
            .I(N__10625));
    LocalMux I__1504 (
            .O(N__10625),
            .I(N__10622));
    Odrv4 I__1503 (
            .O(N__10622),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ));
    InMux I__1502 (
            .O(N__10619),
            .I(N__10615));
    InMux I__1501 (
            .O(N__10618),
            .I(N__10612));
    LocalMux I__1500 (
            .O(N__10615),
            .I(N__10609));
    LocalMux I__1499 (
            .O(N__10612),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ));
    Odrv4 I__1498 (
            .O(N__10609),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ));
    CascadeMux I__1497 (
            .O(N__10604),
            .I(N__10601));
    InMux I__1496 (
            .O(N__10601),
            .I(N__10598));
    LocalMux I__1495 (
            .O(N__10598),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_13 ));
    InMux I__1494 (
            .O(N__10595),
            .I(N__10591));
    InMux I__1493 (
            .O(N__10594),
            .I(N__10588));
    LocalMux I__1492 (
            .O(N__10591),
            .I(N__10585));
    LocalMux I__1491 (
            .O(N__10588),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ));
    Odrv4 I__1490 (
            .O(N__10585),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ));
    CascadeMux I__1489 (
            .O(N__10580),
            .I(N__10577));
    InMux I__1488 (
            .O(N__10577),
            .I(N__10574));
    LocalMux I__1487 (
            .O(N__10574),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_14 ));
    InMux I__1486 (
            .O(N__10571),
            .I(N__10567));
    InMux I__1485 (
            .O(N__10570),
            .I(N__10564));
    LocalMux I__1484 (
            .O(N__10567),
            .I(N__10561));
    LocalMux I__1483 (
            .O(N__10564),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv12 I__1482 (
            .O(N__10561),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ));
    CascadeMux I__1481 (
            .O(N__10556),
            .I(N__10553));
    InMux I__1480 (
            .O(N__10553),
            .I(N__10550));
    LocalMux I__1479 (
            .O(N__10550),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_15 ));
    InMux I__1478 (
            .O(N__10547),
            .I(N__10543));
    InMux I__1477 (
            .O(N__10546),
            .I(N__10540));
    LocalMux I__1476 (
            .O(N__10543),
            .I(N__10537));
    LocalMux I__1475 (
            .O(N__10540),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv12 I__1474 (
            .O(N__10537),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ));
    CascadeMux I__1473 (
            .O(N__10532),
            .I(N__10529));
    InMux I__1472 (
            .O(N__10529),
            .I(N__10526));
    LocalMux I__1471 (
            .O(N__10526),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_16 ));
    InMux I__1470 (
            .O(N__10523),
            .I(N__10519));
    InMux I__1469 (
            .O(N__10522),
            .I(N__10516));
    LocalMux I__1468 (
            .O(N__10519),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ));
    LocalMux I__1467 (
            .O(N__10516),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ));
    CascadeMux I__1466 (
            .O(N__10511),
            .I(N__10508));
    InMux I__1465 (
            .O(N__10508),
            .I(N__10505));
    LocalMux I__1464 (
            .O(N__10505),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_17 ));
    InMux I__1463 (
            .O(N__10502),
            .I(N__10498));
    InMux I__1462 (
            .O(N__10501),
            .I(N__10495));
    LocalMux I__1461 (
            .O(N__10498),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__1460 (
            .O(N__10495),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ));
    CascadeMux I__1459 (
            .O(N__10490),
            .I(N__10487));
    InMux I__1458 (
            .O(N__10487),
            .I(N__10484));
    LocalMux I__1457 (
            .O(N__10484),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_18 ));
    InMux I__1456 (
            .O(N__10481),
            .I(N__10477));
    InMux I__1455 (
            .O(N__10480),
            .I(N__10474));
    LocalMux I__1454 (
            .O(N__10477),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__1453 (
            .O(N__10474),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ));
    CascadeMux I__1452 (
            .O(N__10469),
            .I(N__10466));
    InMux I__1451 (
            .O(N__10466),
            .I(N__10463));
    LocalMux I__1450 (
            .O(N__10463),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_19 ));
    InMux I__1449 (
            .O(N__10460),
            .I(N__10456));
    InMux I__1448 (
            .O(N__10459),
            .I(N__10453));
    LocalMux I__1447 (
            .O(N__10456),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__1446 (
            .O(N__10453),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ));
    CascadeMux I__1445 (
            .O(N__10448),
            .I(N__10445));
    InMux I__1444 (
            .O(N__10445),
            .I(N__10442));
    LocalMux I__1443 (
            .O(N__10442),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_5 ));
    InMux I__1442 (
            .O(N__10439),
            .I(N__10435));
    InMux I__1441 (
            .O(N__10438),
            .I(N__10432));
    LocalMux I__1440 (
            .O(N__10435),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__1439 (
            .O(N__10432),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ));
    CascadeMux I__1438 (
            .O(N__10427),
            .I(N__10424));
    InMux I__1437 (
            .O(N__10424),
            .I(N__10421));
    LocalMux I__1436 (
            .O(N__10421),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_6 ));
    InMux I__1435 (
            .O(N__10418),
            .I(N__10414));
    InMux I__1434 (
            .O(N__10417),
            .I(N__10411));
    LocalMux I__1433 (
            .O(N__10414),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__1432 (
            .O(N__10411),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ));
    CascadeMux I__1431 (
            .O(N__10406),
            .I(N__10403));
    InMux I__1430 (
            .O(N__10403),
            .I(N__10400));
    LocalMux I__1429 (
            .O(N__10400),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_7 ));
    InMux I__1428 (
            .O(N__10397),
            .I(N__10393));
    InMux I__1427 (
            .O(N__10396),
            .I(N__10390));
    LocalMux I__1426 (
            .O(N__10393),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__1425 (
            .O(N__10390),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ));
    CascadeMux I__1424 (
            .O(N__10385),
            .I(N__10382));
    InMux I__1423 (
            .O(N__10382),
            .I(N__10379));
    LocalMux I__1422 (
            .O(N__10379),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_8 ));
    InMux I__1421 (
            .O(N__10376),
            .I(N__10373));
    LocalMux I__1420 (
            .O(N__10373),
            .I(N__10369));
    InMux I__1419 (
            .O(N__10372),
            .I(N__10366));
    Odrv4 I__1418 (
            .O(N__10369),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__1417 (
            .O(N__10366),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ));
    CascadeMux I__1416 (
            .O(N__10361),
            .I(N__10358));
    InMux I__1415 (
            .O(N__10358),
            .I(N__10355));
    LocalMux I__1414 (
            .O(N__10355),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_9 ));
    InMux I__1413 (
            .O(N__10352),
            .I(N__10349));
    LocalMux I__1412 (
            .O(N__10349),
            .I(N__10345));
    InMux I__1411 (
            .O(N__10348),
            .I(N__10342));
    Odrv4 I__1410 (
            .O(N__10345),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__1409 (
            .O(N__10342),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ));
    CascadeMux I__1408 (
            .O(N__10337),
            .I(N__10334));
    InMux I__1407 (
            .O(N__10334),
            .I(N__10331));
    LocalMux I__1406 (
            .O(N__10331),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_10 ));
    InMux I__1405 (
            .O(N__10328),
            .I(N__10325));
    LocalMux I__1404 (
            .O(N__10325),
            .I(N__10321));
    InMux I__1403 (
            .O(N__10324),
            .I(N__10318));
    Odrv4 I__1402 (
            .O(N__10321),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__1401 (
            .O(N__10318),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ));
    CascadeMux I__1400 (
            .O(N__10313),
            .I(N__10310));
    InMux I__1399 (
            .O(N__10310),
            .I(N__10307));
    LocalMux I__1398 (
            .O(N__10307),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_11 ));
    InMux I__1397 (
            .O(N__10304),
            .I(N__10300));
    InMux I__1396 (
            .O(N__10303),
            .I(N__10297));
    LocalMux I__1395 (
            .O(N__10300),
            .I(N__10294));
    LocalMux I__1394 (
            .O(N__10297),
            .I(N__10291));
    Odrv4 I__1393 (
            .O(N__10294),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__1392 (
            .O(N__10291),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ));
    CascadeMux I__1391 (
            .O(N__10286),
            .I(N__10283));
    InMux I__1390 (
            .O(N__10283),
            .I(N__10280));
    LocalMux I__1389 (
            .O(N__10280),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_12 ));
    InMux I__1388 (
            .O(N__10277),
            .I(N__10274));
    LocalMux I__1387 (
            .O(N__10274),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13 ));
    CascadeMux I__1386 (
            .O(N__10271),
            .I(N__10268));
    InMux I__1385 (
            .O(N__10268),
            .I(N__10265));
    LocalMux I__1384 (
            .O(N__10265),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8 ));
    InMux I__1383 (
            .O(N__10262),
            .I(N__10259));
    LocalMux I__1382 (
            .O(N__10259),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5 ));
    CascadeMux I__1381 (
            .O(N__10256),
            .I(N__10253));
    InMux I__1380 (
            .O(N__10253),
            .I(N__10250));
    LocalMux I__1379 (
            .O(N__10250),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4 ));
    InMux I__1378 (
            .O(N__10247),
            .I(N__10244));
    LocalMux I__1377 (
            .O(N__10244),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2 ));
    InMux I__1376 (
            .O(N__10241),
            .I(N__10237));
    InMux I__1375 (
            .O(N__10240),
            .I(N__10233));
    LocalMux I__1374 (
            .O(N__10237),
            .I(N__10230));
    InMux I__1373 (
            .O(N__10236),
            .I(N__10227));
    LocalMux I__1372 (
            .O(N__10233),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__1371 (
            .O(N__10230),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__1370 (
            .O(N__10227),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ));
    CascadeMux I__1369 (
            .O(N__10220),
            .I(N__10217));
    InMux I__1368 (
            .O(N__10217),
            .I(N__10214));
    LocalMux I__1367 (
            .O(N__10214),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_1 ));
    InMux I__1366 (
            .O(N__10211),
            .I(N__10207));
    InMux I__1365 (
            .O(N__10210),
            .I(N__10204));
    LocalMux I__1364 (
            .O(N__10207),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__1363 (
            .O(N__10204),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__1362 (
            .O(N__10199),
            .I(N__10196));
    LocalMux I__1361 (
            .O(N__10196),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_2 ));
    InMux I__1360 (
            .O(N__10193),
            .I(N__10189));
    InMux I__1359 (
            .O(N__10192),
            .I(N__10186));
    LocalMux I__1358 (
            .O(N__10189),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__1357 (
            .O(N__10186),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ));
    CascadeMux I__1356 (
            .O(N__10181),
            .I(N__10178));
    InMux I__1355 (
            .O(N__10178),
            .I(N__10175));
    LocalMux I__1354 (
            .O(N__10175),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_3 ));
    InMux I__1353 (
            .O(N__10172),
            .I(N__10168));
    InMux I__1352 (
            .O(N__10171),
            .I(N__10165));
    LocalMux I__1351 (
            .O(N__10168),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__1350 (
            .O(N__10165),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ));
    CascadeMux I__1349 (
            .O(N__10160),
            .I(N__10157));
    InMux I__1348 (
            .O(N__10157),
            .I(N__10154));
    LocalMux I__1347 (
            .O(N__10154),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_4 ));
    InMux I__1346 (
            .O(N__10151),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ));
    CascadeMux I__1345 (
            .O(N__10148),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_ ));
    CascadeMux I__1344 (
            .O(N__10145),
            .I(N__10142));
    InMux I__1343 (
            .O(N__10142),
            .I(N__10139));
    LocalMux I__1342 (
            .O(N__10139),
            .I(N__10136));
    Span4Mux_s3_h I__1341 (
            .O(N__10136),
            .I(N__10133));
    Odrv4 I__1340 (
            .O(N__10133),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ));
    InMux I__1339 (
            .O(N__10130),
            .I(N__10126));
    InMux I__1338 (
            .O(N__10129),
            .I(N__10122));
    LocalMux I__1337 (
            .O(N__10126),
            .I(N__10119));
    InMux I__1336 (
            .O(N__10125),
            .I(N__10116));
    LocalMux I__1335 (
            .O(N__10122),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__1334 (
            .O(N__10119),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__1333 (
            .O(N__10116),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__1332 (
            .O(N__10109),
            .I(N__10106));
    LocalMux I__1331 (
            .O(N__10106),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0 ));
    InMux I__1330 (
            .O(N__10103),
            .I(N__10100));
    LocalMux I__1329 (
            .O(N__10100),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16 ));
    CascadeMux I__1328 (
            .O(N__10097),
            .I(N__10094));
    InMux I__1327 (
            .O(N__10094),
            .I(N__10091));
    LocalMux I__1326 (
            .O(N__10091),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15 ));
    InMux I__1325 (
            .O(N__10088),
            .I(N__10085));
    LocalMux I__1324 (
            .O(N__10085),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14 ));
    CascadeMux I__1323 (
            .O(N__10082),
            .I(N__10079));
    InMux I__1322 (
            .O(N__10079),
            .I(N__10076));
    LocalMux I__1321 (
            .O(N__10076),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6 ));
    InMux I__1320 (
            .O(N__10073),
            .I(N__10070));
    LocalMux I__1319 (
            .O(N__10070),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7 ));
    CascadeMux I__1318 (
            .O(N__10067),
            .I(N__10064));
    InMux I__1317 (
            .O(N__10064),
            .I(N__10061));
    LocalMux I__1316 (
            .O(N__10061),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3 ));
    InMux I__1315 (
            .O(N__10058),
            .I(N__10054));
    InMux I__1314 (
            .O(N__10057),
            .I(N__10051));
    LocalMux I__1313 (
            .O(N__10054),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    LocalMux I__1312 (
            .O(N__10051),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    CascadeMux I__1311 (
            .O(N__10046),
            .I(N__10043));
    InMux I__1310 (
            .O(N__10043),
            .I(N__10040));
    LocalMux I__1309 (
            .O(N__10040),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    InMux I__1308 (
            .O(N__10037),
            .I(N__10033));
    InMux I__1307 (
            .O(N__10036),
            .I(N__10030));
    LocalMux I__1306 (
            .O(N__10033),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    LocalMux I__1305 (
            .O(N__10030),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    CascadeMux I__1304 (
            .O(N__10025),
            .I(N__10022));
    InMux I__1303 (
            .O(N__10022),
            .I(N__10019));
    LocalMux I__1302 (
            .O(N__10019),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    InMux I__1301 (
            .O(N__10016),
            .I(N__10012));
    InMux I__1300 (
            .O(N__10015),
            .I(N__10009));
    LocalMux I__1299 (
            .O(N__10012),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    LocalMux I__1298 (
            .O(N__10009),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    CascadeMux I__1297 (
            .O(N__10004),
            .I(N__10001));
    InMux I__1296 (
            .O(N__10001),
            .I(N__9998));
    LocalMux I__1295 (
            .O(N__9998),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    InMux I__1294 (
            .O(N__9995),
            .I(N__9991));
    InMux I__1293 (
            .O(N__9994),
            .I(N__9988));
    LocalMux I__1292 (
            .O(N__9991),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    LocalMux I__1291 (
            .O(N__9988),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    CascadeMux I__1290 (
            .O(N__9983),
            .I(N__9980));
    InMux I__1289 (
            .O(N__9980),
            .I(N__9977));
    LocalMux I__1288 (
            .O(N__9977),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ));
    InMux I__1287 (
            .O(N__9974),
            .I(N__9971));
    LocalMux I__1286 (
            .O(N__9971),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    InMux I__1285 (
            .O(N__9968),
            .I(N__9964));
    InMux I__1284 (
            .O(N__9967),
            .I(N__9961));
    LocalMux I__1283 (
            .O(N__9964),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__1282 (
            .O(N__9961),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    CascadeMux I__1281 (
            .O(N__9956),
            .I(N__9953));
    InMux I__1280 (
            .O(N__9953),
            .I(N__9950));
    LocalMux I__1279 (
            .O(N__9950),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ));
    InMux I__1278 (
            .O(N__9947),
            .I(N__9944));
    LocalMux I__1277 (
            .O(N__9944),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    InMux I__1276 (
            .O(N__9941),
            .I(N__9937));
    InMux I__1275 (
            .O(N__9940),
            .I(N__9934));
    LocalMux I__1274 (
            .O(N__9937),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    LocalMux I__1273 (
            .O(N__9934),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    CascadeMux I__1272 (
            .O(N__9929),
            .I(N__9926));
    InMux I__1271 (
            .O(N__9926),
            .I(N__9923));
    LocalMux I__1270 (
            .O(N__9923),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ));
    InMux I__1269 (
            .O(N__9920),
            .I(N__9917));
    LocalMux I__1268 (
            .O(N__9917),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ));
    InMux I__1267 (
            .O(N__9914),
            .I(N__9910));
    InMux I__1266 (
            .O(N__9913),
            .I(N__9907));
    LocalMux I__1265 (
            .O(N__9910),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    LocalMux I__1264 (
            .O(N__9907),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    CascadeMux I__1263 (
            .O(N__9902),
            .I(N__9899));
    InMux I__1262 (
            .O(N__9899),
            .I(N__9896));
    LocalMux I__1261 (
            .O(N__9896),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ));
    InMux I__1260 (
            .O(N__9893),
            .I(N__9889));
    InMux I__1259 (
            .O(N__9892),
            .I(N__9886));
    LocalMux I__1258 (
            .O(N__9889),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__1257 (
            .O(N__9886),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    CascadeMux I__1256 (
            .O(N__9881),
            .I(N__9878));
    InMux I__1255 (
            .O(N__9878),
            .I(N__9875));
    LocalMux I__1254 (
            .O(N__9875),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    InMux I__1253 (
            .O(N__9872),
            .I(N__9868));
    InMux I__1252 (
            .O(N__9871),
            .I(N__9865));
    LocalMux I__1251 (
            .O(N__9868),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__1250 (
            .O(N__9865),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    CascadeMux I__1249 (
            .O(N__9860),
            .I(N__9857));
    InMux I__1248 (
            .O(N__9857),
            .I(N__9854));
    LocalMux I__1247 (
            .O(N__9854),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    InMux I__1246 (
            .O(N__9851),
            .I(N__9847));
    InMux I__1245 (
            .O(N__9850),
            .I(N__9844));
    LocalMux I__1244 (
            .O(N__9847),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__1243 (
            .O(N__9844),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    CascadeMux I__1242 (
            .O(N__9839),
            .I(N__9836));
    InMux I__1241 (
            .O(N__9836),
            .I(N__9833));
    LocalMux I__1240 (
            .O(N__9833),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    InMux I__1239 (
            .O(N__9830),
            .I(N__9826));
    InMux I__1238 (
            .O(N__9829),
            .I(N__9823));
    LocalMux I__1237 (
            .O(N__9826),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    LocalMux I__1236 (
            .O(N__9823),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    CascadeMux I__1235 (
            .O(N__9818),
            .I(N__9815));
    InMux I__1234 (
            .O(N__9815),
            .I(N__9812));
    LocalMux I__1233 (
            .O(N__9812),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    InMux I__1232 (
            .O(N__9809),
            .I(N__9805));
    InMux I__1231 (
            .O(N__9808),
            .I(N__9802));
    LocalMux I__1230 (
            .O(N__9805),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    LocalMux I__1229 (
            .O(N__9802),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    CascadeMux I__1228 (
            .O(N__9797),
            .I(N__9794));
    InMux I__1227 (
            .O(N__9794),
            .I(N__9791));
    LocalMux I__1226 (
            .O(N__9791),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    InMux I__1225 (
            .O(N__9788),
            .I(N__9784));
    InMux I__1224 (
            .O(N__9787),
            .I(N__9781));
    LocalMux I__1223 (
            .O(N__9784),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    LocalMux I__1222 (
            .O(N__9781),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    CascadeMux I__1221 (
            .O(N__9776),
            .I(N__9773));
    InMux I__1220 (
            .O(N__9773),
            .I(N__9770));
    LocalMux I__1219 (
            .O(N__9770),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    InMux I__1218 (
            .O(N__9767),
            .I(N__9763));
    InMux I__1217 (
            .O(N__9766),
            .I(N__9760));
    LocalMux I__1216 (
            .O(N__9763),
            .I(N__9757));
    LocalMux I__1215 (
            .O(N__9760),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv4 I__1214 (
            .O(N__9757),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    CascadeMux I__1213 (
            .O(N__9752),
            .I(N__9749));
    InMux I__1212 (
            .O(N__9749),
            .I(N__9746));
    LocalMux I__1211 (
            .O(N__9746),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    InMux I__1210 (
            .O(N__9743),
            .I(N__9739));
    InMux I__1209 (
            .O(N__9742),
            .I(N__9736));
    LocalMux I__1208 (
            .O(N__9739),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    LocalMux I__1207 (
            .O(N__9736),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    CascadeMux I__1206 (
            .O(N__9731),
            .I(N__9728));
    InMux I__1205 (
            .O(N__9728),
            .I(N__9725));
    LocalMux I__1204 (
            .O(N__9725),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    CascadeMux I__1203 (
            .O(N__9722),
            .I(N__9717));
    CascadeMux I__1202 (
            .O(N__9721),
            .I(N__9714));
    CascadeMux I__1201 (
            .O(N__9720),
            .I(N__9711));
    InMux I__1200 (
            .O(N__9717),
            .I(N__9688));
    InMux I__1199 (
            .O(N__9714),
            .I(N__9688));
    InMux I__1198 (
            .O(N__9711),
            .I(N__9688));
    InMux I__1197 (
            .O(N__9710),
            .I(N__9679));
    InMux I__1196 (
            .O(N__9709),
            .I(N__9679));
    InMux I__1195 (
            .O(N__9708),
            .I(N__9679));
    InMux I__1194 (
            .O(N__9707),
            .I(N__9679));
    InMux I__1193 (
            .O(N__9706),
            .I(N__9668));
    InMux I__1192 (
            .O(N__9705),
            .I(N__9668));
    InMux I__1191 (
            .O(N__9704),
            .I(N__9668));
    InMux I__1190 (
            .O(N__9703),
            .I(N__9668));
    InMux I__1189 (
            .O(N__9702),
            .I(N__9651));
    InMux I__1188 (
            .O(N__9701),
            .I(N__9651));
    InMux I__1187 (
            .O(N__9700),
            .I(N__9651));
    InMux I__1186 (
            .O(N__9699),
            .I(N__9651));
    InMux I__1185 (
            .O(N__9698),
            .I(N__9651));
    InMux I__1184 (
            .O(N__9697),
            .I(N__9651));
    InMux I__1183 (
            .O(N__9696),
            .I(N__9651));
    InMux I__1182 (
            .O(N__9695),
            .I(N__9651));
    LocalMux I__1181 (
            .O(N__9688),
            .I(N__9646));
    LocalMux I__1180 (
            .O(N__9679),
            .I(N__9646));
    InMux I__1179 (
            .O(N__9678),
            .I(N__9638));
    InMux I__1178 (
            .O(N__9677),
            .I(N__9638));
    LocalMux I__1177 (
            .O(N__9668),
            .I(N__9631));
    LocalMux I__1176 (
            .O(N__9651),
            .I(N__9631));
    Span4Mux_s3_h I__1175 (
            .O(N__9646),
            .I(N__9631));
    InMux I__1174 (
            .O(N__9645),
            .I(N__9626));
    InMux I__1173 (
            .O(N__9644),
            .I(N__9626));
    InMux I__1172 (
            .O(N__9643),
            .I(N__9623));
    LocalMux I__1171 (
            .O(N__9638),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__1170 (
            .O(N__9631),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    LocalMux I__1169 (
            .O(N__9626),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    LocalMux I__1168 (
            .O(N__9623),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    CascadeMux I__1167 (
            .O(N__9614),
            .I(N__9595));
    InMux I__1166 (
            .O(N__9613),
            .I(N__9575));
    InMux I__1165 (
            .O(N__9612),
            .I(N__9575));
    InMux I__1164 (
            .O(N__9611),
            .I(N__9575));
    InMux I__1163 (
            .O(N__9610),
            .I(N__9575));
    InMux I__1162 (
            .O(N__9609),
            .I(N__9575));
    InMux I__1161 (
            .O(N__9608),
            .I(N__9575));
    InMux I__1160 (
            .O(N__9607),
            .I(N__9575));
    InMux I__1159 (
            .O(N__9606),
            .I(N__9575));
    InMux I__1158 (
            .O(N__9605),
            .I(N__9560));
    InMux I__1157 (
            .O(N__9604),
            .I(N__9560));
    InMux I__1156 (
            .O(N__9603),
            .I(N__9560));
    InMux I__1155 (
            .O(N__9602),
            .I(N__9560));
    InMux I__1154 (
            .O(N__9601),
            .I(N__9560));
    InMux I__1153 (
            .O(N__9600),
            .I(N__9560));
    InMux I__1152 (
            .O(N__9599),
            .I(N__9560));
    CascadeMux I__1151 (
            .O(N__9598),
            .I(N__9557));
    InMux I__1150 (
            .O(N__9595),
            .I(N__9547));
    InMux I__1149 (
            .O(N__9594),
            .I(N__9547));
    InMux I__1148 (
            .O(N__9593),
            .I(N__9547));
    InMux I__1147 (
            .O(N__9592),
            .I(N__9547));
    LocalMux I__1146 (
            .O(N__9575),
            .I(N__9542));
    LocalMux I__1145 (
            .O(N__9560),
            .I(N__9542));
    InMux I__1144 (
            .O(N__9557),
            .I(N__9534));
    InMux I__1143 (
            .O(N__9556),
            .I(N__9534));
    LocalMux I__1142 (
            .O(N__9547),
            .I(N__9531));
    Span4Mux_v I__1141 (
            .O(N__9542),
            .I(N__9528));
    InMux I__1140 (
            .O(N__9541),
            .I(N__9523));
    InMux I__1139 (
            .O(N__9540),
            .I(N__9523));
    InMux I__1138 (
            .O(N__9539),
            .I(N__9520));
    LocalMux I__1137 (
            .O(N__9534),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__1136 (
            .O(N__9531),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__1135 (
            .O(N__9528),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    LocalMux I__1134 (
            .O(N__9523),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    LocalMux I__1133 (
            .O(N__9520),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    InMux I__1132 (
            .O(N__9509),
            .I(N__9494));
    InMux I__1131 (
            .O(N__9508),
            .I(N__9494));
    InMux I__1130 (
            .O(N__9507),
            .I(N__9494));
    InMux I__1129 (
            .O(N__9506),
            .I(N__9494));
    InMux I__1128 (
            .O(N__9505),
            .I(N__9476));
    InMux I__1127 (
            .O(N__9504),
            .I(N__9469));
    InMux I__1126 (
            .O(N__9503),
            .I(N__9469));
    LocalMux I__1125 (
            .O(N__9494),
            .I(N__9466));
    InMux I__1124 (
            .O(N__9493),
            .I(N__9449));
    InMux I__1123 (
            .O(N__9492),
            .I(N__9449));
    InMux I__1122 (
            .O(N__9491),
            .I(N__9449));
    InMux I__1121 (
            .O(N__9490),
            .I(N__9449));
    InMux I__1120 (
            .O(N__9489),
            .I(N__9449));
    InMux I__1119 (
            .O(N__9488),
            .I(N__9449));
    InMux I__1118 (
            .O(N__9487),
            .I(N__9449));
    InMux I__1117 (
            .O(N__9486),
            .I(N__9449));
    InMux I__1116 (
            .O(N__9485),
            .I(N__9434));
    InMux I__1115 (
            .O(N__9484),
            .I(N__9434));
    InMux I__1114 (
            .O(N__9483),
            .I(N__9434));
    InMux I__1113 (
            .O(N__9482),
            .I(N__9434));
    InMux I__1112 (
            .O(N__9481),
            .I(N__9434));
    InMux I__1111 (
            .O(N__9480),
            .I(N__9434));
    InMux I__1110 (
            .O(N__9479),
            .I(N__9434));
    LocalMux I__1109 (
            .O(N__9476),
            .I(N__9431));
    InMux I__1108 (
            .O(N__9475),
            .I(N__9426));
    InMux I__1107 (
            .O(N__9474),
            .I(N__9426));
    LocalMux I__1106 (
            .O(N__9469),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__1105 (
            .O(N__9466),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__1104 (
            .O(N__9449),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__1103 (
            .O(N__9434),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__1102 (
            .O(N__9431),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__1101 (
            .O(N__9426),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    CascadeMux I__1100 (
            .O(N__9413),
            .I(N__9403));
    CascadeMux I__1099 (
            .O(N__9412),
            .I(N__9400));
    CascadeMux I__1098 (
            .O(N__9411),
            .I(N__9397));
    CascadeMux I__1097 (
            .O(N__9410),
            .I(N__9394));
    CascadeMux I__1096 (
            .O(N__9409),
            .I(N__9387));
    CascadeMux I__1095 (
            .O(N__9408),
            .I(N__9384));
    CascadeMux I__1094 (
            .O(N__9407),
            .I(N__9381));
    CascadeMux I__1093 (
            .O(N__9406),
            .I(N__9378));
    InMux I__1092 (
            .O(N__9403),
            .I(N__9360));
    InMux I__1091 (
            .O(N__9400),
            .I(N__9360));
    InMux I__1090 (
            .O(N__9397),
            .I(N__9360));
    InMux I__1089 (
            .O(N__9394),
            .I(N__9360));
    InMux I__1088 (
            .O(N__9393),
            .I(N__9351));
    InMux I__1087 (
            .O(N__9392),
            .I(N__9351));
    InMux I__1086 (
            .O(N__9391),
            .I(N__9351));
    InMux I__1085 (
            .O(N__9390),
            .I(N__9351));
    InMux I__1084 (
            .O(N__9387),
            .I(N__9339));
    InMux I__1083 (
            .O(N__9384),
            .I(N__9339));
    InMux I__1082 (
            .O(N__9381),
            .I(N__9339));
    InMux I__1081 (
            .O(N__9378),
            .I(N__9339));
    InMux I__1080 (
            .O(N__9377),
            .I(N__9334));
    InMux I__1079 (
            .O(N__9376),
            .I(N__9334));
    InMux I__1078 (
            .O(N__9375),
            .I(N__9325));
    InMux I__1077 (
            .O(N__9374),
            .I(N__9325));
    InMux I__1076 (
            .O(N__9373),
            .I(N__9325));
    InMux I__1075 (
            .O(N__9372),
            .I(N__9325));
    InMux I__1074 (
            .O(N__9371),
            .I(N__9318));
    InMux I__1073 (
            .O(N__9370),
            .I(N__9318));
    InMux I__1072 (
            .O(N__9369),
            .I(N__9318));
    LocalMux I__1071 (
            .O(N__9360),
            .I(N__9313));
    LocalMux I__1070 (
            .O(N__9351),
            .I(N__9313));
    InMux I__1069 (
            .O(N__9350),
            .I(N__9310));
    InMux I__1068 (
            .O(N__9349),
            .I(N__9305));
    InMux I__1067 (
            .O(N__9348),
            .I(N__9305));
    LocalMux I__1066 (
            .O(N__9339),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__1065 (
            .O(N__9334),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__1064 (
            .O(N__9325),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__1063 (
            .O(N__9318),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__1062 (
            .O(N__9313),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__1061 (
            .O(N__9310),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__1060 (
            .O(N__9305),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    CascadeMux I__1059 (
            .O(N__9290),
            .I(N__9287));
    InMux I__1058 (
            .O(N__9287),
            .I(N__9284));
    LocalMux I__1057 (
            .O(N__9284),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    CascadeMux I__1056 (
            .O(N__9281),
            .I(N__9278));
    InMux I__1055 (
            .O(N__9278),
            .I(N__9274));
    InMux I__1054 (
            .O(N__9277),
            .I(N__9271));
    LocalMux I__1053 (
            .O(N__9274),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__1052 (
            .O(N__9271),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    CascadeMux I__1051 (
            .O(N__9266),
            .I(N__9263));
    InMux I__1050 (
            .O(N__9263),
            .I(N__9260));
    LocalMux I__1049 (
            .O(N__9260),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    InMux I__1048 (
            .O(N__9257),
            .I(N__9254));
    LocalMux I__1047 (
            .O(N__9254),
            .I(N__9250));
    InMux I__1046 (
            .O(N__9253),
            .I(N__9247));
    Odrv4 I__1045 (
            .O(N__9250),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__1044 (
            .O(N__9247),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    CascadeMux I__1043 (
            .O(N__9242),
            .I(N__9239));
    InMux I__1042 (
            .O(N__9239),
            .I(N__9236));
    LocalMux I__1041 (
            .O(N__9236),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    InMux I__1040 (
            .O(N__9233),
            .I(N__9229));
    InMux I__1039 (
            .O(N__9232),
            .I(N__9226));
    LocalMux I__1038 (
            .O(N__9229),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__1037 (
            .O(N__9226),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    CascadeMux I__1036 (
            .O(N__9221),
            .I(N__9218));
    InMux I__1035 (
            .O(N__9218),
            .I(N__9215));
    LocalMux I__1034 (
            .O(N__9215),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    InMux I__1033 (
            .O(N__9212),
            .I(N__9208));
    InMux I__1032 (
            .O(N__9211),
            .I(N__9205));
    LocalMux I__1031 (
            .O(N__9208),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    LocalMux I__1030 (
            .O(N__9205),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    CascadeMux I__1029 (
            .O(N__9200),
            .I(N__9197));
    InMux I__1028 (
            .O(N__9197),
            .I(N__9194));
    LocalMux I__1027 (
            .O(N__9194),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ));
    InMux I__1026 (
            .O(N__9191),
            .I(N__9187));
    InMux I__1025 (
            .O(N__9190),
            .I(N__9184));
    LocalMux I__1024 (
            .O(N__9187),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    LocalMux I__1023 (
            .O(N__9184),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    CascadeMux I__1022 (
            .O(N__9179),
            .I(N__9176));
    InMux I__1021 (
            .O(N__9176),
            .I(N__9173));
    LocalMux I__1020 (
            .O(N__9173),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ));
    InMux I__1019 (
            .O(N__9170),
            .I(N__9167));
    LocalMux I__1018 (
            .O(N__9167),
            .I(N__9164));
    Span4Mux_v I__1017 (
            .O(N__9164),
            .I(N__9161));
    Odrv4 I__1016 (
            .O(N__9161),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    InMux I__1015 (
            .O(N__9158),
            .I(N__9154));
    InMux I__1014 (
            .O(N__9157),
            .I(N__9151));
    LocalMux I__1013 (
            .O(N__9154),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__1012 (
            .O(N__9151),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    CascadeMux I__1011 (
            .O(N__9146),
            .I(N__9143));
    InMux I__1010 (
            .O(N__9143),
            .I(N__9140));
    LocalMux I__1009 (
            .O(N__9140),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ));
    InMux I__1008 (
            .O(N__9137),
            .I(N__9133));
    InMux I__1007 (
            .O(N__9136),
            .I(N__9130));
    LocalMux I__1006 (
            .O(N__9133),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__1005 (
            .O(N__9130),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    CascadeMux I__1004 (
            .O(N__9125),
            .I(N__9122));
    InMux I__1003 (
            .O(N__9122),
            .I(N__9119));
    LocalMux I__1002 (
            .O(N__9119),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ));
    InMux I__1001 (
            .O(N__9116),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ));
    CascadeMux I__1000 (
            .O(N__9113),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_ ));
    CascadeMux I__999 (
            .O(N__9110),
            .I(N__9107));
    InMux I__998 (
            .O(N__9107),
            .I(N__9104));
    LocalMux I__997 (
            .O(N__9104),
            .I(N__9101));
    Span4Mux_v I__996 (
            .O(N__9101),
            .I(N__9098));
    Odrv4 I__995 (
            .O(N__9098),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ));
    InMux I__994 (
            .O(N__9095),
            .I(N__9092));
    LocalMux I__993 (
            .O(N__9092),
            .I(N__9089));
    Odrv4 I__992 (
            .O(N__9089),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ));
    CascadeMux I__991 (
            .O(N__9086),
            .I(N__9083));
    InMux I__990 (
            .O(N__9083),
            .I(N__9079));
    InMux I__989 (
            .O(N__9082),
            .I(N__9076));
    LocalMux I__988 (
            .O(N__9079),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__987 (
            .O(N__9076),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    CascadeMux I__986 (
            .O(N__9071),
            .I(N__9068));
    InMux I__985 (
            .O(N__9068),
            .I(N__9065));
    LocalMux I__984 (
            .O(N__9065),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    InMux I__983 (
            .O(N__9062),
            .I(N__9058));
    InMux I__982 (
            .O(N__9061),
            .I(N__9055));
    LocalMux I__981 (
            .O(N__9058),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__980 (
            .O(N__9055),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    CascadeMux I__979 (
            .O(N__9050),
            .I(N__9047));
    InMux I__978 (
            .O(N__9047),
            .I(N__9044));
    LocalMux I__977 (
            .O(N__9044),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    InMux I__976 (
            .O(N__9041),
            .I(N__9037));
    InMux I__975 (
            .O(N__9040),
            .I(N__9034));
    LocalMux I__974 (
            .O(N__9037),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__973 (
            .O(N__9034),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    CascadeMux I__972 (
            .O(N__9029),
            .I(N__9026));
    InMux I__971 (
            .O(N__9026),
            .I(N__9023));
    LocalMux I__970 (
            .O(N__9023),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    InMux I__969 (
            .O(N__9020),
            .I(N__9016));
    InMux I__968 (
            .O(N__9019),
            .I(N__9013));
    LocalMux I__967 (
            .O(N__9016),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__966 (
            .O(N__9013),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    CascadeMux I__965 (
            .O(N__9008),
            .I(N__9005));
    InMux I__964 (
            .O(N__9005),
            .I(N__9002));
    LocalMux I__963 (
            .O(N__9002),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    InMux I__962 (
            .O(N__8999),
            .I(N__8995));
    InMux I__961 (
            .O(N__8998),
            .I(N__8992));
    LocalMux I__960 (
            .O(N__8995),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    LocalMux I__959 (
            .O(N__8992),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    CascadeMux I__958 (
            .O(N__8987),
            .I(N__8984));
    InMux I__957 (
            .O(N__8984),
            .I(N__8981));
    LocalMux I__956 (
            .O(N__8981),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    InMux I__955 (
            .O(N__8978),
            .I(N__8974));
    InMux I__954 (
            .O(N__8977),
            .I(N__8971));
    LocalMux I__953 (
            .O(N__8974),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    LocalMux I__952 (
            .O(N__8971),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    CascadeMux I__951 (
            .O(N__8966),
            .I(N__8963));
    InMux I__950 (
            .O(N__8963),
            .I(N__8960));
    LocalMux I__949 (
            .O(N__8960),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    InMux I__948 (
            .O(N__8957),
            .I(N__8953));
    InMux I__947 (
            .O(N__8956),
            .I(N__8950));
    LocalMux I__946 (
            .O(N__8953),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__945 (
            .O(N__8950),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    CascadeMux I__944 (
            .O(N__8945),
            .I(N__8942));
    InMux I__943 (
            .O(N__8942),
            .I(N__8939));
    LocalMux I__942 (
            .O(N__8939),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    InMux I__941 (
            .O(N__8936),
            .I(N__8932));
    InMux I__940 (
            .O(N__8935),
            .I(N__8929));
    LocalMux I__939 (
            .O(N__8932),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__938 (
            .O(N__8929),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    CascadeMux I__937 (
            .O(N__8924),
            .I(N__8921));
    InMux I__936 (
            .O(N__8921),
            .I(N__8918));
    LocalMux I__935 (
            .O(N__8918),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    InMux I__934 (
            .O(N__8915),
            .I(N__8911));
    InMux I__933 (
            .O(N__8914),
            .I(N__8907));
    LocalMux I__932 (
            .O(N__8911),
            .I(N__8904));
    InMux I__931 (
            .O(N__8910),
            .I(N__8901));
    LocalMux I__930 (
            .O(N__8907),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__929 (
            .O(N__8904),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__928 (
            .O(N__8901),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    CascadeMux I__927 (
            .O(N__8894),
            .I(N__8891));
    InMux I__926 (
            .O(N__8891),
            .I(N__8888));
    LocalMux I__925 (
            .O(N__8888),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    InMux I__924 (
            .O(N__8885),
            .I(N__8881));
    InMux I__923 (
            .O(N__8884),
            .I(N__8878));
    LocalMux I__922 (
            .O(N__8881),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__921 (
            .O(N__8878),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    CascadeMux I__920 (
            .O(N__8873),
            .I(N__8870));
    InMux I__919 (
            .O(N__8870),
            .I(N__8867));
    LocalMux I__918 (
            .O(N__8867),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    InMux I__917 (
            .O(N__8864),
            .I(N__8860));
    InMux I__916 (
            .O(N__8863),
            .I(N__8857));
    LocalMux I__915 (
            .O(N__8860),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__914 (
            .O(N__8857),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    CascadeMux I__913 (
            .O(N__8852),
            .I(N__8849));
    InMux I__912 (
            .O(N__8849),
            .I(N__8846));
    LocalMux I__911 (
            .O(N__8846),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    InMux I__910 (
            .O(N__8843),
            .I(N__8839));
    InMux I__909 (
            .O(N__8842),
            .I(N__8836));
    LocalMux I__908 (
            .O(N__8839),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__907 (
            .O(N__8836),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    CascadeMux I__906 (
            .O(N__8831),
            .I(N__8828));
    InMux I__905 (
            .O(N__8828),
            .I(N__8825));
    LocalMux I__904 (
            .O(N__8825),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    InMux I__903 (
            .O(N__8822),
            .I(N__8818));
    InMux I__902 (
            .O(N__8821),
            .I(N__8815));
    LocalMux I__901 (
            .O(N__8818),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__900 (
            .O(N__8815),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    CascadeMux I__899 (
            .O(N__8810),
            .I(N__8807));
    InMux I__898 (
            .O(N__8807),
            .I(N__8804));
    LocalMux I__897 (
            .O(N__8804),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    InMux I__896 (
            .O(N__8801),
            .I(N__8797));
    InMux I__895 (
            .O(N__8800),
            .I(N__8794));
    LocalMux I__894 (
            .O(N__8797),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__893 (
            .O(N__8794),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    CascadeMux I__892 (
            .O(N__8789),
            .I(N__8786));
    InMux I__891 (
            .O(N__8786),
            .I(N__8783));
    LocalMux I__890 (
            .O(N__8783),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    InMux I__889 (
            .O(N__8780),
            .I(N__8776));
    InMux I__888 (
            .O(N__8779),
            .I(N__8773));
    LocalMux I__887 (
            .O(N__8776),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__886 (
            .O(N__8773),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__885 (
            .O(N__8768),
            .I(N__8765));
    LocalMux I__884 (
            .O(N__8765),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ));
    CascadeMux I__883 (
            .O(N__8762),
            .I(N__8759));
    InMux I__882 (
            .O(N__8759),
            .I(N__8756));
    LocalMux I__881 (
            .O(N__8756),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    CascadeMux I__880 (
            .O(N__8753),
            .I(N__8750));
    InMux I__879 (
            .O(N__8750),
            .I(N__8747));
    LocalMux I__878 (
            .O(N__8747),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18 ));
    InMux I__877 (
            .O(N__8744),
            .I(N__8741));
    LocalMux I__876 (
            .O(N__8741),
            .I(N__8738));
    Odrv4 I__875 (
            .O(N__8738),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11 ));
    CascadeMux I__874 (
            .O(N__8735),
            .I(\phase_controller_slave.stoper_hc.time_passed11_cascade_ ));
    CascadeMux I__873 (
            .O(N__8732),
            .I(N__8729));
    InMux I__872 (
            .O(N__8729),
            .I(N__8726));
    LocalMux I__871 (
            .O(N__8726),
            .I(N__8723));
    Span4Mux_h I__870 (
            .O(N__8723),
            .I(N__8720));
    Odrv4 I__869 (
            .O(N__8720),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0 ));
    InMux I__868 (
            .O(N__8717),
            .I(N__8714));
    LocalMux I__867 (
            .O(N__8714),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0 ));
    InMux I__866 (
            .O(N__8711),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ));
    InMux I__865 (
            .O(N__8708),
            .I(bfn_2_25_0_));
    InMux I__864 (
            .O(N__8705),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ));
    InMux I__863 (
            .O(N__8702),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17 ));
    InMux I__862 (
            .O(N__8699),
            .I(N__8696));
    LocalMux I__861 (
            .O(N__8696),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17 ));
    InMux I__860 (
            .O(N__8693),
            .I(N__8690));
    LocalMux I__859 (
            .O(N__8690),
            .I(N__8687));
    Odrv4 I__858 (
            .O(N__8687),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12 ));
    InMux I__857 (
            .O(N__8684),
            .I(N__8681));
    LocalMux I__856 (
            .O(N__8681),
            .I(N__8678));
    Odrv4 I__855 (
            .O(N__8678),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9 ));
    InMux I__854 (
            .O(N__8675),
            .I(N__8672));
    LocalMux I__853 (
            .O(N__8672),
            .I(N__8669));
    Odrv4 I__852 (
            .O(N__8669),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10 ));
    InMux I__851 (
            .O(N__8666),
            .I(N__8663));
    LocalMux I__850 (
            .O(N__8663),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19 ));
    InMux I__849 (
            .O(N__8660),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ));
    InMux I__848 (
            .O(N__8657),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ));
    InMux I__847 (
            .O(N__8654),
            .I(bfn_2_24_0_));
    InMux I__846 (
            .O(N__8651),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ));
    InMux I__845 (
            .O(N__8648),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ));
    InMux I__844 (
            .O(N__8645),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ));
    InMux I__843 (
            .O(N__8642),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ));
    InMux I__842 (
            .O(N__8639),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ));
    InMux I__841 (
            .O(N__8636),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ));
    InMux I__840 (
            .O(N__8633),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ));
    InMux I__839 (
            .O(N__8630),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ));
    InMux I__838 (
            .O(N__8627),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ));
    InMux I__837 (
            .O(N__8624),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ));
    InMux I__836 (
            .O(N__8621),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ));
    InMux I__835 (
            .O(N__8618),
            .I(N__8615));
    LocalMux I__834 (
            .O(N__8615),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ));
    InMux I__833 (
            .O(N__8612),
            .I(N__8609));
    LocalMux I__832 (
            .O(N__8609),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ));
    InMux I__831 (
            .O(N__8606),
            .I(N__8603));
    LocalMux I__830 (
            .O(N__8603),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ));
    InMux I__829 (
            .O(N__8600),
            .I(N__8597));
    LocalMux I__828 (
            .O(N__8597),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ));
    InMux I__827 (
            .O(N__8594),
            .I(N__8591));
    LocalMux I__826 (
            .O(N__8591),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ));
    InMux I__825 (
            .O(N__8588),
            .I(N__8585));
    LocalMux I__824 (
            .O(N__8585),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ));
    InMux I__823 (
            .O(N__8582),
            .I(N__8579));
    LocalMux I__822 (
            .O(N__8579),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ));
    InMux I__821 (
            .O(N__8576),
            .I(N__8573));
    LocalMux I__820 (
            .O(N__8573),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ));
    InMux I__819 (
            .O(N__8570),
            .I(N__8567));
    LocalMux I__818 (
            .O(N__8567),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ));
    InMux I__817 (
            .O(N__8564),
            .I(N__8561));
    LocalMux I__816 (
            .O(N__8561),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ));
    InMux I__815 (
            .O(N__8558),
            .I(N__8555));
    LocalMux I__814 (
            .O(N__8555),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ));
    InMux I__813 (
            .O(N__8552),
            .I(N__8549));
    LocalMux I__812 (
            .O(N__8549),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ));
    InMux I__811 (
            .O(N__8546),
            .I(N__8543));
    LocalMux I__810 (
            .O(N__8543),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ));
    InMux I__809 (
            .O(N__8540),
            .I(N__8537));
    LocalMux I__808 (
            .O(N__8537),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ));
    InMux I__807 (
            .O(N__8534),
            .I(N__8531));
    LocalMux I__806 (
            .O(N__8531),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ));
    InMux I__805 (
            .O(N__8528),
            .I(N__8525));
    LocalMux I__804 (
            .O(N__8525),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ));
    InMux I__803 (
            .O(N__8522),
            .I(N__8519));
    LocalMux I__802 (
            .O(N__8519),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ));
    InMux I__801 (
            .O(N__8516),
            .I(N__8513));
    LocalMux I__800 (
            .O(N__8513),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ));
    InMux I__799 (
            .O(N__8510),
            .I(N__8507));
    LocalMux I__798 (
            .O(N__8507),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ));
    InMux I__797 (
            .O(N__8504),
            .I(N__8501));
    LocalMux I__796 (
            .O(N__8501),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ));
    CascadeMux I__795 (
            .O(N__8498),
            .I(N__8495));
    InMux I__794 (
            .O(N__8495),
            .I(N__8492));
    LocalMux I__793 (
            .O(N__8492),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ));
    InMux I__792 (
            .O(N__8489),
            .I(N__8486));
    LocalMux I__791 (
            .O(N__8486),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0 ));
    CascadeMux I__790 (
            .O(N__8483),
            .I(\phase_controller_inst1.stoper_tr.time_passed11_cascade_ ));
    CascadeMux I__789 (
            .O(N__8480),
            .I(N__8477));
    InMux I__788 (
            .O(N__8477),
            .I(N__8474));
    LocalMux I__787 (
            .O(N__8474),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ));
    CascadeMux I__786 (
            .O(N__8471),
            .I(\phase_controller_inst1.stoper_hc.time_passed11_cascade_ ));
    CascadeMux I__785 (
            .O(N__8468),
            .I(N__8465));
    InMux I__784 (
            .O(N__8465),
            .I(N__8462));
    LocalMux I__783 (
            .O(N__8462),
            .I(N__8459));
    Span4Mux_s2_h I__782 (
            .O(N__8459),
            .I(N__8456));
    Odrv4 I__781 (
            .O(N__8456),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ));
    InMux I__780 (
            .O(N__8453),
            .I(N__8450));
    LocalMux I__779 (
            .O(N__8450),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ));
    CascadeMux I__778 (
            .O(N__8447),
            .I(N__8444));
    InMux I__777 (
            .O(N__8444),
            .I(N__8441));
    LocalMux I__776 (
            .O(N__8441),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ));
    InMux I__775 (
            .O(N__8438),
            .I(N__8435));
    LocalMux I__774 (
            .O(N__8435),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ));
    CascadeMux I__773 (
            .O(N__8432),
            .I(N__8429));
    InMux I__772 (
            .O(N__8429),
            .I(N__8426));
    LocalMux I__771 (
            .O(N__8426),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ));
    InMux I__770 (
            .O(N__8423),
            .I(N__8420));
    LocalMux I__769 (
            .O(N__8420),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ));
    CascadeMux I__768 (
            .O(N__8417),
            .I(N__8414));
    InMux I__767 (
            .O(N__8414),
            .I(N__8411));
    LocalMux I__766 (
            .O(N__8411),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ));
    InMux I__765 (
            .O(N__8408),
            .I(N__8405));
    LocalMux I__764 (
            .O(N__8405),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ));
    CascadeMux I__763 (
            .O(N__8402),
            .I(N__8399));
    InMux I__762 (
            .O(N__8399),
            .I(N__8396));
    LocalMux I__761 (
            .O(N__8396),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ));
    InMux I__760 (
            .O(N__8393),
            .I(N__8390));
    LocalMux I__759 (
            .O(N__8390),
            .I(rgb_drv_RNOZ0));
    InMux I__758 (
            .O(N__8387),
            .I(N__8384));
    LocalMux I__757 (
            .O(N__8384),
            .I(N_39_i_i));
    InMux I__756 (
            .O(N__8381),
            .I(N__8378));
    LocalMux I__755 (
            .O(N__8378),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ));
    InMux I__754 (
            .O(N__8375),
            .I(N__8372));
    LocalMux I__753 (
            .O(N__8372),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ));
    InMux I__752 (
            .O(N__8369),
            .I(N__8366));
    LocalMux I__751 (
            .O(N__8366),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ));
    InMux I__750 (
            .O(N__8363),
            .I(N__8360));
    LocalMux I__749 (
            .O(N__8360),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ));
    InMux I__748 (
            .O(N__8357),
            .I(N__8354));
    LocalMux I__747 (
            .O(N__8354),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ));
    InMux I__746 (
            .O(N__8351),
            .I(N__8348));
    LocalMux I__745 (
            .O(N__8348),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ));
    InMux I__744 (
            .O(N__8345),
            .I(N__8342));
    LocalMux I__743 (
            .O(N__8342),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ));
    InMux I__742 (
            .O(N__8339),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ));
    InMux I__741 (
            .O(N__8336),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ));
    InMux I__740 (
            .O(N__8333),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ));
    InMux I__739 (
            .O(N__8330),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ));
    InMux I__738 (
            .O(N__8327),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ));
    InMux I__737 (
            .O(N__8324),
            .I(bfn_1_19_0_));
    InMux I__736 (
            .O(N__8321),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ));
    InMux I__735 (
            .O(N__8318),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ));
    InMux I__734 (
            .O(N__8315),
            .I(N__8312));
    LocalMux I__733 (
            .O(N__8312),
            .I(N__8309));
    Span12Mux_s3_v I__732 (
            .O(N__8309),
            .I(N__8306));
    Span12Mux_h I__731 (
            .O(N__8306),
            .I(N__8303));
    Span12Mux_h I__730 (
            .O(N__8303),
            .I(N__8297));
    InMux I__729 (
            .O(N__8302),
            .I(N__8294));
    InMux I__728 (
            .O(N__8301),
            .I(N__8291));
    InMux I__727 (
            .O(N__8300),
            .I(N__8288));
    Odrv12 I__726 (
            .O(N__8297),
            .I(CONSTANT_ONE_NET));
    LocalMux I__725 (
            .O(N__8294),
            .I(CONSTANT_ONE_NET));
    LocalMux I__724 (
            .O(N__8291),
            .I(CONSTANT_ONE_NET));
    LocalMux I__723 (
            .O(N__8288),
            .I(CONSTANT_ONE_NET));
    InMux I__722 (
            .O(N__8279),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ));
    InMux I__721 (
            .O(N__8276),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ));
    InMux I__720 (
            .O(N__8273),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ));
    InMux I__719 (
            .O(N__8270),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ));
    InMux I__718 (
            .O(N__8267),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ));
    InMux I__717 (
            .O(N__8264),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ));
    InMux I__716 (
            .O(N__8261),
            .I(bfn_1_18_0_));
    InMux I__715 (
            .O(N__8258),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ));
    InMux I__714 (
            .O(N__8255),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ));
    InMux I__713 (
            .O(N__8252),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ));
    InMux I__712 (
            .O(N__8249),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ));
    InMux I__711 (
            .O(N__8246),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ));
    InMux I__710 (
            .O(N__8243),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ));
    InMux I__709 (
            .O(N__8240),
            .I(bfn_1_16_0_));
    InMux I__708 (
            .O(N__8237),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ));
    InMux I__707 (
            .O(N__8234),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ));
    InMux I__706 (
            .O(N__8231),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ));
    InMux I__705 (
            .O(N__8228),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ));
    InMux I__704 (
            .O(N__8225),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ));
    InMux I__703 (
            .O(N__8222),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ));
    InMux I__702 (
            .O(N__8219),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ));
    InMux I__701 (
            .O(N__8216),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ));
    InMux I__700 (
            .O(N__8213),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ));
    InMux I__699 (
            .O(N__8210),
            .I(bfn_1_15_0_));
    InMux I__698 (
            .O(N__8207),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ));
    InMux I__697 (
            .O(N__8204),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ));
    InMux I__696 (
            .O(N__8201),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ));
    InMux I__695 (
            .O(N__8198),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ));
    defparam IN_MUX_bfv_8_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_17_0_));
    defparam IN_MUX_bfv_8_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_18_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_8_18_0_));
    defparam IN_MUX_bfv_8_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_19_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_8_19_0_));
    defparam IN_MUX_bfv_2_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_23_0_));
    defparam IN_MUX_bfv_2_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_24_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_2_24_0_));
    defparam IN_MUX_bfv_2_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_25_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_2_25_0_));
    defparam IN_MUX_bfv_1_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_17_0_));
    defparam IN_MUX_bfv_1_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_18_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_1_18_0_));
    defparam IN_MUX_bfv_1_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_19_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_1_19_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_1_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_16_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_1_16_0_));
    defparam IN_MUX_bfv_5_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_17_0_));
    defparam IN_MUX_bfv_5_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_18_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_5_18_0_));
    defparam IN_MUX_bfv_5_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_19_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_5_19_0_));
    defparam IN_MUX_bfv_3_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_25_0_));
    defparam IN_MUX_bfv_3_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_26_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_3_26_0_));
    defparam IN_MUX_bfv_3_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_27_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_3_27_0_));
    defparam IN_MUX_bfv_3_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_19_0_));
    defparam IN_MUX_bfv_3_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_20_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_3_20_0_));
    defparam IN_MUX_bfv_3_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_21_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_3_21_0_));
    defparam IN_MUX_bfv_3_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_15_0_));
    defparam IN_MUX_bfv_3_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_16_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_3_16_0_));
    defparam IN_MUX_bfv_3_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_17_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_3_17_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_9_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_16_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_9_16_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_8_15_0_));
    defparam IN_MUX_bfv_8_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_16_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_8_16_0_));
    defparam IN_MUX_bfv_10_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_21_0_));
    defparam IN_MUX_bfv_10_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_22_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_10_22_0_));
    defparam IN_MUX_bfv_10_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_23_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_10_23_0_));
    defparam IN_MUX_bfv_10_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_24_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_10_24_0_));
    defparam IN_MUX_bfv_9_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_21_0_));
    defparam IN_MUX_bfv_9_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_22_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_9_22_0_));
    defparam IN_MUX_bfv_9_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_23_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_9_23_0_));
    defparam IN_MUX_bfv_9_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_24_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_9_24_0_));
    ICE_GB \delay_measurement_inst.delay_tr_timer.running_RNICNBI_0  (
            .USERSIGNALTOGLOBALBUFFER(N__19934),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_tr_timer.N_255_i_g ));
    ICE_GB \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0  (
            .USERSIGNALTOGLOBALBUFFER(N__20702),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_hc_timer.N_253_i_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__8300),
            .CLKHFEN(N__8302),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__8301),
            .RGB2PWM(N__8387),
            .RGB1(rgb_g),
            .CURREN(N__8315),
            .RGB2(rgb_b),
            .RGB1PWM(N__8393),
            .RGB0PWM(N__20466),
            .RGB0(rgb_r));
    ICE_GB \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_0  (
            .USERSIGNALTOGLOBALBUFFER(N__20048),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_tr_timer.N_256_i_g ));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_1_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_1_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(N__8915),
            .in2(N__9110),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_14_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_1_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_1_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_1_14_1  (
            .in0(_gnd_net_),
            .in1(N__8885),
            .in2(_gnd_net_),
            .in3(N__8198),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_1_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_1_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(N__8864),
            .in2(N__8468),
            .in3(N__8228),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_1_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_1_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_1_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_1_14_3  (
            .in0(_gnd_net_),
            .in1(N__8843),
            .in2(_gnd_net_),
            .in3(N__8225),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_1_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_1_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(N__8822),
            .in2(_gnd_net_),
            .in3(N__8222),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_1_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_1_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_1_14_5  (
            .in0(_gnd_net_),
            .in1(N__8801),
            .in2(_gnd_net_),
            .in3(N__8219),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_1_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_1_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_1_14_6  (
            .in0(_gnd_net_),
            .in1(N__8780),
            .in2(_gnd_net_),
            .in3(N__8216),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_1_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_1_14_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9086),
            .in3(N__8213),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_1_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_1_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(N__9062),
            .in2(_gnd_net_),
            .in3(N__8210),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_1_15_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_1_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_1_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_1_15_1  (
            .in0(_gnd_net_),
            .in1(N__9041),
            .in2(_gnd_net_),
            .in3(N__8207),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_1_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_1_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_1_15_2  (
            .in0(_gnd_net_),
            .in1(N__9020),
            .in2(_gnd_net_),
            .in3(N__8204),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_1_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_1_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(N__8999),
            .in2(_gnd_net_),
            .in3(N__8201),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_1_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_1_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_1_15_4  (
            .in0(_gnd_net_),
            .in1(N__8978),
            .in2(_gnd_net_),
            .in3(N__8252),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_1_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_1_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_1_15_5  (
            .in0(_gnd_net_),
            .in1(N__8957),
            .in2(_gnd_net_),
            .in3(N__8249),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_1_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_1_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_1_15_6  (
            .in0(_gnd_net_),
            .in1(N__8936),
            .in2(_gnd_net_),
            .in3(N__8246),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_1_15_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_1_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_1_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_1_15_7  (
            .in0(_gnd_net_),
            .in1(N__9212),
            .in2(_gnd_net_),
            .in3(N__8243),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_1_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_1_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_1_16_0  (
            .in0(_gnd_net_),
            .in1(N__9191),
            .in2(_gnd_net_),
            .in3(N__8240),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_1_16_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_1_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_1_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_1_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_1_16_1  (
            .in0(_gnd_net_),
            .in1(N__9158),
            .in2(_gnd_net_),
            .in3(N__8237),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_1_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_1_16_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_1_16_2  (
            .in0(_gnd_net_),
            .in1(N__9137),
            .in2(_gnd_net_),
            .in3(N__8234),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_1_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_1_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_1_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_1_17_0  (
            .in0(_gnd_net_),
            .in1(N__10130),
            .in2(N__10145),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_17_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_1_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_1_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_1_17_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_1_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9281),
            .in3(N__8231),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_1_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_1_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_1_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_1_17_2  (
            .in0(_gnd_net_),
            .in1(N__9257),
            .in2(N__8480),
            .in3(N__8279),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_1_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_1_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_1_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_1_17_3  (
            .in0(_gnd_net_),
            .in1(N__9233),
            .in2(_gnd_net_),
            .in3(N__8276),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_1_17_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_1_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_1_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_1_17_4  (
            .in0(_gnd_net_),
            .in1(N__9893),
            .in2(_gnd_net_),
            .in3(N__8273),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_1_17_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_1_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_1_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_1_17_5  (
            .in0(_gnd_net_),
            .in1(N__9872),
            .in2(_gnd_net_),
            .in3(N__8270),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_1_17_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_1_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_1_17_6  (
            .in0(_gnd_net_),
            .in1(N__9851),
            .in2(_gnd_net_),
            .in3(N__8267),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_1_17_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_1_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_1_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_1_17_7  (
            .in0(_gnd_net_),
            .in1(N__9830),
            .in2(_gnd_net_),
            .in3(N__8264),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_1_18_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_1_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_1_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_1_18_0  (
            .in0(_gnd_net_),
            .in1(N__9809),
            .in2(_gnd_net_),
            .in3(N__8261),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ),
            .ltout(),
            .carryin(bfn_1_18_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_1_18_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_1_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_1_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_1_18_1  (
            .in0(_gnd_net_),
            .in1(N__9788),
            .in2(_gnd_net_),
            .in3(N__8258),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_1_18_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_1_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_1_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_1_18_2  (
            .in0(_gnd_net_),
            .in1(N__9766),
            .in2(_gnd_net_),
            .in3(N__8255),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_1_18_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_1_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_1_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_1_18_3  (
            .in0(_gnd_net_),
            .in1(N__9743),
            .in2(_gnd_net_),
            .in3(N__8339),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_1_18_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_1_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_1_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_1_18_4  (
            .in0(_gnd_net_),
            .in1(N__10058),
            .in2(_gnd_net_),
            .in3(N__8336),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_1_18_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_1_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_1_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_1_18_5  (
            .in0(_gnd_net_),
            .in1(N__10037),
            .in2(_gnd_net_),
            .in3(N__8333),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_1_18_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_1_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_1_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_1_18_6  (
            .in0(_gnd_net_),
            .in1(N__10016),
            .in2(_gnd_net_),
            .in3(N__8330),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_1_18_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_1_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_1_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_1_18_7  (
            .in0(_gnd_net_),
            .in1(N__9995),
            .in2(_gnd_net_),
            .in3(N__8327),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_1_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_1_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_1_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_1_19_0  (
            .in0(_gnd_net_),
            .in1(N__9968),
            .in2(_gnd_net_),
            .in3(N__8324),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ),
            .ltout(),
            .carryin(bfn_1_19_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_1_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_1_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_1_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_1_19_1  (
            .in0(_gnd_net_),
            .in1(N__9941),
            .in2(_gnd_net_),
            .in3(N__8321),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_1_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_1_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_1_19_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_1_19_2  (
            .in0(_gnd_net_),
            .in1(N__9914),
            .in2(_gnd_net_),
            .in3(N__8318),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_1_30_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_1_30_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_1_30_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_1_30_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_drv_RNO_LC_1_30_2.C_ON=1'b0;
    defparam rgb_drv_RNO_LC_1_30_2.SEQ_MODE=4'b0000;
    defparam rgb_drv_RNO_LC_1_30_2.LUT_INIT=16'b0101010100000000;
    LogicCell40 rgb_drv_RNO_LC_1_30_2 (
            .in0(N__20465),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13085),
            .lcout(rgb_drv_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_drv_RNO_0_LC_1_30_4.C_ON=1'b0;
    defparam rgb_drv_RNO_0_LC_1_30_4.SEQ_MODE=4'b0000;
    defparam rgb_drv_RNO_0_LC_1_30_4.LUT_INIT=16'b1010101001010101;
    LogicCell40 rgb_drv_RNO_0_LC_1_30_4 (
            .in0(N__20464),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13084),
            .lcout(N_39_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_2_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_2_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_2_14_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_2_14_0  (
            .in0(N__9601),
            .in1(N__11915),
            .in2(N__9722),
            .in3(N__8381),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20942),
            .ce(),
            .sr(N__20382));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_2_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_2_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_2_14_1 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_2_14_1  (
            .in0(N__9710),
            .in1(N__9605),
            .in2(N__11941),
            .in3(N__8375),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20942),
            .ce(),
            .sr(N__20382));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_2_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_2_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_2_14_3 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_2_14_3  (
            .in0(N__9708),
            .in1(N__9603),
            .in2(N__11939),
            .in3(N__8369),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20942),
            .ce(),
            .sr(N__20382));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_2_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_2_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_2_14_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_2_14_4  (
            .in0(N__9599),
            .in1(N__11913),
            .in2(N__9720),
            .in3(N__8363),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20942),
            .ce(),
            .sr(N__20382));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_2_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_2_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_2_14_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_2_14_5  (
            .in0(N__9707),
            .in1(N__9602),
            .in2(N__11938),
            .in3(N__8357),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20942),
            .ce(),
            .sr(N__20382));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_2_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_2_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_2_14_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_2_14_6  (
            .in0(N__9600),
            .in1(N__11914),
            .in2(N__9721),
            .in3(N__8351),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20942),
            .ce(),
            .sr(N__20382));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_2_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_2_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_2_14_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_2_14_7  (
            .in0(N__9709),
            .in1(N__9604),
            .in2(N__11940),
            .in3(N__8345),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20942),
            .ce(),
            .sr(N__20382));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_2_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_2_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_2_15_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_2_15_0  (
            .in0(N__9607),
            .in1(N__9700),
            .in2(N__11933),
            .in3(N__8453),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20940),
            .ce(),
            .sr(N__20390));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_2_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_2_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_2_15_1 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_2_15_1  (
            .in0(N__9695),
            .in1(N__11902),
            .in2(N__8447),
            .in3(N__9610),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20940),
            .ce(),
            .sr(N__20390));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_2_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_2_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_2_15_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_2_15_2  (
            .in0(N__9606),
            .in1(N__9699),
            .in2(N__11932),
            .in3(N__8438),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20940),
            .ce(),
            .sr(N__20390));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_2_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_2_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_2_15_3 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_2_15_3  (
            .in0(N__9696),
            .in1(N__11903),
            .in2(N__8432),
            .in3(N__9611),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20940),
            .ce(),
            .sr(N__20390));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_2_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_2_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_2_15_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_2_15_4  (
            .in0(N__9609),
            .in1(N__9702),
            .in2(N__11935),
            .in3(N__8423),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20940),
            .ce(),
            .sr(N__20390));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_2_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_2_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_2_15_5 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_2_15_5  (
            .in0(N__9697),
            .in1(N__11904),
            .in2(N__8417),
            .in3(N__9612),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20940),
            .ce(),
            .sr(N__20390));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_2_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_2_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_2_15_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_2_15_6  (
            .in0(N__9608),
            .in1(N__9701),
            .in2(N__11934),
            .in3(N__8408),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20940),
            .ce(),
            .sr(N__20390));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_2_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_2_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_2_15_7 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_2_15_7  (
            .in0(N__9698),
            .in1(N__11901),
            .in2(N__8402),
            .in3(N__9613),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20940),
            .ce(),
            .sr(N__20390));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_2_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_2_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_2_16_1 .LUT_INIT=16'b1010100010100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_2_16_1  (
            .in0(N__8489),
            .in1(N__9706),
            .in2(N__9614),
            .in3(N__11912),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20938),
            .ce(),
            .sr(N__20395));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_2_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_2_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_2_16_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_2_16_3  (
            .in0(N__9594),
            .in1(N__9705),
            .in2(N__11937),
            .in3(N__8510),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20938),
            .ce(),
            .sr(N__20395));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_2_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_2_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_2_16_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_2_16_5  (
            .in0(N__9593),
            .in1(N__9704),
            .in2(N__11936),
            .in3(N__8504),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20938),
            .ce(),
            .sr(N__20395));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_2_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_2_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_2_16_7 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_2_16_7  (
            .in0(N__9592),
            .in1(N__9703),
            .in2(N__8498),
            .in3(N__11911),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20938),
            .ce(),
            .sr(N__20395));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_2_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_2_17_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_2_17_1  (
            .in0(N__12169),
            .in1(N__9349),
            .in2(_gnd_net_),
            .in3(N__9475),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_2_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_2_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_2_17_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_2_17_2  (
            .in0(N__11042),
            .in1(N__8914),
            .in2(_gnd_net_),
            .in3(N__11005),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_2_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_2_17_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_2_17_3  (
            .in0(_gnd_net_),
            .in1(N__9348),
            .in2(_gnd_net_),
            .in3(N__9474),
            .lcout(\phase_controller_inst1.stoper_tr.time_passed11 ),
            .ltout(\phase_controller_inst1.stoper_tr.time_passed11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_2_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_2_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_2_17_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_2_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8483),
            .in3(N__11080),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_2_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_2_17_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_2_17_6  (
            .in0(_gnd_net_),
            .in1(N__9643),
            .in2(_gnd_net_),
            .in3(N__9539),
            .lcout(\phase_controller_inst1.stoper_hc.time_passed11 ),
            .ltout(\phase_controller_inst1.stoper_hc.time_passed11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_2_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_2_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_2_17_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_2_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8471),
            .in3(N__11041),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_2_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_2_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_2_18_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_2_18_1  (
            .in0(N__9485),
            .in1(N__12231),
            .in2(N__9413),
            .in3(N__8570),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20933),
            .ce(),
            .sr(N__20405));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_2_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_2_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_2_18_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_2_18_2  (
            .in0(N__9371),
            .in1(N__9484),
            .in2(N__12245),
            .in3(N__8564),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20933),
            .ce(),
            .sr(N__20405));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_2_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_2_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_2_18_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_2_18_3  (
            .in0(N__9482),
            .in1(N__12230),
            .in2(N__9412),
            .in3(N__8558),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20933),
            .ce(),
            .sr(N__20405));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_2_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_2_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_2_18_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_2_18_4  (
            .in0(N__9369),
            .in1(N__9479),
            .in2(N__12243),
            .in3(N__8552),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20933),
            .ce(),
            .sr(N__20405));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_2_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_2_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_2_18_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_2_18_5  (
            .in0(N__9480),
            .in1(N__12228),
            .in2(N__9410),
            .in3(N__8546),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20933),
            .ce(),
            .sr(N__20405));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_2_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_2_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_2_18_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_2_18_6  (
            .in0(N__9370),
            .in1(N__9483),
            .in2(N__12244),
            .in3(N__8540),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20933),
            .ce(),
            .sr(N__20405));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_2_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_2_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_2_18_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_2_18_7  (
            .in0(N__9481),
            .in1(N__12229),
            .in2(N__9411),
            .in3(N__8534),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20933),
            .ce(),
            .sr(N__20405));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_2_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_2_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_2_19_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_2_19_0  (
            .in0(N__9373),
            .in1(N__9488),
            .in2(N__12225),
            .in3(N__8528),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20927),
            .ce(),
            .sr(N__20410));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_2_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_2_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_2_19_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_2_19_1  (
            .in0(N__9487),
            .in1(N__12183),
            .in2(N__9406),
            .in3(N__8522),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20927),
            .ce(),
            .sr(N__20410));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_2_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_2_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_2_19_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_2_19_2  (
            .in0(N__9375),
            .in1(N__9492),
            .in2(N__12227),
            .in3(N__8516),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20927),
            .ce(),
            .sr(N__20410));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_2_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_2_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_2_19_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_2_19_3  (
            .in0(N__9491),
            .in1(N__12185),
            .in2(N__9408),
            .in3(N__8618),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20927),
            .ce(),
            .sr(N__20410));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_2_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_2_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_2_19_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_2_19_4  (
            .in0(N__9372),
            .in1(N__9486),
            .in2(N__12224),
            .in3(N__8612),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20927),
            .ce(),
            .sr(N__20410));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_2_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_2_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_2_19_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_2_19_5  (
            .in0(N__9493),
            .in1(N__12186),
            .in2(N__9409),
            .in3(N__8606),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20927),
            .ce(),
            .sr(N__20410));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_2_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_2_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_2_19_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_2_19_6  (
            .in0(N__9374),
            .in1(N__9490),
            .in2(N__12226),
            .in3(N__8600),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20927),
            .ce(),
            .sr(N__20410));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_2_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_2_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_2_19_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_2_19_7  (
            .in0(N__9489),
            .in1(N__12184),
            .in2(N__9407),
            .in3(N__8594),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20927),
            .ce(),
            .sr(N__20410));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_2_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_2_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_2_20_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_2_20_0  (
            .in0(N__9509),
            .in1(N__9393),
            .in2(N__12220),
            .in3(N__10109),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20923),
            .ce(),
            .sr(N__20413));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_2_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_2_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_2_20_1 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_2_20_1  (
            .in0(N__9392),
            .in1(N__9508),
            .in2(N__12223),
            .in3(N__8588),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20923),
            .ce(),
            .sr(N__20413));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_2_20_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_2_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_2_20_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_2_20_5  (
            .in0(N__9391),
            .in1(N__9507),
            .in2(N__12222),
            .in3(N__8582),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20923),
            .ce(),
            .sr(N__20413));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_2_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_2_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_2_20_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_2_20_7  (
            .in0(N__9390),
            .in1(N__9506),
            .in2(N__12221),
            .in3(N__8576),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20923),
            .ce(),
            .sr(N__20413));
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_2_21_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_2_21_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_2_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_18_LC_2_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16793),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20919),
            .ce(N__11262),
            .sr(N__20415));
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_2_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_2_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_2_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_17_LC_2_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16754),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20919),
            .ce(N__11262),
            .sr(N__20415));
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_2_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_2_21_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_2_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_19_LC_2_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18551),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20919),
            .ce(N__11262),
            .sr(N__20415));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_2_23_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_2_23_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_2_23_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_2_23_0  (
            .in0(_gnd_net_),
            .in1(N__10241),
            .in2(N__10907),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_23_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_2_23_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_2_23_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_2_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_2_23_1  (
            .in0(_gnd_net_),
            .in1(N__10211),
            .in2(_gnd_net_),
            .in3(N__8633),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_2_23_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_2_23_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_2_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_2_23_2  (
            .in0(_gnd_net_),
            .in1(N__10193),
            .in2(N__8732),
            .in3(N__8630),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_2_23_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_2_23_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_2_23_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_2_23_3  (
            .in0(_gnd_net_),
            .in1(N__10172),
            .in2(_gnd_net_),
            .in3(N__8627),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_2_23_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_2_23_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_2_23_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_2_23_4  (
            .in0(_gnd_net_),
            .in1(N__10460),
            .in2(_gnd_net_),
            .in3(N__8624),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_2_23_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_2_23_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_2_23_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_2_23_5  (
            .in0(_gnd_net_),
            .in1(N__10439),
            .in2(_gnd_net_),
            .in3(N__8621),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_2_23_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_2_23_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_2_23_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_2_23_6  (
            .in0(_gnd_net_),
            .in1(N__10418),
            .in2(_gnd_net_),
            .in3(N__8660),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_2_23_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_2_23_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_2_23_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_2_23_7  (
            .in0(_gnd_net_),
            .in1(N__10397),
            .in2(_gnd_net_),
            .in3(N__8657),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_2_24_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_2_24_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_2_24_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_2_24_0  (
            .in0(_gnd_net_),
            .in1(N__10376),
            .in2(_gnd_net_),
            .in3(N__8654),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9 ),
            .ltout(),
            .carryin(bfn_2_24_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_2_24_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_2_24_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_2_24_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_2_24_1  (
            .in0(_gnd_net_),
            .in1(N__10352),
            .in2(_gnd_net_),
            .in3(N__8651),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_2_24_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_2_24_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_2_24_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_2_24_2  (
            .in0(_gnd_net_),
            .in1(N__10328),
            .in2(_gnd_net_),
            .in3(N__8648),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_2_24_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_2_24_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_2_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_2_24_3  (
            .in0(_gnd_net_),
            .in1(N__10304),
            .in2(_gnd_net_),
            .in3(N__8645),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_2_24_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_2_24_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_2_24_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_2_24_4  (
            .in0(_gnd_net_),
            .in1(N__10618),
            .in2(_gnd_net_),
            .in3(N__8642),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_2_24_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_2_24_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_2_24_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_2_24_5  (
            .in0(_gnd_net_),
            .in1(N__10594),
            .in2(_gnd_net_),
            .in3(N__8639),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_2_24_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_2_24_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_2_24_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_2_24_6  (
            .in0(_gnd_net_),
            .in1(N__10570),
            .in2(_gnd_net_),
            .in3(N__8636),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_2_24_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_2_24_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_2_24_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_2_24_7  (
            .in0(_gnd_net_),
            .in1(N__10546),
            .in2(_gnd_net_),
            .in3(N__8711),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_2_25_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_2_25_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_2_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_2_25_0  (
            .in0(_gnd_net_),
            .in1(N__10523),
            .in2(_gnd_net_),
            .in3(N__8708),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17 ),
            .ltout(),
            .carryin(bfn_2_25_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_2_25_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_2_25_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_2_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_2_25_1  (
            .in0(_gnd_net_),
            .in1(N__10502),
            .in2(_gnd_net_),
            .in3(N__8705),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_2_25_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_2_25_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_2_25_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_2_25_2  (
            .in0(_gnd_net_),
            .in1(N__10481),
            .in2(_gnd_net_),
            .in3(N__8702),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_17_LC_2_26_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_17_LC_2_26_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_17_LC_2_26_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_17_LC_2_26_0  (
            .in0(N__10775),
            .in1(N__10874),
            .in2(N__12913),
            .in3(N__8699),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20894),
            .ce(),
            .sr(N__20424));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_12_LC_2_26_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_12_LC_2_26_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_12_LC_2_26_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_12_LC_2_26_1  (
            .in0(N__10871),
            .in1(N__10779),
            .in2(N__12910),
            .in3(N__8693),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20894),
            .ce(),
            .sr(N__20424));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_9_LC_2_26_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_9_LC_2_26_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_9_LC_2_26_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_9_LC_2_26_2  (
            .in0(N__10777),
            .in1(N__10875),
            .in2(N__12914),
            .in3(N__8684),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20894),
            .ce(),
            .sr(N__20424));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_1_LC_2_26_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_1_LC_2_26_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_1_LC_2_26_3 .LUT_INIT=16'b1010100010100010;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_1_LC_2_26_3  (
            .in0(N__8717),
            .in1(N__12892),
            .in2(N__10892),
            .in3(N__10781),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20894),
            .ce(),
            .sr(N__20424));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_10_LC_2_26_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_10_LC_2_26_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_10_LC_2_26_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_10_LC_2_26_4  (
            .in0(N__10774),
            .in1(N__10873),
            .in2(N__12912),
            .in3(N__8675),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20894),
            .ce(),
            .sr(N__20424));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_19_LC_2_26_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_19_LC_2_26_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_19_LC_2_26_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_19_LC_2_26_5  (
            .in0(N__10872),
            .in1(N__10780),
            .in2(N__12911),
            .in3(N__8666),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20894),
            .ce(),
            .sr(N__20424));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_18_LC_2_26_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_18_LC_2_26_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_18_LC_2_26_6 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_18_LC_2_26_6  (
            .in0(N__10776),
            .in1(N__12888),
            .in2(N__8753),
            .in3(N__10879),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20894),
            .ce(),
            .sr(N__20424));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_11_LC_2_26_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_11_LC_2_26_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_11_LC_2_26_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_11_LC_2_26_7  (
            .in0(N__10870),
            .in1(N__10778),
            .in2(N__12909),
            .in3(N__8744),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20894),
            .ce(),
            .sr(N__20424));
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_2_27_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_2_27_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_2_27_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_2_27_2  (
            .in0(_gnd_net_),
            .in1(N__10816),
            .in2(_gnd_net_),
            .in3(N__10709),
            .lcout(\phase_controller_slave.stoper_hc.time_passed11 ),
            .ltout(\phase_controller_slave.stoper_hc.time_passed11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_2_27_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_2_27_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_2_27_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_2_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8735),
            .in3(N__11962),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_2_27_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_2_27_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_2_27_4 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_2_27_4  (
            .in0(N__11963),
            .in1(N__11992),
            .in2(_gnd_net_),
            .in3(N__10240),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.stoper_state_0_LC_2_28_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_0_LC_2_28_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_0_LC_2_28_1 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_0_LC_2_28_1  (
            .in0(N__10720),
            .in1(N__10842),
            .in2(N__12904),
            .in3(N__11964),
            .lcout(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20880),
            .ce(N__20191),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.stoper_state_1_LC_2_28_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_1_LC_2_28_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_1_LC_2_28_6 .LUT_INIT=16'b0000110001010000;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_1_LC_2_28_6  (
            .in0(N__11965),
            .in1(N__12862),
            .in2(N__10880),
            .in3(N__10721),
            .lcout(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20880),
            .ce(N__20191),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_3_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_3_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_3_14_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_LC_3_14_0  (
            .in0(N__11442),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13883),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20941),
            .ce(N__11146),
            .sr(N__20376));
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_3_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_3_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_3_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_18_LC_3_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13934),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20941),
            .ce(N__11146),
            .sr(N__20376));
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_3_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_3_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_3_14_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_8_LC_3_14_6  (
            .in0(N__11443),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13847),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20941),
            .ce(N__11146),
            .sr(N__20376));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_3_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_3_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_3_15_0  (
            .in0(_gnd_net_),
            .in1(N__10643),
            .in2(N__8894),
            .in3(N__8910),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_3_15_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_3_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_3_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_3_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_3_15_1  (
            .in0(_gnd_net_),
            .in1(N__10652),
            .in2(N__8873),
            .in3(N__8884),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_3_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_3_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_3_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_3_15_2  (
            .in0(_gnd_net_),
            .in1(N__10988),
            .in2(N__8852),
            .in3(N__8863),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_3_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_3_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_3_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_3_15_3  (
            .in0(_gnd_net_),
            .in1(N__10634),
            .in2(N__8831),
            .in3(N__8842),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_3_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_3_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_3_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_3_15_4  (
            .in0(_gnd_net_),
            .in1(N__10964),
            .in2(N__8810),
            .in3(N__8821),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_3_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_3_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_3_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_3_15_5  (
            .in0(_gnd_net_),
            .in1(N__10628),
            .in2(N__8789),
            .in3(N__8800),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_3_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_3_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_3_15_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_3_15_6  (
            .in0(N__8779),
            .in1(N__8768),
            .in2(N__8762),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_3_15_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_3_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_3_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_3_15_7  (
            .in0(_gnd_net_),
            .in1(N__9095),
            .in2(N__9071),
            .in3(N__9082),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_3_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_3_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_3_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_3_16_0  (
            .in0(_gnd_net_),
            .in1(N__11156),
            .in2(N__9050),
            .in3(N__9061),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_3_16_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_3_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_3_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_3_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_3_16_1  (
            .in0(_gnd_net_),
            .in1(N__10922),
            .in2(N__9029),
            .in3(N__9040),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_3_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_3_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_3_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_3_16_2  (
            .in0(_gnd_net_),
            .in1(N__10934),
            .in2(N__9008),
            .in3(N__9019),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_3_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_3_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_3_16_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_3_16_3  (
            .in0(N__8998),
            .in1(N__10979),
            .in2(N__8987),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_3_16_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_3_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_3_16_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_3_16_4  (
            .in0(N__8977),
            .in1(N__10949),
            .in2(N__8966),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_3_16_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_3_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_3_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_3_16_5  (
            .in0(_gnd_net_),
            .in1(N__10955),
            .in2(N__8945),
            .in3(N__8956),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_3_16_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_3_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_3_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_3_16_6  (
            .in0(_gnd_net_),
            .in1(N__11165),
            .in2(N__8924),
            .in3(N__8935),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_3_16_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_3_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_3_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_3_16_7  (
            .in0(_gnd_net_),
            .in1(N__10973),
            .in2(N__9200),
            .in3(N__9211),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_3_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_3_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_3_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_3_17_0  (
            .in0(_gnd_net_),
            .in1(N__10940),
            .in2(N__9179),
            .in3(N__9190),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_3_17_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_3_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_3_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_3_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_3_17_1  (
            .in0(_gnd_net_),
            .in1(N__9170),
            .in2(N__9146),
            .in3(N__9157),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_3_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_3_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_3_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_3_17_2  (
            .in0(_gnd_net_),
            .in1(N__10928),
            .in2(N__9125),
            .in3(N__9136),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9116),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_3_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_3_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_3_17_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_3_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9113),
            .in3(N__11004),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_3_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_3_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_3_17_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_3_17_5  (
            .in0(N__9645),
            .in1(N__11882),
            .in2(_gnd_net_),
            .in3(N__9540),
            .lcout(\phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_3_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_3_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_3_17_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_3_17_6  (
            .in0(N__9350),
            .in1(N__12170),
            .in2(_gnd_net_),
            .in3(N__9505),
            .lcout(\phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_3_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_3_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_3_17_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_3_17_7  (
            .in0(N__9644),
            .in1(N__11881),
            .in2(_gnd_net_),
            .in3(N__9541),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_3_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_3_18_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_3_18_0 .LUT_INIT=16'b0000110001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_1_LC_3_18_0  (
            .in0(N__11044),
            .in1(N__11928),
            .in2(N__9598),
            .in3(N__9678),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20928),
            .ce(N__20195),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_3_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_3_18_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_3_18_1 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_0_LC_3_18_1  (
            .in0(N__9677),
            .in1(N__9556),
            .in2(N__11942),
            .in3(N__11043),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20928),
            .ce(N__20195),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_3_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_3_18_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_3_18_2 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_0_LC_3_18_2  (
            .in0(N__9376),
            .in1(N__9503),
            .in2(N__12241),
            .in3(N__11075),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20928),
            .ce(N__20195),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_3_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_3_18_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_3_18_6 .LUT_INIT=16'b0010000001100100;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_1_LC_3_18_6  (
            .in0(N__9377),
            .in1(N__9504),
            .in2(N__12242),
            .in3(N__11076),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20928),
            .ce(N__20195),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_3_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_3_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_3_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_3_19_0  (
            .in0(_gnd_net_),
            .in1(N__11216),
            .in2(N__9290),
            .in3(N__10125),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_3_19_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_3_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_3_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_3_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_3_19_1  (
            .in0(_gnd_net_),
            .in1(N__11210),
            .in2(N__9266),
            .in3(N__9277),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_3_19_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_3_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_3_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_3_19_2  (
            .in0(_gnd_net_),
            .in1(N__11237),
            .in2(N__9242),
            .in3(N__9253),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_3_19_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_3_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_3_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_3_19_3  (
            .in0(_gnd_net_),
            .in1(N__11228),
            .in2(N__9221),
            .in3(N__9232),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_3_19_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_3_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_3_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_3_19_4  (
            .in0(_gnd_net_),
            .in1(N__11204),
            .in2(N__9881),
            .in3(N__9892),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_3_19_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_3_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_3_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_3_19_5  (
            .in0(_gnd_net_),
            .in1(N__11222),
            .in2(N__9860),
            .in3(N__9871),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_3_19_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_3_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_3_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_3_19_6  (
            .in0(_gnd_net_),
            .in1(N__11174),
            .in2(N__9839),
            .in3(N__9850),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_3_19_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_3_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_3_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_3_19_7  (
            .in0(_gnd_net_),
            .in1(N__11198),
            .in2(N__9818),
            .in3(N__9829),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_3_20_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_3_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_3_20_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_3_20_0  (
            .in0(_gnd_net_),
            .in1(N__11297),
            .in2(N__9797),
            .in3(N__9808),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_3_20_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_3_20_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_3_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_3_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_3_20_1  (
            .in0(_gnd_net_),
            .in1(N__11279),
            .in2(N__9776),
            .in3(N__9787),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_3_20_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_3_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_3_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_3_20_2  (
            .in0(_gnd_net_),
            .in1(N__11303),
            .in2(N__9752),
            .in3(N__9767),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_3_20_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_3_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_3_20_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_3_20_3  (
            .in0(_gnd_net_),
            .in1(N__11309),
            .in2(N__9731),
            .in3(N__9742),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_3_20_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_3_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_3_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_3_20_4  (
            .in0(_gnd_net_),
            .in1(N__11183),
            .in2(N__10046),
            .in3(N__10057),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_3_20_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_3_20_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_3_20_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_3_20_5  (
            .in0(_gnd_net_),
            .in1(N__11288),
            .in2(N__10025),
            .in3(N__10036),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_3_20_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_3_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_3_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_3_20_6  (
            .in0(_gnd_net_),
            .in1(N__11189),
            .in2(N__10004),
            .in3(N__10015),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_3_20_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_3_20_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_3_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_3_20_7  (
            .in0(_gnd_net_),
            .in1(N__11318),
            .in2(N__9983),
            .in3(N__9994),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_3_21_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_3_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_3_21_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_3_21_0  (
            .in0(_gnd_net_),
            .in1(N__9974),
            .in2(N__9956),
            .in3(N__9967),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_3_21_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_3_21_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_3_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_3_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_3_21_1  (
            .in0(_gnd_net_),
            .in1(N__9947),
            .in2(N__9929),
            .in3(N__9940),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_3_21_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_3_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_3_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_3_21_2  (
            .in0(_gnd_net_),
            .in1(N__9920),
            .in2(N__9902),
            .in3(N__9913),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10151),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_3_21_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_3_21_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_3_21_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_3_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10148),
            .in3(N__11116),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_3_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_3_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_3_21_7 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_3_21_7  (
            .in0(N__11117),
            .in1(N__11071),
            .in2(_gnd_net_),
            .in3(N__10129),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_16_LC_3_23_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_16_LC_3_23_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_16_LC_3_23_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_16_LC_3_23_0  (
            .in0(N__10764),
            .in1(N__10883),
            .in2(N__12903),
            .in3(N__10103),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20902),
            .ce(),
            .sr(N__20416));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_15_LC_3_23_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_15_LC_3_23_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_15_LC_3_23_1 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_15_LC_3_23_1  (
            .in0(N__10881),
            .in1(N__12854),
            .in2(N__10097),
            .in3(N__10765),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20902),
            .ce(),
            .sr(N__20416));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_14_LC_3_23_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_14_LC_3_23_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_14_LC_3_23_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_14_LC_3_23_2  (
            .in0(N__10763),
            .in1(N__10882),
            .in2(N__12902),
            .in3(N__10088),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20902),
            .ce(),
            .sr(N__20416));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_6_LC_3_24_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_6_LC_3_24_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_6_LC_3_24_0 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_6_LC_3_24_0  (
            .in0(N__10886),
            .in1(N__12880),
            .in2(N__10082),
            .in3(N__10772),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20898),
            .ce(),
            .sr(N__20419));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_7_LC_3_24_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_7_LC_3_24_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_7_LC_3_24_1 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_7_LC_3_24_1  (
            .in0(N__10769),
            .in1(N__10891),
            .in2(N__12908),
            .in3(N__10073),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20898),
            .ce(),
            .sr(N__20419));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_3_LC_3_24_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_3_LC_3_24_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_3_LC_3_24_2 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_3_LC_3_24_2  (
            .in0(N__10884),
            .in1(N__12878),
            .in2(N__10067),
            .in3(N__10770),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20898),
            .ce(),
            .sr(N__20419));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_13_LC_3_24_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_13_LC_3_24_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_13_LC_3_24_3 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_13_LC_3_24_3  (
            .in0(N__10766),
            .in1(N__10888),
            .in2(N__12905),
            .in3(N__10277),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20898),
            .ce(),
            .sr(N__20419));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_8_LC_3_24_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_8_LC_3_24_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_8_LC_3_24_4 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_8_LC_3_24_4  (
            .in0(N__10887),
            .in1(N__12881),
            .in2(N__10271),
            .in3(N__10773),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20898),
            .ce(),
            .sr(N__20419));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_5_LC_3_24_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_5_LC_3_24_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_5_LC_3_24_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_5_LC_3_24_5  (
            .in0(N__10768),
            .in1(N__10890),
            .in2(N__12907),
            .in3(N__10262),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20898),
            .ce(),
            .sr(N__20419));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_4_LC_3_24_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_4_LC_3_24_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_4_LC_3_24_6 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_4_LC_3_24_6  (
            .in0(N__10885),
            .in1(N__12879),
            .in2(N__10256),
            .in3(N__10771),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20898),
            .ce(),
            .sr(N__20419));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_2_LC_3_24_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_2_LC_3_24_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_2_LC_3_24_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_2_LC_3_24_7  (
            .in0(N__10767),
            .in1(N__10889),
            .in2(N__12906),
            .in3(N__10247),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20898),
            .ce(),
            .sr(N__20419));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_3_25_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_3_25_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_3_25_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_3_25_0  (
            .in0(_gnd_net_),
            .in1(N__11582),
            .in2(N__10220),
            .in3(N__10236),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_3_25_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_3_25_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_3_25_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_3_25_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_3_25_1  (
            .in0(_gnd_net_),
            .in1(N__10199),
            .in2(N__11534),
            .in3(N__10210),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_3_25_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_3_25_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_3_25_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_3_25_2  (
            .in0(_gnd_net_),
            .in1(N__11450),
            .in2(N__10181),
            .in3(N__10192),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_3_25_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_3_25_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_3_25_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_3_25_3  (
            .in0(_gnd_net_),
            .in1(N__11525),
            .in2(N__10160),
            .in3(N__10171),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_3_25_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_3_25_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_3_25_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_3_25_4  (
            .in0(_gnd_net_),
            .in1(N__11594),
            .in2(N__10448),
            .in3(N__10459),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_3_25_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_3_25_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_3_25_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_3_25_5  (
            .in0(N__10438),
            .in1(N__11564),
            .in2(N__10427),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_3_25_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_3_25_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_3_25_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_3_25_6  (
            .in0(N__10417),
            .in1(N__11576),
            .in2(N__10406),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_3_25_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_3_25_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_3_25_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_3_25_7  (
            .in0(_gnd_net_),
            .in1(N__11369),
            .in2(N__10385),
            .in3(N__10396),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_3_26_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_3_26_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_3_26_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_3_26_0  (
            .in0(_gnd_net_),
            .in1(N__11726),
            .in2(N__10361),
            .in3(N__10372),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_3_26_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_3_26_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_3_26_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_3_26_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_3_26_1  (
            .in0(_gnd_net_),
            .in1(N__11765),
            .in2(N__10337),
            .in3(N__10348),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_3_26_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_3_26_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_3_26_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_3_26_2  (
            .in0(_gnd_net_),
            .in1(N__11663),
            .in2(N__10313),
            .in3(N__10324),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_3_26_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_3_26_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_3_26_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_3_26_3  (
            .in0(_gnd_net_),
            .in1(N__11759),
            .in2(N__10286),
            .in3(N__10303),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_3_26_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_3_26_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_3_26_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_3_26_4  (
            .in0(_gnd_net_),
            .in1(N__11771),
            .in2(N__10604),
            .in3(N__10619),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_3_26_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_3_26_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_3_26_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_3_26_5  (
            .in0(_gnd_net_),
            .in1(N__11618),
            .in2(N__10580),
            .in3(N__10595),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_3_26_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_3_26_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_3_26_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_3_26_6  (
            .in0(_gnd_net_),
            .in1(N__11360),
            .in2(N__10556),
            .in3(N__10571),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_3_26_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_3_26_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_3_26_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_3_26_7  (
            .in0(_gnd_net_),
            .in1(N__11612),
            .in2(N__10532),
            .in3(N__10547),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_3_27_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_3_27_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_3_27_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_3_27_0  (
            .in0(_gnd_net_),
            .in1(N__11600),
            .in2(N__10511),
            .in3(N__10522),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_3_27_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_3_27_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_3_27_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_3_27_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_3_27_1  (
            .in0(_gnd_net_),
            .in1(N__12050),
            .in2(N__10490),
            .in3(N__10501),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_3_27_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_3_27_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_3_27_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_3_27_2  (
            .in0(_gnd_net_),
            .in1(N__11606),
            .in2(N__10469),
            .in3(N__10480),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_27_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_27_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_27_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10913),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_3_27_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_3_27_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_3_27_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_3_27_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10910),
            .in3(N__11991),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_3_27_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_3_27_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_3_27_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_3_27_6  (
            .in0(N__10817),
            .in1(N__12853),
            .in2(_gnd_net_),
            .in3(N__10710),
            .lcout(\phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_3_28_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_3_28_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_3_28_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_3_28_6  (
            .in0(N__12861),
            .in1(N__10818),
            .in2(_gnd_net_),
            .in3(N__10711),
            .lcout(\phase_controller_slave.stoper_hc.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_3_30_2.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_3_30_2.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_3_30_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_3_30_2 (
            .in0(N__10679),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_4_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_4_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_4_15_0 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_2_LC_4_15_0  (
            .in0(N__11558),
            .in1(N__13343),
            .in2(N__11444),
            .in3(N__11515),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20936),
            .ce(N__11147),
            .sr(N__20377));
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_4_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_4_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_4_15_1 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_1_LC_4_15_1  (
            .in0(N__11514),
            .in1(N__11434),
            .in2(N__13652),
            .in3(N__11557),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20936),
            .ce(N__11147),
            .sr(N__20377));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_4_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_4_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_4_15_2 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_LC_4_15_2  (
            .in0(N__11439),
            .in1(N__11517),
            .in2(_gnd_net_),
            .in3(N__13703),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20936),
            .ce(N__11147),
            .sr(N__20377));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_4_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_4_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_4_15_3 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_LC_4_15_3  (
            .in0(N__11519),
            .in1(N__11441),
            .in2(_gnd_net_),
            .in3(N__14099),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20936),
            .ce(N__11147),
            .sr(N__20377));
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_4_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_4_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_4_15_4 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_3_LC_4_15_4  (
            .in0(N__11438),
            .in1(N__11516),
            .in2(N__13742),
            .in3(N__11468),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20936),
            .ce(N__11147),
            .sr(N__20377));
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_4_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_4_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_4_15_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_12_LC_4_15_5  (
            .in0(_gnd_net_),
            .in1(N__11712),
            .in2(_gnd_net_),
            .in3(N__13772),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20936),
            .ce(N__11147),
            .sr(N__20377));
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_4_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_4_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_4_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_16_LC_4_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14024),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20936),
            .ce(N__11147),
            .sr(N__20377));
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_4_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_4_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_4_15_7 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_5_LC_4_15_7  (
            .in0(N__11518),
            .in1(N__13382),
            .in2(_gnd_net_),
            .in3(N__11440),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20936),
            .ce(N__11147),
            .sr(N__20377));
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_4_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_4_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_4_16_0 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_14_LC_4_16_0  (
            .in0(N__13555),
            .in1(N__11650),
            .in2(_gnd_net_),
            .in3(N__13979),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20934),
            .ce(N__11145),
            .sr(N__20383));
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_4_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_4_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_4_16_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_13_LC_4_16_1  (
            .in0(N__11708),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15776),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20934),
            .ce(N__11145),
            .sr(N__20383));
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_4_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_4_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_4_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_17_LC_4_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14066),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20934),
            .ce(N__11145),
            .sr(N__20383));
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_4_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_4_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_4_16_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_11_LC_4_16_3  (
            .in0(N__11707),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13802),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20934),
            .ce(N__11145),
            .sr(N__20383));
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_4_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_4_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_4_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_19_LC_4_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13498),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20934),
            .ce(N__11145),
            .sr(N__20383));
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_4_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_4_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_4_16_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_10_LC_4_16_5  (
            .in0(N__11706),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13619),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20934),
            .ce(N__11145),
            .sr(N__20383));
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_4_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_4_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_4_16_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_15_LC_4_16_6  (
            .in0(N__13554),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11651),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20934),
            .ce(N__11145),
            .sr(N__20383));
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_4_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_4_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_4_16_7 .LUT_INIT=16'b1010111110101011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_9_LC_4_16_7  (
            .in0(N__13589),
            .in1(N__11750),
            .in2(N__11714),
            .in3(N__13556),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20934),
            .ce(N__11145),
            .sr(N__20383));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_4_LC_4_17_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_4_LC_4_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_4_LC_4_17_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_4_LC_4_17_0  (
            .in0(N__15468),
            .in1(N__15146),
            .in2(N__15342),
            .in3(N__14309),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20929),
            .ce(),
            .sr(N__20391));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_1_LC_4_17_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_1_LC_4_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_1_LC_4_17_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_1_LC_4_17_1  (
            .in0(N__15141),
            .in1(N__15316),
            .in2(N__15479),
            .in3(N__12617),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20929),
            .ce(),
            .sr(N__20391));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_4_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_4_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_4_17_2 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_4_17_2  (
            .in0(N__12378),
            .in1(N__11115),
            .in2(N__11093),
            .in3(N__11081),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20929),
            .ce(),
            .sr(N__20391));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_6_LC_4_17_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_6_LC_4_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_6_LC_4_17_3 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_6_LC_4_17_3  (
            .in0(N__15144),
            .in1(N__15319),
            .in2(N__14243),
            .in3(N__15471),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20929),
            .ce(),
            .sr(N__20391));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_2_LC_4_17_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_2_LC_4_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_2_LC_4_17_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_2_LC_4_17_4  (
            .in0(N__15467),
            .in1(N__15145),
            .in2(N__15341),
            .in3(N__14387),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20929),
            .ce(),
            .sr(N__20391));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_5_LC_4_17_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_5_LC_4_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_5_LC_4_17_5 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_5_LC_4_17_5  (
            .in0(N__15143),
            .in1(N__15318),
            .in2(N__14276),
            .in3(N__15470),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20929),
            .ce(),
            .sr(N__20391));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_4_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_4_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_4_17_6 .LUT_INIT=16'b1100110111000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_4_17_6  (
            .in0(N__11045),
            .in1(N__12314),
            .in2(N__11021),
            .in3(N__11009),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20929),
            .ce(),
            .sr(N__20391));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_3_LC_4_17_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_3_LC_4_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_3_LC_4_17_7 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_3_LC_4_17_7  (
            .in0(N__15142),
            .in1(N__15317),
            .in2(N__14342),
            .in3(N__15469),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20929),
            .ce(),
            .sr(N__20391));
    defparam \phase_controller_slave.stoper_tr.target_time_3_LC_4_18_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_3_LC_4_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_3_LC_4_18_0 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_3_LC_4_18_0  (
            .in0(N__14827),
            .in1(N__14717),
            .in2(N__16420),
            .in3(N__17099),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20924),
            .ce(N__12666),
            .sr(N__20396));
    defparam \phase_controller_slave.stoper_tr.target_time_9_LC_4_18_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_9_LC_4_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_9_LC_4_18_1 .LUT_INIT=16'b1111000011111101;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_9_LC_4_18_1  (
            .in0(N__16564),
            .in1(N__16997),
            .in2(N__16532),
            .in3(N__12737),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20924),
            .ce(N__12666),
            .sr(N__20396));
    defparam \phase_controller_slave.stoper_tr.target_time_8_LC_4_18_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_8_LC_4_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_8_LC_4_18_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_8_LC_4_18_2  (
            .in0(_gnd_net_),
            .in1(N__14720),
            .in2(_gnd_net_),
            .in3(N__18717),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20924),
            .ce(N__12666),
            .sr(N__20396));
    defparam \phase_controller_slave.stoper_tr.target_time_11_LC_4_18_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_11_LC_4_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_11_LC_4_18_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_11_LC_4_18_3  (
            .in0(_gnd_net_),
            .in1(N__12735),
            .in2(_gnd_net_),
            .in3(N__16645),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20924),
            .ce(N__12666),
            .sr(N__20396));
    defparam \phase_controller_slave.stoper_tr.target_time_2_LC_4_18_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_2_LC_4_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_2_LC_4_18_4 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_2_LC_4_18_4  (
            .in0(N__14826),
            .in1(N__14887),
            .in2(N__16460),
            .in3(N__14716),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20924),
            .ce(N__12666),
            .sr(N__20396));
    defparam \phase_controller_slave.stoper_tr.target_time_12_LC_4_18_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_12_LC_4_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_12_LC_4_18_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_12_LC_4_18_5  (
            .in0(_gnd_net_),
            .in1(N__12736),
            .in2(_gnd_net_),
            .in3(N__16672),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20924),
            .ce(N__12666),
            .sr(N__20396));
    defparam \phase_controller_slave.stoper_tr.target_time_6_LC_4_18_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_6_LC_4_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_6_LC_4_18_6 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_6_LC_4_18_6  (
            .in0(N__14828),
            .in1(N__14718),
            .in2(_gnd_net_),
            .in3(N__16819),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20924),
            .ce(N__12666),
            .sr(N__20396));
    defparam \phase_controller_slave.stoper_tr.target_time_7_LC_4_18_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_7_LC_4_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_7_LC_4_18_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_7_LC_4_18_7  (
            .in0(N__14719),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17851),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20924),
            .ce(N__12666),
            .sr(N__20396));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_4_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_4_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_4_19_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_LC_4_19_0  (
            .in0(N__14696),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17855),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20920),
            .ce(N__11269),
            .sr(N__20398));
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_4_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_4_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_4_19_1 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_3_LC_4_19_1  (
            .in0(N__14798),
            .in1(N__14692),
            .in2(N__16421),
            .in3(N__17092),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20920),
            .ce(N__11269),
            .sr(N__20398));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_4_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_4_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_4_19_2 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_LC_4_19_2  (
            .in0(N__14693),
            .in1(N__14799),
            .in2(_gnd_net_),
            .in3(N__17069),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20920),
            .ce(N__11269),
            .sr(N__20398));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_4_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_4_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_4_19_3 .LUT_INIT=16'b0000101000001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_LC_4_19_3  (
            .in0(N__16820),
            .in1(_gnd_net_),
            .in2(N__14815),
            .in3(N__14695),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20920),
            .ce(N__11269),
            .sr(N__20398));
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_4_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_4_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_4_19_4 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_1_LC_4_19_4  (
            .in0(N__14690),
            .in1(N__14794),
            .in2(N__16487),
            .in3(N__14879),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20920),
            .ce(N__11269),
            .sr(N__20398));
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_4_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_4_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_4_19_5 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_2_LC_4_19_5  (
            .in0(N__14880),
            .in1(N__16456),
            .in2(N__14814),
            .in3(N__14691),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20920),
            .ce(N__11269),
            .sr(N__20398));
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_4_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_4_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_4_19_6 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_5_LC_4_19_6  (
            .in0(N__14694),
            .in1(N__14800),
            .in2(_gnd_net_),
            .in3(N__16931),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20920),
            .ce(N__11269),
            .sr(N__20398));
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_4_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_4_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_4_19_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_8_LC_4_19_7  (
            .in0(N__18725),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14697),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20920),
            .ce(N__11269),
            .sr(N__20398));
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_4_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_4_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_4_20_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_15_LC_4_20_0  (
            .in0(N__14759),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17000),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20913),
            .ce(N__11273),
            .sr(N__20406));
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_4_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_4_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_4_20_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_13_LC_4_20_1  (
            .in0(_gnd_net_),
            .in1(N__12726),
            .in2(_gnd_net_),
            .in3(N__16622),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20913),
            .ce(N__11273),
            .sr(N__20406));
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_4_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_4_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_4_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_16_LC_4_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16715),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20913),
            .ce(N__11273),
            .sr(N__20406));
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_4_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_4_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_4_20_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_12_LC_4_20_3  (
            .in0(_gnd_net_),
            .in1(N__12725),
            .in2(_gnd_net_),
            .in3(N__16676),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20913),
            .ce(N__11273),
            .sr(N__20406));
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_4_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_4_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_4_20_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_11_LC_4_20_4  (
            .in0(N__12724),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16652),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20913),
            .ce(N__11273),
            .sr(N__20406));
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_4_20_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_4_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_4_20_5 .LUT_INIT=16'b1111111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_9_LC_4_20_5  (
            .in0(N__16998),
            .in1(N__12727),
            .in2(N__16565),
            .in3(N__16531),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20913),
            .ce(N__11273),
            .sr(N__20406));
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_4_20_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_4_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_4_20_6 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_14_LC_4_20_6  (
            .in0(N__14758),
            .in1(N__16999),
            .in2(_gnd_net_),
            .in3(N__17039),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20913),
            .ce(N__11273),
            .sr(N__20406));
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_4_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_4_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_4_20_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_10_LC_4_20_7  (
            .in0(_gnd_net_),
            .in1(N__12723),
            .in2(_gnd_net_),
            .in3(N__16592),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20913),
            .ce(N__11273),
            .sr(N__20406));
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_4_21_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_4_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_4_21_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_4_21_1  (
            .in0(N__15221),
            .in1(N__15466),
            .in2(_gnd_net_),
            .in3(N__15140),
            .lcout(\phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_4_3_LC_4_22_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_4_3_LC_4_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_4_3_LC_4_22_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_4_3_LC_4_22_0  (
            .in0(N__13973),
            .in1(N__13377),
            .in2(N__13553),
            .in3(N__13692),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_3_3_LC_4_22_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_3_3_LC_4_22_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_3_3_LC_4_22_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_3_3_LC_4_22_2  (
            .in0(N__13922),
            .in1(N__14061),
            .in2(N__13499),
            .in3(N__14019),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_3Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_3_LC_4_22_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_3_LC_4_22_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_3_LC_4_22_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a2_3_LC_4_22_3  (
            .in0(N__11354),
            .in1(N__11327),
            .in2(N__11348),
            .in3(N__11339),
            .lcout(\phase_controller_inst1.stoper_hc.N_144 ),
            .ltout(\phase_controller_inst1.stoper_hc.N_144_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a3_1_LC_4_22_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a3_1_LC_4_22_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a3_1_LC_4_22_4 .LUT_INIT=16'b0101000011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_f0_0_a3_1_LC_4_22_4  (
            .in0(N__13725),
            .in1(_gnd_net_),
            .in2(N__11345),
            .in3(N__13332),
            .lcout(\phase_controller_inst1.stoper_hc.N_122 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_0_6_LC_4_22_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_0_6_LC_4_22_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_0_6_LC_4_22_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_0_6_LC_4_22_5  (
            .in0(N__13761),
            .in1(N__13791),
            .in2(N__15771),
            .in3(N__13611),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_0Z0Z_6 ),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_9_LC_4_22_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_9_LC_4_22_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_9_LC_4_22_6 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_9_LC_4_22_6  (
            .in0(N__13584),
            .in1(_gnd_net_),
            .in2(N__11342),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2Z0Z_9 ),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2_6_LC_4_22_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2_6_LC_4_22_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2_6_LC_4_22_7 .LUT_INIT=16'b1011101010111011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2_6_LC_4_22_7  (
            .in0(N__11634),
            .in1(N__13540),
            .in2(N__11333),
            .in3(N__13974),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_i_o2_15_LC_4_23_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_i_o2_15_LC_4_23_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_i_o2_15_LC_4_23_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_i_o2_15_LC_4_23_1  (
            .in0(N__13926),
            .in1(N__14054),
            .in2(N__13490),
            .in3(N__14015),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_6_i_o2Z0Z_15 ),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_6_i_o2Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2_9_LC_4_23_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2_9_LC_4_23_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2_9_LC_4_23_2 .LUT_INIT=16'b1111000111110001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2_9_LC_4_23_2  (
            .in0(N__13541),
            .in1(N__13966),
            .in2(N__11330),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_o2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_1_6_LC_4_23_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_1_6_LC_4_23_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_1_6_LC_4_23_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_1_6_LC_4_23_6  (
            .in0(N__13881),
            .in1(N__13846),
            .in2(_gnd_net_),
            .in3(N__14088),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_1Z0Z_6 ),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a3_0_6_LC_4_23_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a3_0_6_LC_4_23_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a3_0_6_LC_4_23_7 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a3_0_6_LC_4_23_7  (
            .in0(N__11742),
            .in1(_gnd_net_),
            .in2(N__11321),
            .in3(N__13542),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_6_f1_0_i_i_a3_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.target_time_5_LC_4_24_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_5_LC_4_24_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_5_LC_4_24_0 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_5_LC_4_24_0  (
            .in0(N__11403),
            .in1(N__11493),
            .in2(_gnd_net_),
            .in3(N__13378),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20895),
            .ce(N__12044),
            .sr(N__20417));
    defparam \phase_controller_slave.stoper_hc.target_time_1_LC_4_24_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_1_LC_4_24_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_1_LC_4_24_1 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_1_LC_4_24_1  (
            .in0(N__11489),
            .in1(N__11397),
            .in2(N__13648),
            .in3(N__11555),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20895),
            .ce(N__12044),
            .sr(N__20417));
    defparam \phase_controller_slave.stoper_hc.target_time_7_LC_4_24_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_7_LC_4_24_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_7_LC_4_24_2 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_7_LC_4_24_2  (
            .in0(N__13882),
            .in1(_gnd_net_),
            .in2(N__11415),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20895),
            .ce(N__12044),
            .sr(N__20417));
    defparam \phase_controller_slave.stoper_hc.target_time_6_LC_4_24_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_6_LC_4_24_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_6_LC_4_24_3 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_6_LC_4_24_3  (
            .in0(N__11494),
            .in1(N__11404),
            .in2(_gnd_net_),
            .in3(N__14095),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20895),
            .ce(N__12044),
            .sr(N__20417));
    defparam \phase_controller_slave.stoper_hc.target_time_2_LC_4_24_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_2_LC_4_24_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_2_LC_4_24_4 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_2_LC_4_24_4  (
            .in0(N__11556),
            .in1(N__13339),
            .in2(N__11414),
            .in3(N__11490),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20895),
            .ce(N__12044),
            .sr(N__20417));
    defparam \phase_controller_slave.stoper_hc.target_time_4_LC_4_24_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_4_LC_4_24_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_4_LC_4_24_5 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_4_LC_4_24_5  (
            .in0(N__11492),
            .in1(N__13699),
            .in2(_gnd_net_),
            .in3(N__11402),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20895),
            .ce(N__12044),
            .sr(N__20417));
    defparam \phase_controller_slave.stoper_hc.target_time_3_LC_4_24_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_3_LC_4_24_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_3_LC_4_24_6 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_3_LC_4_24_6  (
            .in0(N__11401),
            .in1(N__11491),
            .in2(N__13741),
            .in3(N__11467),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20895),
            .ce(N__12044),
            .sr(N__20417));
    defparam \phase_controller_slave.stoper_hc.target_time_8_LC_4_24_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_8_LC_4_24_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_8_LC_4_24_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_8_LC_4_24_7  (
            .in0(_gnd_net_),
            .in1(N__11408),
            .in2(_gnd_net_),
            .in3(N__13842),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20895),
            .ce(N__12044),
            .sr(N__20417));
    defparam \phase_controller_slave.stoper_hc.target_time_15_LC_4_25_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_15_LC_4_25_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_15_LC_4_25_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_15_LC_4_25_0  (
            .in0(N__11644),
            .in1(N__13550),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20887),
            .ce(N__12042),
            .sr(N__20420));
    defparam \phase_controller_slave.stoper_hc.target_time_13_LC_4_25_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_13_LC_4_25_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_13_LC_4_25_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_13_LC_4_25_1  (
            .in0(N__11702),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15772),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20887),
            .ce(N__12042),
            .sr(N__20420));
    defparam \phase_controller_slave.stoper_hc.target_time_10_LC_4_25_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_10_LC_4_25_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_10_LC_4_25_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_10_LC_4_25_2  (
            .in0(_gnd_net_),
            .in1(N__11699),
            .in2(_gnd_net_),
            .in3(N__13618),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20887),
            .ce(N__12042),
            .sr(N__20420));
    defparam \phase_controller_slave.stoper_hc.target_time_12_LC_4_25_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_12_LC_4_25_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_12_LC_4_25_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_12_LC_4_25_4  (
            .in0(_gnd_net_),
            .in1(N__11701),
            .in2(_gnd_net_),
            .in3(N__13768),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20887),
            .ce(N__12042),
            .sr(N__20420));
    defparam \phase_controller_slave.stoper_hc.target_time_9_LC_4_25_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_9_LC_4_25_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_9_LC_4_25_5 .LUT_INIT=16'b1111111100001011;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_9_LC_4_25_5  (
            .in0(N__13552),
            .in1(N__11749),
            .in2(N__11713),
            .in3(N__13585),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20887),
            .ce(N__12042),
            .sr(N__20420));
    defparam \phase_controller_slave.stoper_hc.target_time_11_LC_4_25_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_11_LC_4_25_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_11_LC_4_25_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_11_LC_4_25_6  (
            .in0(_gnd_net_),
            .in1(N__11700),
            .in2(_gnd_net_),
            .in3(N__13798),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20887),
            .ce(N__12042),
            .sr(N__20420));
    defparam \phase_controller_slave.stoper_hc.target_time_14_LC_4_25_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_14_LC_4_25_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_14_LC_4_25_7 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_14_LC_4_25_7  (
            .in0(N__13551),
            .in1(N__11643),
            .in2(_gnd_net_),
            .in3(N__13975),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20887),
            .ce(N__12042),
            .sr(N__20420));
    defparam \phase_controller_slave.stoper_hc.target_time_16_LC_4_26_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_16_LC_4_26_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_16_LC_4_26_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_16_LC_4_26_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14020),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20881),
            .ce(N__12043),
            .sr(N__20422));
    defparam \phase_controller_slave.stoper_hc.target_time_19_LC_4_27_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_19_LC_4_27_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_19_LC_4_27_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_19_LC_4_27_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13491),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20875),
            .ce(N__12035),
            .sr(N__20423));
    defparam \phase_controller_slave.stoper_hc.target_time_17_LC_4_27_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_17_LC_4_27_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_17_LC_4_27_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_17_LC_4_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14062),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20875),
            .ce(N__12035),
            .sr(N__20423));
    defparam \phase_controller_slave.stoper_hc.target_time_18_LC_4_27_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_18_LC_4_27_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_18_LC_4_27_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_18_LC_4_27_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13933),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20875),
            .ce(N__12035),
            .sr(N__20423));
    defparam \phase_controller_slave.stoper_hc.time_passed_LC_4_28_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.time_passed_LC_4_28_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.time_passed_LC_4_28_7 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_slave.stoper_hc.time_passed_LC_4_28_7  (
            .in0(N__13281),
            .in1(N__11999),
            .in2(N__11975),
            .in3(N__11966),
            .lcout(\phase_controller_slave.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20870),
            .ce(),
            .sr(N__20425));
    defparam \phase_controller_inst1.state_2_LC_5_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_5_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_5_13_0 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_inst1.state_2_LC_5_13_0  (
            .in0(N__13217),
            .in1(N__12340),
            .in2(N__16890),
            .in3(N__12323),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20939),
            .ce(),
            .sr(N__20368));
    defparam \phase_controller_inst1.state_3_LC_5_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_5_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_5_13_2 .LUT_INIT=16'b1110111011111110;
    LogicCell40 \phase_controller_inst1.state_3_LC_5_13_2  (
            .in0(N__11786),
            .in1(N__12257),
            .in2(N__16891),
            .in3(N__13216),
            .lcout(\phase_controller_inst1.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20939),
            .ce(),
            .sr(N__20368));
    defparam \phase_controller_inst1.state_4_LC_5_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_5_13_3 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_5_13_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst1.state_4_LC_5_13_3  (
            .in0(N__13057),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12285),
            .lcout(\phase_controller_inst1.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20939),
            .ce(),
            .sr(N__20368));
    defparam \phase_controller_inst1.start_timer_hc_LC_5_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_5_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_5_13_7 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_5_13_7  (
            .in0(N__13193),
            .in1(N__12284),
            .in2(N__11888),
            .in3(N__11777),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20939),
            .ce(),
            .sr(N__20368));
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_5_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_5_14_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNI7NN7_0_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(N__12379),
            .in2(_gnd_net_),
            .in3(N__12358),
            .lcout(\phase_controller_inst1.N_107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_RNO_0_3_LC_5_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNO_0_3_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNO_0_3_LC_5_14_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.state_RNO_0_3_LC_5_14_3  (
            .in0(N__13058),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12277),
            .lcout(\phase_controller_inst1.N_110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_5_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_5_14_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_0_LC_5_14_5  (
            .in0(_gnd_net_),
            .in1(N__12339),
            .in2(_gnd_net_),
            .in3(N__12322),
            .lcout(\phase_controller_inst1.N_112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_0_LC_5_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_5_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_5_15_1 .LUT_INIT=16'b1111010001000100;
    LogicCell40 \phase_controller_inst1.state_0_LC_5_15_1  (
            .in0(N__12380),
            .in1(N__12359),
            .in2(N__19915),
            .in3(N__13160),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20935),
            .ce(),
            .sr(N__20373));
    defparam \phase_controller_inst1.T01_LC_5_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.T01_LC_5_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T01_LC_5_15_3 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \phase_controller_inst1.T01_LC_5_15_3  (
            .in0(N__12346),
            .in1(N__13138),
            .in2(N__13016),
            .in3(N__12286),
            .lcout(shift_flag_start),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20935),
            .ce(),
            .sr(N__20373));
    defparam \phase_controller_inst1.state_1_LC_5_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_5_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_5_15_5 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \phase_controller_inst1.state_1_LC_5_15_5  (
            .in0(N__12347),
            .in1(N__12321),
            .in2(N__19914),
            .in3(N__13159),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20935),
            .ce(),
            .sr(N__20373));
    defparam \phase_controller_inst1.start_timer_tr_LC_5_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_5_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_5_15_7 .LUT_INIT=16'b1100110011001110;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_5_15_7  (
            .in0(N__12127),
            .in1(N__13139),
            .in2(N__12290),
            .in3(N__12256),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20935),
            .ce(),
            .sr(N__20373));
    defparam \phase_controller_slave.stoper_tr.target_time_4_LC_5_16_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_4_LC_5_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_4_LC_5_16_5 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_4_LC_5_16_5  (
            .in0(N__14824),
            .in1(N__17068),
            .in2(_gnd_net_),
            .in3(N__14722),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20930),
            .ce(N__12671),
            .sr(N__20378));
    defparam \phase_controller_slave.stoper_tr.target_time_5_LC_5_16_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_5_LC_5_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_5_LC_5_16_6 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_5_LC_5_16_6  (
            .in0(N__14723),
            .in1(N__14825),
            .in2(_gnd_net_),
            .in3(N__16927),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20930),
            .ce(N__12671),
            .sr(N__20378));
    defparam \phase_controller_slave.stoper_tr.target_time_1_LC_5_16_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_1_LC_5_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_1_LC_5_16_7 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_1_LC_5_16_7  (
            .in0(N__14823),
            .in1(N__14721),
            .in2(N__16483),
            .in3(N__14888),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20930),
            .ce(N__12671),
            .sr(N__20378));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_5_17_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_5_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_5_17_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_5_17_0  (
            .in0(N__14433),
            .in1(N__12089),
            .in2(N__12080),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_5_17_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_5_17_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_5_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_5_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_5_17_1  (
            .in0(_gnd_net_),
            .in1(N__12071),
            .in2(N__12059),
            .in3(N__14398),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_5_17_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_5_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_5_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_5_17_2  (
            .in0(_gnd_net_),
            .in1(N__12497),
            .in2(N__12491),
            .in3(N__14368),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_5_17_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_5_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_5_17_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_5_17_3  (
            .in0(N__14320),
            .in1(N__12482),
            .in2(N__12476),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_5_17_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_5_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_5_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_5_17_4  (
            .in0(_gnd_net_),
            .in1(N__12467),
            .in2(N__12461),
            .in3(N__14287),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_5_17_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_5_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_5_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_5_17_5  (
            .in0(_gnd_net_),
            .in1(N__12452),
            .in2(N__12446),
            .in3(N__14254),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_5_17_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_5_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_5_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_5_17_6  (
            .in0(_gnd_net_),
            .in1(N__12437),
            .in2(N__12428),
            .in3(N__14225),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_5_17_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_5_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_5_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_5_17_7  (
            .in0(_gnd_net_),
            .in1(N__12419),
            .in2(N__12413),
            .in3(N__14651),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_5_18_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_5_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_5_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_5_18_0  (
            .in0(_gnd_net_),
            .in1(N__12404),
            .in2(N__12398),
            .in3(N__14621),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_5_18_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_5_18_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_5_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_5_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_5_18_1  (
            .in0(_gnd_net_),
            .in1(N__12599),
            .in2(N__12389),
            .in3(N__14597),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_5_18_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_5_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_5_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_5_18_2  (
            .in0(_gnd_net_),
            .in1(N__12584),
            .in2(N__12575),
            .in3(N__14570),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_5_18_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_5_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_5_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_5_18_3  (
            .in0(_gnd_net_),
            .in1(N__12566),
            .in2(N__12560),
            .in3(N__14546),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_5_18_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_5_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_5_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_5_18_4  (
            .in0(_gnd_net_),
            .in1(N__12695),
            .in2(N__12551),
            .in3(N__14516),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_5_18_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_5_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_5_18_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_5_18_5  (
            .in0(N__14492),
            .in1(N__12755),
            .in2(N__12542),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_5_18_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_5_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_5_18_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_5_18_6  (
            .in0(N__14465),
            .in1(N__12746),
            .in2(N__12533),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_5_18_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_5_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_5_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_5_18_7  (
            .in0(_gnd_net_),
            .in1(N__12608),
            .in2(N__12524),
            .in3(N__14987),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_5_19_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_5_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_5_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_5_19_0  (
            .in0(_gnd_net_),
            .in1(N__12677),
            .in2(N__12515),
            .in3(N__14960),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_5_19_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_5_19_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_5_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_5_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_5_19_1  (
            .in0(_gnd_net_),
            .in1(N__12686),
            .in2(N__12506),
            .in3(N__14936),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_5_19_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_5_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_5_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_5_19_2  (
            .in0(_gnd_net_),
            .in1(N__12590),
            .in2(N__12632),
            .in3(N__14912),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_5_19_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_5_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_5_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_5_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12623),
            .lcout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_5_19_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_5_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_5_19_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_5_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12620),
            .in3(N__14846),
            .lcout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_5_19_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_5_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_5_19_5 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_5_19_5  (
            .in0(N__14848),
            .in1(N__15168),
            .in2(_gnd_net_),
            .in3(N__14441),
            .lcout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_5_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_5_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_5_19_6 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_5_19_6  (
            .in0(N__14745),
            .in1(N__16994),
            .in2(_gnd_net_),
            .in3(N__17031),
            .lcout(\phase_controller_inst1.stoper_tr.N_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_5_19_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_5_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_5_19_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_5_19_7  (
            .in0(N__14847),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15167),
            .lcout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.target_time_16_LC_5_20_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_16_LC_5_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_16_LC_5_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_16_LC_5_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16711),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20907),
            .ce(N__12667),
            .sr(N__20399));
    defparam \phase_controller_slave.stoper_tr.target_time_10_LC_5_20_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_10_LC_5_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_10_LC_5_20_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_10_LC_5_20_1  (
            .in0(N__12721),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16588),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20907),
            .ce(N__12667),
            .sr(N__20399));
    defparam \phase_controller_slave.stoper_tr.target_time_19_LC_5_20_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_19_LC_5_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_19_LC_5_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_19_LC_5_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18547),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20907),
            .ce(N__12667),
            .sr(N__20399));
    defparam \phase_controller_slave.stoper_tr.target_time_14_LC_5_20_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_14_LC_5_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_14_LC_5_20_3 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_14_LC_5_20_3  (
            .in0(N__14756),
            .in1(N__16996),
            .in2(_gnd_net_),
            .in3(N__17038),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20907),
            .ce(N__12667),
            .sr(N__20399));
    defparam \phase_controller_slave.stoper_tr.target_time_15_LC_5_20_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_15_LC_5_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_15_LC_5_20_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_15_LC_5_20_4  (
            .in0(N__16995),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14757),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20907),
            .ce(N__12667),
            .sr(N__20399));
    defparam \phase_controller_slave.stoper_tr.target_time_13_LC_5_20_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_13_LC_5_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_13_LC_5_20_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_13_LC_5_20_5  (
            .in0(N__12722),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16618),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20907),
            .ce(N__12667),
            .sr(N__20399));
    defparam \phase_controller_slave.stoper_tr.target_time_18_LC_5_20_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_18_LC_5_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_18_LC_5_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_18_LC_5_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16792),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20907),
            .ce(N__12667),
            .sr(N__20399));
    defparam \phase_controller_slave.stoper_tr.target_time_17_LC_5_20_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_17_LC_5_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_17_LC_5_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_17_LC_5_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16750),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20907),
            .ce(N__12667),
            .sr(N__20399));
    defparam \phase_controller_slave.stoper_tr.time_passed_LC_5_21_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.time_passed_LC_5_21_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.time_passed_LC_5_21_2 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_slave.stoper_tr.time_passed_LC_5_21_2  (
            .in0(N__13126),
            .in1(N__14852),
            .in2(N__13445),
            .in3(N__15177),
            .lcout(\phase_controller_slave.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20903),
            .ce(),
            .sr(N__20407));
    defparam \phase_controller_slave.state_4_LC_5_22_3 .C_ON=1'b0;
    defparam \phase_controller_slave.state_4_LC_5_22_3 .SEQ_MODE=4'b1011;
    defparam \phase_controller_slave.state_4_LC_5_22_3 .LUT_INIT=16'b1010111011101110;
    LogicCell40 \phase_controller_slave.state_4_LC_5_22_3  (
            .in0(N__13094),
            .in1(N__12927),
            .in2(N__13083),
            .in3(N__13015),
            .lcout(\phase_controller_slave.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20899),
            .ce(),
            .sr(N__20411));
    defparam \phase_controller_slave.start_timer_tr_LC_5_22_4 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_tr_LC_5_22_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.start_timer_tr_LC_5_22_4 .LUT_INIT=16'b1010101010101110;
    LogicCell40 \phase_controller_slave.start_timer_tr_LC_5_22_4  (
            .in0(N__12638),
            .in1(N__15235),
            .in2(N__12936),
            .in3(N__13093),
            .lcout(\phase_controller_slave.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20899),
            .ce(),
            .sr(N__20411));
    defparam \phase_controller_slave.state_0_LC_5_22_7 .C_ON=1'b0;
    defparam \phase_controller_slave.state_0_LC_5_22_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_0_LC_5_22_7 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \phase_controller_slave.state_0_LC_5_22_7  (
            .in0(N__13417),
            .in1(N__13125),
            .in2(N__15707),
            .in3(N__13106),
            .lcout(\phase_controller_slave.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20899),
            .ce(),
            .sr(N__20411));
    defparam \phase_controller_slave.start_timer_tr_RNO_0_LC_5_23_3 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_tr_RNO_0_LC_5_23_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.start_timer_tr_RNO_0_LC_5_23_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.start_timer_tr_RNO_0_LC_5_23_3  (
            .in0(_gnd_net_),
            .in1(N__15699),
            .in2(_gnd_net_),
            .in3(N__13416),
            .lcout(\phase_controller_slave.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.state_RNIVDE2_0_LC_5_23_5 .C_ON=1'b0;
    defparam \phase_controller_slave.state_RNIVDE2_0_LC_5_23_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.state_RNIVDE2_0_LC_5_23_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.state_RNIVDE2_0_LC_5_23_5  (
            .in0(_gnd_net_),
            .in1(N__13127),
            .in2(_gnd_net_),
            .in3(N__13105),
            .lcout(\phase_controller_slave.state_RNIVDE2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.state_RNO_0_3_LC_5_24_1 .C_ON=1'b0;
    defparam \phase_controller_slave.state_RNO_0_3_LC_5_24_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.state_RNO_0_3_LC_5_24_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.state_RNO_0_3_LC_5_24_1  (
            .in0(N__13071),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13014),
            .lcout(\phase_controller_slave.state_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D2_LC_5_24_3.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_5_24_3.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_5_24_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D2_LC_5_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12977),
            .lcout(il_max_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20888),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.start_timer_hc_RNO_1_LC_5_24_4 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_hc_RNO_1_LC_5_24_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.start_timer_hc_RNO_1_LC_5_24_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.start_timer_hc_RNO_1_LC_5_24_4  (
            .in0(_gnd_net_),
            .in1(N__17264),
            .in2(_gnd_net_),
            .in3(N__12960),
            .lcout(\phase_controller_slave.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_24_5.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_24_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_24_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D1_LC_5_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12992),
            .lcout(il_max_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20888),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.state_1_LC_5_25_0 .C_ON=1'b0;
    defparam \phase_controller_slave.state_1_LC_5_25_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_1_LC_5_25_0 .LUT_INIT=16'b1010111000001100;
    LogicCell40 \phase_controller_slave.state_1_LC_5_25_0  (
            .in0(N__13288),
            .in1(N__15695),
            .in2(N__13421),
            .in3(N__13306),
            .lcout(\phase_controller_slave.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20882),
            .ce(),
            .sr(N__20418));
    defparam \phase_controller_slave.state_3_LC_5_25_1 .C_ON=1'b0;
    defparam \phase_controller_slave.state_3_LC_5_25_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_3_LC_5_25_1 .LUT_INIT=16'b1010000010101100;
    LogicCell40 \phase_controller_slave.state_3_LC_5_25_1  (
            .in0(N__12971),
            .in1(N__17265),
            .in2(N__12941),
            .in3(N__12961),
            .lcout(\phase_controller_slave.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20882),
            .ce(),
            .sr(N__20418));
    defparam \phase_controller_slave.state_2_LC_5_25_5 .C_ON=1'b0;
    defparam \phase_controller_slave.state_2_LC_5_25_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_2_LC_5_25_5 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \phase_controller_slave.state_2_LC_5_25_5  (
            .in0(N__17266),
            .in1(N__13289),
            .in2(N__13307),
            .in3(N__12962),
            .lcout(\phase_controller_slave.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20882),
            .ce(),
            .sr(N__20418));
    defparam \phase_controller_slave.start_timer_hc_LC_5_25_6 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_hc_LC_5_25_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.start_timer_hc_LC_5_25_6 .LUT_INIT=16'b1100110011001110;
    LogicCell40 \phase_controller_slave.start_timer_hc_LC_5_25_6  (
            .in0(N__12799),
            .in1(N__12947),
            .in2(N__13262),
            .in3(N__12940),
            .lcout(\phase_controller_slave.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20882),
            .ce(),
            .sr(N__20418));
    defparam \phase_controller_slave.start_timer_hc_RNO_0_LC_5_26_3 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_hc_RNO_0_LC_5_26_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.start_timer_hc_RNO_0_LC_5_26_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.start_timer_hc_RNO_0_LC_5_26_3  (
            .in0(_gnd_net_),
            .in1(N__13302),
            .in2(_gnd_net_),
            .in3(N__13282),
            .lcout(\phase_controller_slave.start_timer_hc_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D1_LC_7_12_0.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_7_12_0.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_7_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D1_LC_7_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13250),
            .lcout(il_max_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20937),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D1_LC_7_12_1.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_7_12_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_7_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MIN_D1_LC_7_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13235),
            .lcout(il_min_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20937),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D2_LC_7_12_7.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_7_12_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_7_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D2_LC_7_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13223),
            .lcout(il_max_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20937),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_7_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_7_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_1_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__16889),
            .in2(_gnd_net_),
            .in3(N__13204),
            .lcout(\phase_controller_inst1.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D2_LC_7_14_3.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_7_14_3.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_7_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D2_LC_7_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13166),
            .lcout(il_min_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20931),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D1_LC_7_14_5.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_7_14_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_7_14_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH1_MIN_D1_LC_7_14_5 (
            .in0(N__13184),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_min_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20931),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_RNIR0JF_1_LC_7_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNIR0JF_1_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNIR0JF_1_LC_7_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNIR0JF_1_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(N__19910),
            .in2(_gnd_net_),
            .in3(N__13150),
            .lcout(\phase_controller_inst1.T01_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_8_LC_7_17_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_8_LC_7_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_8_LC_7_17_0 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_8_LC_7_17_0  (
            .in0(N__15147),
            .in1(N__15330),
            .in2(N__14633),
            .in3(N__15459),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20914),
            .ce(),
            .sr(N__20374));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_7_LC_7_17_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_7_LC_7_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_7_LC_7_17_1 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_7_LC_7_17_1  (
            .in0(N__15458),
            .in1(N__15148),
            .in2(N__15346),
            .in3(N__14210),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20914),
            .ce(),
            .sr(N__20374));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_16_LC_7_18_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_16_LC_7_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_16_LC_7_18_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_16_LC_7_18_0  (
            .in0(N__15453),
            .in1(N__15135),
            .in2(N__15336),
            .in3(N__14969),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20908),
            .ce(),
            .sr(N__20379));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_12_LC_7_18_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_12_LC_7_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_12_LC_7_18_1 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_12_LC_7_18_1  (
            .in0(N__15130),
            .in1(N__15304),
            .in2(N__14528),
            .in3(N__15456),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20908),
            .ce(),
            .sr(N__20379));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_15_LC_7_18_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_15_LC_7_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_15_LC_7_18_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_15_LC_7_18_2  (
            .in0(N__15452),
            .in1(N__15134),
            .in2(N__15335),
            .in3(N__14450),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20908),
            .ce(),
            .sr(N__20379));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_14_LC_7_18_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_14_LC_7_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_14_LC_7_18_3 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_14_LC_7_18_3  (
            .in0(N__15132),
            .in1(N__15306),
            .in2(N__14477),
            .in3(N__15457),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20908),
            .ce(),
            .sr(N__20379));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_11_LC_7_18_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_11_LC_7_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_11_LC_7_18_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_11_LC_7_18_4  (
            .in0(N__15451),
            .in1(N__15133),
            .in2(N__15334),
            .in3(N__14555),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20908),
            .ce(),
            .sr(N__20379));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_13_LC_7_18_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_13_LC_7_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_13_LC_7_18_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_13_LC_7_18_5  (
            .in0(N__15131),
            .in1(N__15305),
            .in2(N__15478),
            .in3(N__14501),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20908),
            .ce(),
            .sr(N__20379));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_9_LC_7_18_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_9_LC_7_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_9_LC_7_18_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_9_LC_7_18_6  (
            .in0(N__15454),
            .in1(N__15136),
            .in2(N__15337),
            .in3(N__14606),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20908),
            .ce(),
            .sr(N__20379));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_10_LC_7_18_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_10_LC_7_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_10_LC_7_18_7 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_10_LC_7_18_7  (
            .in0(N__15129),
            .in1(N__15303),
            .in2(N__14582),
            .in3(N__15455),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20908),
            .ce(),
            .sr(N__20379));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_19_LC_7_19_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_19_LC_7_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_19_LC_7_19_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_19_LC_7_19_0  (
            .in0(N__15105),
            .in1(N__15434),
            .in2(N__15344),
            .in3(N__14894),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20904),
            .ce(),
            .sr(N__20384));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_17_LC_7_19_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_17_LC_7_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_17_LC_7_19_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_17_LC_7_19_6  (
            .in0(N__15104),
            .in1(N__15433),
            .in2(N__15343),
            .in3(N__14945),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20904),
            .ce(),
            .sr(N__20384));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_18_LC_7_19_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_18_LC_7_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_18_LC_7_19_7 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_18_LC_7_19_7  (
            .in0(N__15432),
            .in1(N__15320),
            .in2(N__15149),
            .in3(N__14921),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20904),
            .ce(),
            .sr(N__20384));
    defparam \phase_controller_slave.stoper_tr.stoper_state_1_LC_7_20_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_1_LC_7_20_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_1_LC_7_20_7 .LUT_INIT=16'b0010000001100100;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_1_LC_7_20_7  (
            .in0(N__15435),
            .in1(N__15107),
            .in2(N__15345),
            .in3(N__15184),
            .lcout(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20900),
            .ce(N__20190),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGUTL_6_LC_7_21_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGUTL_6_LC_7_21_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGUTL_6_LC_7_21_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGUTL_6_LC_7_21_0  (
            .in0(_gnd_net_),
            .in1(N__18845),
            .in2(_gnd_net_),
            .in3(N__18326),
            .lcout(\delay_measurement_inst.delay_hc_reg_3_0_a2_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_7_21_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_7_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_7_21_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_7_21_1  (
            .in0(N__15285),
            .in1(N__15420),
            .in2(_gnd_net_),
            .in3(N__15103),
            .lcout(\phase_controller_slave.stoper_tr.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_7_21_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_7_21_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_7_21_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_7_21_3  (
            .in0(_gnd_net_),
            .in1(N__18373),
            .in2(_gnd_net_),
            .in3(N__18415),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_232_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D2_LC_7_21_7.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_7_21_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_7_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MIN_D2_LC_7_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13430),
            .lcout(il_min_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20896),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_esr_5_LC_7_22_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_5_LC_7_22_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_5_LC_7_22_0 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_5_LC_7_22_0  (
            .in0(N__15831),
            .in1(N__13670),
            .in2(N__15539),
            .in3(N__18377),
            .lcout(measured_delay_hc_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20889),
            .ce(N__15740),
            .sr(N__20400));
    defparam \delay_measurement_inst.delay_hc_reg_esr_2_LC_7_22_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_2_LC_7_22_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_2_LC_7_22_1 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_2_LC_7_22_1  (
            .in0(N__15002),
            .in1(N__15532),
            .in2(N__13673),
            .in3(N__15829),
            .lcout(measured_delay_hc_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20889),
            .ce(N__15740),
            .sr(N__20400));
    defparam \delay_measurement_inst.delay_hc_reg_esr_11_LC_7_22_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_11_LC_7_22_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_11_LC_7_22_2 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_11_LC_7_22_2  (
            .in0(N__15802),
            .in1(N__19569),
            .in2(_gnd_net_),
            .in3(N__19046),
            .lcout(measured_delay_hc_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20889),
            .ce(N__15740),
            .sr(N__20400));
    defparam \delay_measurement_inst.delay_hc_reg_esr_12_LC_7_22_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_12_LC_7_22_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_12_LC_7_22_3 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_12_LC_7_22_3  (
            .in0(N__19568),
            .in1(N__15803),
            .in2(_gnd_net_),
            .in3(N__19007),
            .lcout(measured_delay_hc_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20889),
            .ce(N__15740),
            .sr(N__20400));
    defparam \delay_measurement_inst.delay_hc_reg_ess_3_LC_7_22_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_ess_3_LC_7_22_4 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_hc_reg_ess_3_LC_7_22_4 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_ess_3_LC_7_22_4  (
            .in0(N__15833),
            .in1(N__15538),
            .in2(N__18467),
            .in3(N__13672),
            .lcout(measured_delay_hc_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20889),
            .ce(N__15740),
            .sr(N__20400));
    defparam \delay_measurement_inst.delay_hc_reg_esr_4_LC_7_22_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_4_LC_7_22_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_4_LC_7_22_5 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_4_LC_7_22_5  (
            .in0(N__13669),
            .in1(N__15533),
            .in2(N__18425),
            .in3(N__15830),
            .lcout(measured_delay_hc_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20889),
            .ce(N__15740),
            .sr(N__20400));
    defparam \delay_measurement_inst.delay_hc_reg_ess_1_LC_7_22_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_ess_1_LC_7_22_6 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_hc_reg_ess_1_LC_7_22_6 .LUT_INIT=16'b1111000010000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_ess_1_LC_7_22_6  (
            .in0(N__15832),
            .in1(N__13671),
            .in2(N__15035),
            .in3(N__15537),
            .lcout(measured_delay_hc_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20889),
            .ce(N__15740),
            .sr(N__20400));
    defparam \delay_measurement_inst.delay_hc_reg_esr_10_LC_7_22_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_10_LC_7_22_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_10_LC_7_22_7 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_10_LC_7_22_7  (
            .in0(N__19567),
            .in1(N__15801),
            .in2(_gnd_net_),
            .in3(N__19085),
            .lcout(measured_delay_hc_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20889),
            .ce(N__15740),
            .sr(N__20400));
    defparam \delay_measurement_inst.delay_hc_reg_esr_9_LC_7_23_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_9_LC_7_23_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_9_LC_7_23_0 .LUT_INIT=16'b0011000000110001;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_9_LC_7_23_0  (
            .in0(N__19558),
            .in1(N__15548),
            .in2(N__19154),
            .in3(N__15800),
            .lcout(measured_delay_hc_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20883),
            .ce(N__15732),
            .sr(N__20408));
    defparam \delay_measurement_inst.delay_hc_reg_esr_15_LC_7_23_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_15_LC_7_23_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_15_LC_7_23_1 .LUT_INIT=16'b1100000011001000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_15_LC_7_23_1  (
            .in0(N__15500),
            .in1(N__18853),
            .in2(N__19571),
            .in3(N__19829),
            .lcout(measured_delay_hc_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20883),
            .ce(N__15732),
            .sr(N__20408));
    defparam \delay_measurement_inst.delay_hc_reg_esr_19_LC_7_23_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_19_LC_7_23_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_19_LC_7_23_2 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_19_LC_7_23_2  (
            .in0(N__19826),
            .in1(N__19562),
            .in2(_gnd_net_),
            .in3(N__19309),
            .lcout(measured_delay_hc_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20883),
            .ce(N__15732),
            .sr(N__20408));
    defparam \delay_measurement_inst.delay_hc_reg_esr_6_LC_7_23_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_6_LC_7_23_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_6_LC_7_23_3 .LUT_INIT=16'b1111010011110101;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_6_LC_7_23_3  (
            .in0(N__15529),
            .in1(N__18854),
            .in2(N__18335),
            .in3(N__15828),
            .lcout(measured_delay_hc_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20883),
            .ce(N__15732),
            .sr(N__20408));
    defparam \delay_measurement_inst.delay_hc_reg_esr_17_LC_7_23_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_17_LC_7_23_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_17_LC_7_23_4 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_17_LC_7_23_4  (
            .in0(N__19825),
            .in1(N__19561),
            .in2(_gnd_net_),
            .in3(N__19408),
            .lcout(measured_delay_hc_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20883),
            .ce(N__15732),
            .sr(N__20408));
    defparam \delay_measurement_inst.delay_hc_reg_esr_16_LC_7_23_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_16_LC_7_23_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_16_LC_7_23_5 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_16_LC_7_23_5  (
            .in0(N__19559),
            .in1(N__19459),
            .in2(_gnd_net_),
            .in3(N__19827),
            .lcout(measured_delay_hc_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20883),
            .ce(N__15732),
            .sr(N__20408));
    defparam \delay_measurement_inst.delay_hc_reg_esr_14_LC_7_23_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_14_LC_7_23_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_14_LC_7_23_6 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_14_LC_7_23_6  (
            .in0(N__19557),
            .in1(N__15799),
            .in2(_gnd_net_),
            .in3(N__18916),
            .lcout(measured_delay_hc_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20883),
            .ce(N__15732),
            .sr(N__20408));
    defparam \delay_measurement_inst.delay_hc_reg_esr_18_LC_7_23_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_18_LC_7_23_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_18_LC_7_23_7 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_18_LC_7_23_7  (
            .in0(N__19560),
            .in1(N__19355),
            .in2(_gnd_net_),
            .in3(N__19828),
            .lcout(measured_delay_hc_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20883),
            .ce(N__15732),
            .sr(N__20408));
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_7_24_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_7_24_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_7_24_0 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_7_LC_7_24_0  (
            .in0(N__13871),
            .in1(N__15530),
            .in2(N__18281),
            .in3(N__15559),
            .lcout(measured_delay_hc_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20876),
            .ce(),
            .sr(N__20412));
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_7_24_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_7_24_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_7_24_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_8_LC_7_24_2  (
            .in0(N__13838),
            .in1(N__15531),
            .in2(N__18236),
            .in3(N__15560),
            .lcout(measured_delay_hc_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20876),
            .ce(),
            .sr(N__20412));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_8_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_8_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_8_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_8_13_0  (
            .in0(N__17559),
            .in1(N__17232),
            .in2(_gnd_net_),
            .in3(N__13808),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__20932),
            .ce(N__14171),
            .sr(N__20353));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_8_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_8_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_8_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_8_13_1  (
            .in0(N__17554),
            .in1(N__17211),
            .in2(_gnd_net_),
            .in3(N__13805),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__20932),
            .ce(N__14171),
            .sr(N__20353));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_8_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_8_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_8_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_8_13_2  (
            .in0(N__17560),
            .in1(N__15657),
            .in2(_gnd_net_),
            .in3(N__14126),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__20932),
            .ce(N__14171),
            .sr(N__20353));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_8_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_8_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_8_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_8_13_3  (
            .in0(N__17555),
            .in1(N__15633),
            .in2(_gnd_net_),
            .in3(N__14123),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__20932),
            .ce(N__14171),
            .sr(N__20353));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_8_13_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_8_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_8_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_8_13_4  (
            .in0(N__17561),
            .in1(N__15611),
            .in2(_gnd_net_),
            .in3(N__14120),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__20932),
            .ce(N__14171),
            .sr(N__20353));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_8_13_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_8_13_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_8_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_8_13_5  (
            .in0(N__17556),
            .in1(N__16037),
            .in2(_gnd_net_),
            .in3(N__14117),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__20932),
            .ce(N__14171),
            .sr(N__20353));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_8_13_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_8_13_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_8_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_8_13_6  (
            .in0(N__17558),
            .in1(N__16017),
            .in2(_gnd_net_),
            .in3(N__14114),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__20932),
            .ce(N__14171),
            .sr(N__20353));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_8_13_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_8_13_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_8_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_8_13_7  (
            .in0(N__17557),
            .in1(N__15993),
            .in2(_gnd_net_),
            .in3(N__14111),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__20932),
            .ce(N__14171),
            .sr(N__20353));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_8_14_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_8_14_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_8_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_8_14_0  (
            .in0(N__17532),
            .in1(N__15970),
            .in2(_gnd_net_),
            .in3(N__14108),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__20925),
            .ce(N__14172),
            .sr(N__20355));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_8_14_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_8_14_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_8_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_8_14_1  (
            .in0(N__17567),
            .in1(N__15949),
            .in2(_gnd_net_),
            .in3(N__14105),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__20925),
            .ce(N__14172),
            .sr(N__20355));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_8_14_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_8_14_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_8_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_8_14_2  (
            .in0(N__17529),
            .in1(N__15927),
            .in2(_gnd_net_),
            .in3(N__14102),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__20925),
            .ce(N__14172),
            .sr(N__20355));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_8_14_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_8_14_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_8_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_8_14_3  (
            .in0(N__17564),
            .in1(N__15903),
            .in2(_gnd_net_),
            .in3(N__14156),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__20925),
            .ce(N__14172),
            .sr(N__20355));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_8_14_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_8_14_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_8_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_8_14_4  (
            .in0(N__17530),
            .in1(N__15881),
            .in2(_gnd_net_),
            .in3(N__14153),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__20925),
            .ce(N__14172),
            .sr(N__20355));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_8_14_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_8_14_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_8_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_8_14_5  (
            .in0(N__17565),
            .in1(N__15863),
            .in2(_gnd_net_),
            .in3(N__14150),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__20925),
            .ce(N__14172),
            .sr(N__20355));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_8_14_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_8_14_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_8_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_8_14_6  (
            .in0(N__17531),
            .in1(N__16209),
            .in2(_gnd_net_),
            .in3(N__14147),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__20925),
            .ce(N__14172),
            .sr(N__20355));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_8_14_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_8_14_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_8_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_8_14_7  (
            .in0(N__17566),
            .in1(N__16185),
            .in2(_gnd_net_),
            .in3(N__14144),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__20925),
            .ce(N__14172),
            .sr(N__20355));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_8_15_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_8_15_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_8_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_8_15_0  (
            .in0(N__17542),
            .in1(N__16162),
            .in2(_gnd_net_),
            .in3(N__14141),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_8_15_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__20921),
            .ce(N__14173),
            .sr(N__20361));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_8_15_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_8_15_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_8_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_8_15_1  (
            .in0(N__17546),
            .in1(N__16141),
            .in2(_gnd_net_),
            .in3(N__14138),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__20921),
            .ce(N__14173),
            .sr(N__20361));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_8_15_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_8_15_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_8_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_8_15_2  (
            .in0(N__17543),
            .in1(N__16119),
            .in2(_gnd_net_),
            .in3(N__14135),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__20921),
            .ce(N__14173),
            .sr(N__20361));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_8_15_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_8_15_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_8_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_8_15_3  (
            .in0(N__17547),
            .in1(N__16095),
            .in2(_gnd_net_),
            .in3(N__14132),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__20921),
            .ce(N__14173),
            .sr(N__20361));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_8_15_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_8_15_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_8_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_8_15_4  (
            .in0(N__17544),
            .in1(N__16073),
            .in2(_gnd_net_),
            .in3(N__14129),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__20921),
            .ce(N__14173),
            .sr(N__20361));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_8_15_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_8_15_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_8_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_8_15_5  (
            .in0(N__17548),
            .in1(N__16055),
            .in2(_gnd_net_),
            .in3(N__14201),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__20921),
            .ce(N__14173),
            .sr(N__20361));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_8_15_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_8_15_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_8_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_8_15_6  (
            .in0(N__17545),
            .in1(N__16374),
            .in2(_gnd_net_),
            .in3(N__14198),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__20921),
            .ce(N__14173),
            .sr(N__20361));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_8_15_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_8_15_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_8_15_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_8_15_7  (
            .in0(N__17549),
            .in1(N__16350),
            .in2(_gnd_net_),
            .in3(N__14195),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__20921),
            .ce(N__14173),
            .sr(N__20361));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_8_16_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_8_16_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_8_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_8_16_0  (
            .in0(N__17550),
            .in1(N__16327),
            .in2(_gnd_net_),
            .in3(N__14192),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_8_16_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__20915),
            .ce(N__14174),
            .sr(N__20369));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_8_16_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_8_16_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_8_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_8_16_1  (
            .in0(N__17562),
            .in1(N__16306),
            .in2(_gnd_net_),
            .in3(N__14189),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__20915),
            .ce(N__14174),
            .sr(N__20369));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_8_16_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_8_16_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_8_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_8_16_2  (
            .in0(N__17551),
            .in1(N__16272),
            .in2(_gnd_net_),
            .in3(N__14186),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__20915),
            .ce(N__14174),
            .sr(N__20369));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_8_16_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_8_16_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_8_16_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_8_16_3  (
            .in0(N__17563),
            .in1(N__16236),
            .in2(_gnd_net_),
            .in3(N__14183),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__20915),
            .ce(N__14174),
            .sr(N__20369));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_8_16_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_8_16_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_8_16_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_8_16_4  (
            .in0(N__17552),
            .in1(N__16286),
            .in2(_gnd_net_),
            .in3(N__14180),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__20915),
            .ce(N__14174),
            .sr(N__20369));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_8_16_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_8_16_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_8_16_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_8_16_5  (
            .in0(N__16250),
            .in1(N__17553),
            .in2(_gnd_net_),
            .in3(N__14177),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20915),
            .ce(N__14174),
            .sr(N__20369));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_8_17_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_8_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_8_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_8_17_0  (
            .in0(_gnd_net_),
            .in1(N__14440),
            .in2(N__14417),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_17_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_8_17_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_8_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_8_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_8_17_1  (
            .in0(_gnd_net_),
            .in1(N__14402),
            .in2(_gnd_net_),
            .in3(N__14375),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_8_17_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_8_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_8_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_8_17_2  (
            .in0(_gnd_net_),
            .in1(N__14372),
            .in2(N__14357),
            .in3(N__14330),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_8_17_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_8_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_8_17_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_8_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14327),
            .in3(N__14297),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_8_17_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_8_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_8_17_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_8_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14294),
            .in3(N__14261),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_8_17_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_8_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_8_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_8_17_5  (
            .in0(_gnd_net_),
            .in1(N__14258),
            .in2(_gnd_net_),
            .in3(N__14228),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_8_17_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_8_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_8_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_8_17_6  (
            .in0(_gnd_net_),
            .in1(N__14224),
            .in2(_gnd_net_),
            .in3(N__14204),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_8_17_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_8_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_8_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_8_17_7  (
            .in0(_gnd_net_),
            .in1(N__14650),
            .in2(_gnd_net_),
            .in3(N__14624),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_8_18_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_8_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_8_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_8_18_0  (
            .in0(_gnd_net_),
            .in1(N__14620),
            .in2(_gnd_net_),
            .in3(N__14600),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9 ),
            .ltout(),
            .carryin(bfn_8_18_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_8_18_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_8_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_8_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_8_18_1  (
            .in0(_gnd_net_),
            .in1(N__14596),
            .in2(_gnd_net_),
            .in3(N__14573),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_8_18_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_8_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_8_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_8_18_2  (
            .in0(_gnd_net_),
            .in1(N__14569),
            .in2(_gnd_net_),
            .in3(N__14549),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_8_18_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_8_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_8_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_8_18_3  (
            .in0(_gnd_net_),
            .in1(N__14542),
            .in2(_gnd_net_),
            .in3(N__14519),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_8_18_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_8_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_8_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_8_18_4  (
            .in0(_gnd_net_),
            .in1(N__14515),
            .in2(_gnd_net_),
            .in3(N__14495),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_8_18_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_8_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_8_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_8_18_5  (
            .in0(_gnd_net_),
            .in1(N__14491),
            .in2(_gnd_net_),
            .in3(N__14468),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_8_18_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_8_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_8_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_8_18_6  (
            .in0(_gnd_net_),
            .in1(N__14464),
            .in2(_gnd_net_),
            .in3(N__14444),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_8_18_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_8_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_8_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_8_18_7  (
            .in0(_gnd_net_),
            .in1(N__14983),
            .in2(_gnd_net_),
            .in3(N__14963),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_8_19_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_8_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_8_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_8_19_0  (
            .in0(_gnd_net_),
            .in1(N__14959),
            .in2(_gnd_net_),
            .in3(N__14939),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17 ),
            .ltout(),
            .carryin(bfn_8_19_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_8_19_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_8_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_8_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_8_19_1  (
            .in0(_gnd_net_),
            .in1(N__14935),
            .in2(_gnd_net_),
            .in3(N__14915),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_8_19_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_8_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_8_19_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_8_19_2  (
            .in0(_gnd_net_),
            .in1(N__14911),
            .in2(_gnd_net_),
            .in3(N__14897),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_8_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_8_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_8_19_3 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_8_19_3  (
            .in0(N__16401),
            .in1(N__16449),
            .in2(_gnd_net_),
            .in3(N__17085),
            .lcout(\phase_controller_inst1.stoper_tr.N_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_8_19_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_8_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_8_19_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_8_19_4  (
            .in0(_gnd_net_),
            .in1(N__15398),
            .in2(_gnd_net_),
            .in3(N__15074),
            .lcout(\phase_controller_slave.stoper_tr.time_passed11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_8_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_8_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_8_19_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_8_19_5  (
            .in0(N__16548),
            .in1(N__16964),
            .in2(_gnd_net_),
            .in3(N__17111),
            .lcout(\phase_controller_inst1.stoper_tr.N_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_8_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_8_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_8_19_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_8_19_6  (
            .in0(N__16698),
            .in1(N__16778),
            .in2(N__18546),
            .in3(N__16737),
            .lcout(\phase_controller_inst1.stoper_tr.N_32 ),
            .ltout(\phase_controller_inst1.stoper_tr.N_32_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_8_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_8_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_8_19_7 .LUT_INIT=16'b1111001111110001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_8_19_7  (
            .in0(N__17022),
            .in1(N__16965),
            .in2(N__14726),
            .in3(N__16493),
            .lcout(\phase_controller_inst1.stoper_tr.N_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.stoper_state_0_LC_8_20_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_0_LC_8_20_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_0_LC_8_20_2 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_0_LC_8_20_2  (
            .in0(N__15436),
            .in1(N__15106),
            .in2(N__15347),
            .in3(N__15185),
            .lcout(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20897),
            .ce(N__20189),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_8_21_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_8_21_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_8_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_8_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18443),
            .lcout(\delay_measurement_inst.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20890),
            .ce(N__19496),
            .sr(N__20392));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_8_21_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_8_21_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_8_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_8_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18485),
            .lcout(\delay_measurement_inst.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20890),
            .ce(N__19496),
            .sr(N__20392));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNID3EH4_1_LC_8_22_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNID3EH4_1_LC_8_22_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNID3EH4_1_LC_8_22_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNID3EH4_1_LC_8_22_0  (
            .in0(N__15008),
            .in1(N__15498),
            .in2(N__15017),
            .in3(N__15590),
            .lcout(\delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_8_22_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_8_22_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_8_22_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_8_22_1  (
            .in0(N__19003),
            .in1(N__19045),
            .in2(N__18964),
            .in3(N__19084),
            .lcout(\delay_measurement_inst.N_243 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_6_LC_8_22_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_6_LC_8_22_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_6_LC_8_22_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_6_LC_8_22_2  (
            .in0(_gnd_net_),
            .in1(N__19145),
            .in2(_gnd_net_),
            .in3(N__18331),
            .lcout(\delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3GIH1_1_LC_8_22_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3GIH1_1_LC_8_22_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3GIH1_1_LC_8_22_3 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3GIH1_1_LC_8_22_3  (
            .in0(N__18910),
            .in1(N__18462),
            .in2(N__15034),
            .in3(N__15001),
            .lcout(\delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3HO31_6_LC_8_22_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3HO31_6_LC_8_22_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3HO31_6_LC_8_22_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3HO31_6_LC_8_22_4  (
            .in0(N__18837),
            .in1(N__19144),
            .in2(_gnd_net_),
            .in3(N__18330),
            .lcout(\delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0TRB1_18_LC_8_22_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0TRB1_18_LC_8_22_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0TRB1_18_LC_8_22_5 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0TRB1_18_LC_8_22_5  (
            .in0(N__19347),
            .in1(N__18463),
            .in2(N__19310),
            .in3(N__15000),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0QNN2_16_LC_8_22_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0QNN2_16_LC_8_22_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0QNN2_16_LC_8_22_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0QNN2_16_LC_8_22_6  (
            .in0(N__19404),
            .in1(N__19460),
            .in2(N__15593),
            .in3(N__15589),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2PJ34_14_LC_8_22_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2PJ34_14_LC_8_22_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2PJ34_14_LC_8_22_7 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2PJ34_14_LC_8_22_7  (
            .in0(N__15581),
            .in1(N__18911),
            .in2(N__15575),
            .in3(N__18838),
            .lcout(\delay_measurement_inst.delay_hc_timer.un3_elapsed_time_hc_0_a4_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4ESID_31_LC_8_23_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4ESID_31_LC_8_23_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4ESID_31_LC_8_23_0 .LUT_INIT=16'b0000000100001111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4ESID_31_LC_8_23_0  (
            .in0(N__15572),
            .in1(N__15566),
            .in2(N__19570),
            .in3(N__15827),
            .lcout(\delay_measurement_inst.un3_elapsed_time_hc_0_i ),
            .ltout(\delay_measurement_inst.un3_elapsed_time_hc_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBNQQD_31_LC_8_23_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBNQQD_31_LC_8_23_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBNQQD_31_LC_8_23_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBNQQD_31_LC_8_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15551),
            .in3(N__20463),
            .lcout(\delay_measurement_inst.un3_elapsed_time_hc_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_esr_RNO_0_9_LC_8_23_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_RNO_0_9_LC_8_23_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_RNO_0_9_LC_8_23_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_RNO_0_9_LC_8_23_2  (
            .in0(N__19824),
            .in1(N__15845),
            .in2(N__19153),
            .in3(N__18851),
            .lcout(\delay_measurement_inst.N_219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4TEU1_14_LC_8_23_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4TEU1_14_LC_8_23_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4TEU1_14_LC_8_23_3 .LUT_INIT=16'b0000001100100011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4TEU1_14_LC_8_23_3  (
            .in0(N__15844),
            .in1(N__18839),
            .in2(N__18917),
            .in3(N__19146),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.N_237_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE5L06_31_LC_8_23_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE5L06_31_LC_8_23_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE5L06_31_LC_8_23_4 .LUT_INIT=16'b1101110111011100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE5L06_31_LC_8_23_4  (
            .in0(N__19823),
            .in1(N__19566),
            .in2(N__15542),
            .in3(N__15499),
            .lcout(\delay_measurement_inst.N_209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_8_23_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_8_23_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_8_23_5 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_8_23_5  (
            .in0(N__19458),
            .in1(N__19308),
            .in2(N__19409),
            .in3(N__19354),
            .lcout(\delay_measurement_inst.N_207 ),
            .ltout(\delay_measurement_inst.N_207_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBM7A4_14_LC_8_23_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBM7A4_14_LC_8_23_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBM7A4_14_LC_8_23_6 .LUT_INIT=16'b0101000001010001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBM7A4_14_LC_8_23_6  (
            .in0(N__19822),
            .in1(N__18852),
            .in2(N__15482),
            .in3(N__18915),
            .lcout(\delay_measurement_inst.N_216_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN2LL4_7_LC_8_23_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN2LL4_7_LC_8_23_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN2LL4_7_LC_8_23_7 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN2LL4_7_LC_8_23_7  (
            .in0(N__15843),
            .in1(N__18277),
            .in2(N__18235),
            .in3(N__19821),
            .lcout(\delay_measurement_inst.N_247 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_esr_13_LC_8_24_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_13_LC_8_24_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_13_LC_8_24_1 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_13_LC_8_24_1  (
            .in0(N__19553),
            .in1(N__15798),
            .in2(_gnd_net_),
            .in3(N__18965),
            .lcout(measured_delay_hc_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20871),
            .ce(N__15739),
            .sr(N__20409));
    defparam \phase_controller_slave.S2_LC_8_26_3 .C_ON=1'b0;
    defparam \phase_controller_slave.S2_LC_8_26_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.S2_LC_8_26_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.S2_LC_8_26_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15706),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20866),
            .ce(),
            .sr(N__20414));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_9_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_9_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_9_13_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__17233),
            .in2(N__15658),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__20926),
            .ce(N__17194),
            .sr(N__20352));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_9_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_9_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_9_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(N__17212),
            .in2(N__15634),
            .in3(N__15662),
            .lcout(\delay_measurement_inst.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__20926),
            .ce(N__17194),
            .sr(N__20352));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_9_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_9_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_9_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__15609),
            .in2(N__15659),
            .in3(N__15638),
            .lcout(\delay_measurement_inst.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__20926),
            .ce(N__17194),
            .sr(N__20352));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_9_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_9_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_9_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__16035),
            .in2(N__15635),
            .in3(N__15614),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__20926),
            .ce(N__17194),
            .sr(N__20352));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_9_13_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_9_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_9_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(N__15610),
            .in2(N__16018),
            .in3(N__15596),
            .lcout(\delay_measurement_inst.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__20926),
            .ce(N__17194),
            .sr(N__20352));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_9_13_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_9_13_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_9_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(N__16036),
            .in2(N__15994),
            .in3(N__16022),
            .lcout(\delay_measurement_inst.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__20926),
            .ce(N__17194),
            .sr(N__20352));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_9_13_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_9_13_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_9_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__15969),
            .in2(N__16019),
            .in3(N__15998),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__20926),
            .ce(N__17194),
            .sr(N__20352));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_9_13_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_9_13_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_9_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(N__15948),
            .in2(N__15995),
            .in3(N__15974),
            .lcout(\delay_measurement_inst.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__20926),
            .ce(N__17194),
            .sr(N__20352));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_9_14_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_9_14_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_9_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__15971),
            .in2(N__15928),
            .in3(N__15953),
            .lcout(\delay_measurement_inst.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__20922),
            .ce(N__17193),
            .sr(N__20354));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_9_14_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_9_14_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_9_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__15950),
            .in2(N__15904),
            .in3(N__15932),
            .lcout(\delay_measurement_inst.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__20922),
            .ce(N__17193),
            .sr(N__20354));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_9_14_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_9_14_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_9_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(N__15879),
            .in2(N__15929),
            .in3(N__15908),
            .lcout(\delay_measurement_inst.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__20922),
            .ce(N__17193),
            .sr(N__20354));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_9_14_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_9_14_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_9_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__15861),
            .in2(N__15905),
            .in3(N__15884),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__20922),
            .ce(N__17193),
            .sr(N__20354));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_9_14_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_9_14_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_9_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(N__15880),
            .in2(N__16210),
            .in3(N__15866),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__20922),
            .ce(N__17193),
            .sr(N__20354));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_9_14_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_9_14_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_9_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(N__15862),
            .in2(N__16186),
            .in3(N__15848),
            .lcout(\delay_measurement_inst.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__20922),
            .ce(N__17193),
            .sr(N__20354));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_9_14_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_9_14_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_9_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__16161),
            .in2(N__16211),
            .in3(N__16190),
            .lcout(\delay_measurement_inst.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__20922),
            .ce(N__17193),
            .sr(N__20354));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_9_14_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_9_14_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_9_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(N__16140),
            .in2(N__16187),
            .in3(N__16166),
            .lcout(\delay_measurement_inst.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__20922),
            .ce(N__17193),
            .sr(N__20354));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_9_15_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_9_15_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_9_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__16163),
            .in2(N__16120),
            .in3(N__16145),
            .lcout(\delay_measurement_inst.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__20916),
            .ce(N__17192),
            .sr(N__20356));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_9_15_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_9_15_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_9_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__16142),
            .in2(N__16096),
            .in3(N__16124),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__20916),
            .ce(N__17192),
            .sr(N__20356));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_9_15_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_9_15_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_9_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__16071),
            .in2(N__16121),
            .in3(N__16100),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__20916),
            .ce(N__17192),
            .sr(N__20356));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_9_15_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_9_15_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_9_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__16053),
            .in2(N__16097),
            .in3(N__16076),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__20916),
            .ce(N__17192),
            .sr(N__20356));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_9_15_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_9_15_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_9_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(N__16072),
            .in2(N__16375),
            .in3(N__16058),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__20916),
            .ce(N__17192),
            .sr(N__20356));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_9_15_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_9_15_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_9_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(N__16054),
            .in2(N__16351),
            .in3(N__16040),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__20916),
            .ce(N__17192),
            .sr(N__20356));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_9_15_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_9_15_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_9_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(N__16326),
            .in2(N__16376),
            .in3(N__16355),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__20916),
            .ce(N__17192),
            .sr(N__20356));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_9_15_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_9_15_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_9_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(N__16305),
            .in2(N__16352),
            .in3(N__16331),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__20916),
            .ce(N__17192),
            .sr(N__20356));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_9_16_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_9_16_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_9_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(N__16328),
            .in2(N__16273),
            .in3(N__16310),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_9_16_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__20909),
            .ce(N__17191),
            .sr(N__20362));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_9_16_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_9_16_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_9_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(N__16307),
            .in2(N__16237),
            .in3(N__16289),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__20909),
            .ce(N__17191),
            .sr(N__20362));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_9_16_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_9_16_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_9_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(N__16285),
            .in2(N__16274),
            .in3(N__16253),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__20909),
            .ce(N__17191),
            .sr(N__20362));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_9_16_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_9_16_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_9_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(N__16249),
            .in2(N__16238),
            .in3(N__16217),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__20909),
            .ce(N__17191),
            .sr(N__20362));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_9_16_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_9_16_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_9_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16214),
            .lcout(\delay_measurement_inst.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20909),
            .ce(N__17191),
            .sr(N__20362));
    defparam \delay_measurement_inst.delay_tr_reg_esr_15_LC_9_17_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_15_LC_9_17_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_15_LC_9_17_0 .LUT_INIT=16'b1100000011001000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_15_LC_9_17_0  (
            .in0(N__18023),
            .in1(N__17941),
            .in2(N__18688),
            .in3(N__18579),
            .lcout(measured_delay_tr_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20905),
            .ce(N__18501),
            .sr(N__20370));
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_9_17_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_9_17_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_9_17_1 .LUT_INIT=16'b0010001000100011;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_9_LC_9_17_1  (
            .in0(N__18105),
            .in1(N__18203),
            .in2(N__18689),
            .in3(N__18147),
            .lcout(measured_delay_tr_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20905),
            .ce(N__18501),
            .sr(N__20370));
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_9_17_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_9_17_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_9_17_2 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_4_LC_9_17_2  (
            .in0(N__18193),
            .in1(N__18775),
            .in2(N__17903),
            .in3(N__17417),
            .lcout(measured_delay_tr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20905),
            .ce(N__18501),
            .sr(N__20370));
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_9_17_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_9_17_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_9_17_3 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_5_LC_9_17_3  (
            .in0(N__18776),
            .in1(N__18194),
            .in2(N__17438),
            .in3(N__17899),
            .lcout(measured_delay_tr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20905),
            .ce(N__18501),
            .sr(N__20370));
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_9_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_9_17_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_9_17_4 .LUT_INIT=16'b1111000011111101;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_6_LC_9_17_4  (
            .in0(N__18195),
            .in1(N__17942),
            .in2(N__17981),
            .in3(N__18777),
            .lcout(measured_delay_tr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20905),
            .ce(N__18501),
            .sr(N__20370));
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_9_17_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_9_17_5 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_9_17_5 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_ess_1_LC_9_17_5  (
            .in0(N__18778),
            .in1(N__18196),
            .in2(N__17375),
            .in3(N__17900),
            .lcout(measured_delay_tr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20905),
            .ce(N__18501),
            .sr(N__20370));
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_9_17_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_9_17_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_9_17_6 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_2_LC_9_17_6  (
            .in0(N__18192),
            .in1(N__18774),
            .in2(N__17902),
            .in3(N__17348),
            .lcout(measured_delay_tr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20905),
            .ce(N__18501),
            .sr(N__20370));
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_9_17_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_9_17_7 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_9_17_7 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_ess_3_LC_9_17_7  (
            .in0(N__18779),
            .in1(N__18197),
            .in2(N__17402),
            .in3(N__17901),
            .lcout(measured_delay_tr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20905),
            .ce(N__18501),
            .sr(N__20370));
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_9_18_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_9_18_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_9_18_0 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_10_LC_9_18_0  (
            .in0(N__18676),
            .in1(N__18148),
            .in2(_gnd_net_),
            .in3(N__17654),
            .lcout(measured_delay_tr_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20901),
            .ce(N__18505),
            .sr(N__20372));
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_9_18_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_9_18_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_9_18_1 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_12_LC_9_18_1  (
            .in0(N__18150),
            .in1(N__18678),
            .in2(_gnd_net_),
            .in3(N__17716),
            .lcout(measured_delay_tr_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20901),
            .ce(N__18505),
            .sr(N__20372));
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_9_18_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_9_18_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_9_18_2 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_16_LC_9_18_2  (
            .in0(N__18681),
            .in1(N__17792),
            .in2(_gnd_net_),
            .in3(N__18591),
            .lcout(measured_delay_tr_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20901),
            .ce(N__18505),
            .sr(N__20372));
    defparam \delay_measurement_inst.delay_tr_reg_esr_14_LC_9_18_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_14_LC_9_18_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_14_LC_9_18_3 .LUT_INIT=16'b1010101110101011;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_14_LC_9_18_3  (
            .in0(N__18059),
            .in1(N__18680),
            .in2(N__18155),
            .in3(_gnd_net_),
            .lcout(measured_delay_tr_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20901),
            .ce(N__18505),
            .sr(N__20372));
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_9_18_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_9_18_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_9_18_4 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_17_LC_9_18_4  (
            .in0(N__17774),
            .in1(N__18683),
            .in2(_gnd_net_),
            .in3(N__18592),
            .lcout(measured_delay_tr_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20901),
            .ce(N__18505),
            .sr(N__20372));
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_9_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_9_18_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_9_18_5 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_18_LC_9_18_5  (
            .in0(N__18593),
            .in1(N__18682),
            .in2(_gnd_net_),
            .in3(N__17750),
            .lcout(measured_delay_tr_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20901),
            .ce(N__18505),
            .sr(N__20372));
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_9_18_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_9_18_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_9_18_6 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_11_LC_9_18_6  (
            .in0(N__18677),
            .in1(N__18149),
            .in2(_gnd_net_),
            .in3(N__17695),
            .lcout(measured_delay_tr_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20901),
            .ce(N__18505),
            .sr(N__20372));
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_9_18_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_9_18_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_9_18_7 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_13_LC_9_18_7  (
            .in0(N__18151),
            .in1(N__18679),
            .in2(_gnd_net_),
            .in3(N__17675),
            .lcout(measured_delay_tr_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20901),
            .ce(N__18505),
            .sr(N__20372));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_9_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_9_19_0 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_9_19_0  (
            .in0(N__16807),
            .in1(_gnd_net_),
            .in2(N__17850),
            .in3(N__18707),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_9_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_9_19_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_9_19_1  (
            .in0(N__16782),
            .in1(N__16736),
            .in2(N__18527),
            .in3(N__16697),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_9_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_9_19_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_9_19_4  (
            .in0(N__16665),
            .in1(N__16638),
            .in2(N__16611),
            .in3(N__16576),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_0_6 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_9_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_9_19_5 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_9_19_5  (
            .in0(N__16515),
            .in1(_gnd_net_),
            .in2(N__16496),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_9 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_9_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_9_19_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_9_19_6  (
            .in0(N__16904),
            .in1(N__17120),
            .in2(N__17114),
            .in3(N__17110),
            .lcout(\phase_controller_inst1.stoper_tr.N_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_9_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_9_19_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_9_19_7  (
            .in0(N__17061),
            .in1(N__17016),
            .in2(N__16963),
            .in3(N__16920),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.S1_LC_9_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_9_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_9_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S1_LC_9_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16898),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20891),
            .ce(),
            .sr(N__20380));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_9_21_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_9_21_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_9_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_9_21_0  (
            .in0(N__20523),
            .in1(N__18483),
            .in2(_gnd_net_),
            .in3(N__16838),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_9_21_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__20884),
            .ce(N__20651),
            .sr(N__20385));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_9_21_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_9_21_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_9_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_9_21_1  (
            .in0(N__20582),
            .in1(N__18441),
            .in2(_gnd_net_),
            .in3(N__16835),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__20884),
            .ce(N__20651),
            .sr(N__20385));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_9_21_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_9_21_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_9_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_9_21_2  (
            .in0(N__20524),
            .in1(N__18396),
            .in2(_gnd_net_),
            .in3(N__16832),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__20884),
            .ce(N__20651),
            .sr(N__20385));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_9_21_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_9_21_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_9_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_9_21_3  (
            .in0(N__20583),
            .in1(N__18354),
            .in2(_gnd_net_),
            .in3(N__16829),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__20884),
            .ce(N__20651),
            .sr(N__20385));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_9_21_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_9_21_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_9_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_9_21_4  (
            .in0(N__20525),
            .in1(N__18296),
            .in2(_gnd_net_),
            .in3(N__16826),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__20884),
            .ce(N__20651),
            .sr(N__20385));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_9_21_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_9_21_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_9_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_9_21_5  (
            .in0(N__20584),
            .in1(N__18251),
            .in2(_gnd_net_),
            .in3(N__16823),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__20884),
            .ce(N__20651),
            .sr(N__20385));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_9_21_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_9_21_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_9_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_9_21_6  (
            .in0(N__20526),
            .in1(N__19173),
            .in2(_gnd_net_),
            .in3(N__17147),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__20884),
            .ce(N__20651),
            .sr(N__20385));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_9_21_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_9_21_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_9_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_9_21_7  (
            .in0(N__20585),
            .in1(N__19104),
            .in2(_gnd_net_),
            .in3(N__17144),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__20884),
            .ce(N__20651),
            .sr(N__20385));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_9_22_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_9_22_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_9_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_9_22_0  (
            .in0(N__20581),
            .in1(N__19063),
            .in2(_gnd_net_),
            .in3(N__17141),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_9_22_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__20877),
            .ce(N__20659),
            .sr(N__20393));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_9_22_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_9_22_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_9_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_9_22_1  (
            .in0(N__20593),
            .in1(N__19024),
            .in2(_gnd_net_),
            .in3(N__17138),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__20877),
            .ce(N__20659),
            .sr(N__20393));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_9_22_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_9_22_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_9_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_9_22_2  (
            .in0(N__20578),
            .in1(N__18984),
            .in2(_gnd_net_),
            .in3(N__17135),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__20877),
            .ce(N__20659),
            .sr(N__20393));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_9_22_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_9_22_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_9_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_9_22_3  (
            .in0(N__20590),
            .in1(N__18936),
            .in2(_gnd_net_),
            .in3(N__17132),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__20877),
            .ce(N__20659),
            .sr(N__20393));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_9_22_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_9_22_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_9_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_9_22_4  (
            .in0(N__20579),
            .in1(N__18869),
            .in2(_gnd_net_),
            .in3(N__17129),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__20877),
            .ce(N__20659),
            .sr(N__20393));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_9_22_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_9_22_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_9_22_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_9_22_5  (
            .in0(N__20591),
            .in1(N__19475),
            .in2(_gnd_net_),
            .in3(N__17126),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__20877),
            .ce(N__20659),
            .sr(N__20393));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_9_22_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_9_22_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_9_22_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_9_22_6  (
            .in0(N__20580),
            .in1(N__19428),
            .in2(_gnd_net_),
            .in3(N__17123),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__20877),
            .ce(N__20659),
            .sr(N__20393));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_9_22_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_9_22_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_9_22_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_9_22_7  (
            .in0(N__20592),
            .in1(N__19374),
            .in2(_gnd_net_),
            .in3(N__17174),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__20877),
            .ce(N__20659),
            .sr(N__20393));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_9_23_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_9_23_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_9_23_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_9_23_0  (
            .in0(N__20594),
            .in1(N__19327),
            .in2(_gnd_net_),
            .in3(N__17171),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_9_23_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__20872),
            .ce(N__20658),
            .sr(N__20397));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_9_23_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_9_23_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_9_23_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_9_23_1  (
            .in0(N__20586),
            .in1(N__19276),
            .in2(_gnd_net_),
            .in3(N__17168),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__20872),
            .ce(N__20658),
            .sr(N__20397));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_9_23_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_9_23_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_9_23_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_9_23_2  (
            .in0(N__20595),
            .in1(N__19254),
            .in2(_gnd_net_),
            .in3(N__17165),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__20872),
            .ce(N__20658),
            .sr(N__20397));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_9_23_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_9_23_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_9_23_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_9_23_3  (
            .in0(N__20587),
            .in1(N__19230),
            .in2(_gnd_net_),
            .in3(N__17162),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__20872),
            .ce(N__20658),
            .sr(N__20397));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_9_23_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_9_23_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_9_23_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_9_23_4  (
            .in0(N__20596),
            .in1(N__19208),
            .in2(_gnd_net_),
            .in3(N__17159),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__20872),
            .ce(N__20658),
            .sr(N__20397));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_9_23_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_9_23_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_9_23_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_9_23_5  (
            .in0(N__20588),
            .in1(N__19190),
            .in2(_gnd_net_),
            .in3(N__17156),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__20872),
            .ce(N__20658),
            .sr(N__20397));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_9_23_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_9_23_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_9_23_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_9_23_6  (
            .in0(N__20597),
            .in1(N__19734),
            .in2(_gnd_net_),
            .in3(N__17153),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__20872),
            .ce(N__20658),
            .sr(N__20397));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_9_23_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_9_23_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_9_23_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_9_23_7  (
            .in0(N__20589),
            .in1(N__19710),
            .in2(_gnd_net_),
            .in3(N__17150),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__20872),
            .ce(N__20658),
            .sr(N__20397));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_9_24_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_9_24_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_9_24_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_9_24_0  (
            .in0(N__20527),
            .in1(N__19687),
            .in2(_gnd_net_),
            .in3(N__17294),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_9_24_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__20868),
            .ce(N__20663),
            .sr(N__20401));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_9_24_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_9_24_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_9_24_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_9_24_1  (
            .in0(N__20531),
            .in1(N__19666),
            .in2(_gnd_net_),
            .in3(N__17291),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__20868),
            .ce(N__20663),
            .sr(N__20401));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_9_24_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_9_24_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_9_24_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_9_24_2  (
            .in0(N__20528),
            .in1(N__19632),
            .in2(_gnd_net_),
            .in3(N__17288),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__20868),
            .ce(N__20663),
            .sr(N__20401));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_9_24_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_9_24_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_9_24_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_9_24_3  (
            .in0(N__20532),
            .in1(N__19596),
            .in2(_gnd_net_),
            .in3(N__17285),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__20868),
            .ce(N__20663),
            .sr(N__20401));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_9_24_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_9_24_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_9_24_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_9_24_4  (
            .in0(N__20529),
            .in1(N__19646),
            .in2(_gnd_net_),
            .in3(N__17282),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__20868),
            .ce(N__20663),
            .sr(N__20401));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_9_24_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_9_24_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_9_24_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_9_24_5  (
            .in0(N__19610),
            .in1(N__20530),
            .in2(_gnd_net_),
            .in3(N__17279),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20868),
            .ce(N__20663),
            .sr(N__20401));
    defparam \phase_controller_slave.S1_LC_9_30_2 .C_ON=1'b0;
    defparam \phase_controller_slave.S1_LC_9_30_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.S1_LC_9_30_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.S1_LC_9_30_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17276),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20864),
            .ce(),
            .sr(N__20421));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_10_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_10_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_10_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_10_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17237),
            .lcout(\delay_measurement_inst.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20917),
            .ce(N__17195),
            .sr(N__20351));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_10_13_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_10_13_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_10_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_10_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17216),
            .lcout(\delay_measurement_inst.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20917),
            .ce(N__17195),
            .sr(N__20351));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_10_14_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_10_14_1 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_10_14_1  (
            .in0(N__17745),
            .in1(N__17388),
            .in2(N__18616),
            .in3(N__17337),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5OTB1_6_LC_10_14_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5OTB1_6_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5OTB1_6_LC_10_14_2 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5OTB1_6_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(N__18077),
            .in2(N__17570),
            .in3(N__17960),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_10_14_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_10_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_10_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20071),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_10_14_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_10_14_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(N__17428),
            .in2(_gnd_net_),
            .in3(N__17413),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_177_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIF2PP_1_LC_10_15_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIF2PP_1_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIF2PP_1_LC_10_15_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIF2PP_1_LC_10_15_0  (
            .in0(N__18043),
            .in1(N__17395),
            .in2(N__17371),
            .in3(N__17344),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_10_15_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_10_15_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_10_15_1  (
            .in0(N__17324),
            .in1(N__17318),
            .in2(N__17312),
            .in3(N__17303),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC841_7_LC_10_15_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC841_7_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC841_7_LC_10_15_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC841_7_LC_10_15_2  (
            .in0(N__17871),
            .in1(N__17920),
            .in2(N__18056),
            .in3(N__18741),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQMG82_16_LC_10_15_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQMG82_16_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQMG82_16_LC_10_15_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQMG82_16_LC_10_15_3  (
            .in0(N__17788),
            .in1(N__17769),
            .in2(N__17297),
            .in3(N__17809),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKTUL_6_LC_10_15_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKTUL_6_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKTUL_6_LC_10_15_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKTUL_6_LC_10_15_5  (
            .in0(N__17921),
            .in1(N__18089),
            .in2(_gnd_net_),
            .in3(N__17970),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICHJG3_1_LC_10_15_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICHJG3_1_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICHJG3_1_LC_10_15_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICHJG3_1_LC_10_15_6  (
            .in0(N__17810),
            .in1(N__17801),
            .in2(N__17795),
            .in3(N__18005),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_10_15_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_10_15_7 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_10_15_7  (
            .in0(N__17787),
            .in1(N__18612),
            .in2(N__17773),
            .in3(N__17746),
            .lcout(\delay_measurement_inst.N_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_10_16_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_10_16_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_10_16_2  (
            .in0(_gnd_net_),
            .in1(N__17729),
            .in2(_gnd_net_),
            .in3(N__17723),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_10_16_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_10_16_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_10_16_3  (
            .in0(N__17717),
            .in1(N__17696),
            .in2(N__17674),
            .in3(N__17653),
            .lcout(\delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_10_16_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_10_16_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_10_16_5  (
            .in0(N__17636),
            .in1(N__17630),
            .in2(N__17624),
            .in3(N__17615),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_10_16_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_10_16_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_10_16_6  (
            .in0(N__17609),
            .in1(N__17603),
            .in2(N__17597),
            .in3(N__17594),
            .lcout(\delay_measurement_inst.N_35 ),
            .ltout(\delay_measurement_inst.N_35_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_6_LC_10_16_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_6_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_6_LC_10_16_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_6_LC_10_16_7  (
            .in0(N__18122),
            .in1(N__17588),
            .in2(N__17579),
            .in3(N__17576),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_177 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_10_17_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_10_17_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_10_17_0  (
            .in0(N__18578),
            .in1(N__18127),
            .in2(N__18107),
            .in3(N__17940),
            .lcout(\delay_measurement_inst.N_164 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_10_17_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_10_17_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_10_17_1  (
            .in0(N__18748),
            .in1(N__17878),
            .in2(N__18128),
            .in3(N__18575),
            .lcout(\delay_measurement_inst.N_187 ),
            .ltout(\delay_measurement_inst.N_187_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_10_17_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_10_17_2 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_10_17_2  (
            .in0(N__18176),
            .in1(N__18647),
            .in2(N__18167),
            .in3(N__18164),
            .lcout(\delay_measurement_inst.un3_elapsed_time_tr_0_i ),
            .ltout(\delay_measurement_inst.un3_elapsed_time_tr_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_10_17_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_10_17_3 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_10_17_3  (
            .in0(N__20461),
            .in1(_gnd_net_),
            .in2(N__18158),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_10_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_10_17_4 .LUT_INIT=16'b0101000001010001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_10_17_4  (
            .in0(N__18576),
            .in1(N__17939),
            .in2(N__18022),
            .in3(N__18058),
            .lcout(\delay_measurement_inst.N_162_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_10_17_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_10_17_5 .LUT_INIT=16'b0000001000110011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_10_17_5  (
            .in0(N__18126),
            .in1(N__17937),
            .in2(N__18106),
            .in3(N__18057),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_180_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_10_17_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_10_17_6 .LUT_INIT=16'b1111111101010100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_10_17_6  (
            .in0(N__18577),
            .in1(N__18018),
            .in2(N__17984),
            .in3(N__18648),
            .lcout(\delay_measurement_inst.N_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI654I_6_LC_10_17_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI654I_6_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI654I_6_LC_10_17_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI654I_6_LC_10_17_7  (
            .in0(_gnd_net_),
            .in1(N__17977),
            .in2(_gnd_net_),
            .in3(N__17938),
            .lcout(\delay_measurement_inst.delay_tr_reg_5_0_a2_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_10_18_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_10_18_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_10_18_0 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_7_LC_10_18_0  (
            .in0(N__18772),
            .in1(N__18787),
            .in2(N__17849),
            .in3(N__17879),
            .lcout(measured_delay_tr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20892),
            .ce(),
            .sr(N__20366));
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_10_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_10_18_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_10_18_5 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_8_LC_10_18_5  (
            .in0(N__18788),
            .in1(N__18773),
            .in2(N__18721),
            .in3(N__18749),
            .lcout(measured_delay_tr_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20892),
            .ce(),
            .sr(N__20366));
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_10_19_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_10_19_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_10_19_5 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_19_LC_10_19_5  (
            .in0(N__18687),
            .in1(N__18620),
            .in2(_gnd_net_),
            .in3(N__18590),
            .lcout(measured_delay_tr_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20885),
            .ce(N__18506),
            .sr(N__20371));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_10_21_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_10_21_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_10_21_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_10_21_0  (
            .in0(_gnd_net_),
            .in1(N__18484),
            .in2(N__18397),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_10_21_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__20873),
            .ce(N__19495),
            .sr(N__20375));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_10_21_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_10_21_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_10_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_10_21_1  (
            .in0(_gnd_net_),
            .in1(N__18442),
            .in2(N__18355),
            .in3(N__18401),
            .lcout(\delay_measurement_inst.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__20873),
            .ce(N__19495),
            .sr(N__20375));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_10_21_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_10_21_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_10_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_10_21_2  (
            .in0(_gnd_net_),
            .in1(N__18294),
            .in2(N__18398),
            .in3(N__18359),
            .lcout(\delay_measurement_inst.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__20873),
            .ce(N__19495),
            .sr(N__20375));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_10_21_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_10_21_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_10_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_10_21_3  (
            .in0(_gnd_net_),
            .in1(N__18249),
            .in2(N__18356),
            .in3(N__18299),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__20873),
            .ce(N__19495),
            .sr(N__20375));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_10_21_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_10_21_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_10_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_10_21_4  (
            .in0(_gnd_net_),
            .in1(N__18295),
            .in2(N__19174),
            .in3(N__18254),
            .lcout(\delay_measurement_inst.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__20873),
            .ce(N__19495),
            .sr(N__20375));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_10_21_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_10_21_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_10_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_10_21_5  (
            .in0(_gnd_net_),
            .in1(N__18250),
            .in2(N__19105),
            .in3(N__18206),
            .lcout(\delay_measurement_inst.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__20873),
            .ce(N__19495),
            .sr(N__20375));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_10_21_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_10_21_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_10_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_10_21_6  (
            .in0(_gnd_net_),
            .in1(N__19062),
            .in2(N__19175),
            .in3(N__19109),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__20873),
            .ce(N__19495),
            .sr(N__20375));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_10_21_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_10_21_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_10_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_10_21_7  (
            .in0(_gnd_net_),
            .in1(N__19023),
            .in2(N__19106),
            .in3(N__19067),
            .lcout(\delay_measurement_inst.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__20873),
            .ce(N__19495),
            .sr(N__20375));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_10_22_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_10_22_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_10_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_10_22_0  (
            .in0(_gnd_net_),
            .in1(N__19064),
            .in2(N__18985),
            .in3(N__19028),
            .lcout(\delay_measurement_inst.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_10_22_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__20869),
            .ce(N__19494),
            .sr(N__20381));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_10_22_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_10_22_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_10_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_10_22_1  (
            .in0(_gnd_net_),
            .in1(N__19025),
            .in2(N__18937),
            .in3(N__18989),
            .lcout(\delay_measurement_inst.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__20869),
            .ce(N__19494),
            .sr(N__20381));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_10_22_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_10_22_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_10_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_10_22_2  (
            .in0(_gnd_net_),
            .in1(N__18867),
            .in2(N__18986),
            .in3(N__18941),
            .lcout(\delay_measurement_inst.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__20869),
            .ce(N__19494),
            .sr(N__20381));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_10_22_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_10_22_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_10_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_10_22_3  (
            .in0(_gnd_net_),
            .in1(N__19473),
            .in2(N__18938),
            .in3(N__18872),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__20869),
            .ce(N__19494),
            .sr(N__20381));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_10_22_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_10_22_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_10_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_10_22_4  (
            .in0(_gnd_net_),
            .in1(N__18868),
            .in2(N__19429),
            .in3(N__18791),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__20869),
            .ce(N__19494),
            .sr(N__20381));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_10_22_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_10_22_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_10_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_10_22_5  (
            .in0(_gnd_net_),
            .in1(N__19474),
            .in2(N__19375),
            .in3(N__19433),
            .lcout(\delay_measurement_inst.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__20869),
            .ce(N__19494),
            .sr(N__20381));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_10_22_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_10_22_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_10_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_10_22_6  (
            .in0(_gnd_net_),
            .in1(N__19326),
            .in2(N__19430),
            .in3(N__19379),
            .lcout(\delay_measurement_inst.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__20869),
            .ce(N__19494),
            .sr(N__20381));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_10_22_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_10_22_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_10_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_10_22_7  (
            .in0(_gnd_net_),
            .in1(N__19275),
            .in2(N__19376),
            .in3(N__19331),
            .lcout(\delay_measurement_inst.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__20869),
            .ce(N__19494),
            .sr(N__20381));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_10_23_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_10_23_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_10_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_10_23_0  (
            .in0(_gnd_net_),
            .in1(N__19328),
            .in2(N__19255),
            .in3(N__19280),
            .lcout(\delay_measurement_inst.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_10_23_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__20867),
            .ce(N__19493),
            .sr(N__20389));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_10_23_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_10_23_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_10_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_10_23_1  (
            .in0(_gnd_net_),
            .in1(N__19277),
            .in2(N__19231),
            .in3(N__19259),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__20867),
            .ce(N__19493),
            .sr(N__20389));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_10_23_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_10_23_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_10_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_10_23_2  (
            .in0(_gnd_net_),
            .in1(N__19206),
            .in2(N__19256),
            .in3(N__19235),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__20867),
            .ce(N__19493),
            .sr(N__20389));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_10_23_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_10_23_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_10_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_10_23_3  (
            .in0(_gnd_net_),
            .in1(N__19188),
            .in2(N__19232),
            .in3(N__19211),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__20867),
            .ce(N__19493),
            .sr(N__20389));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_10_23_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_10_23_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_10_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_10_23_4  (
            .in0(_gnd_net_),
            .in1(N__19207),
            .in2(N__19735),
            .in3(N__19193),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__20867),
            .ce(N__19493),
            .sr(N__20389));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_10_23_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_10_23_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_10_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_10_23_5  (
            .in0(_gnd_net_),
            .in1(N__19189),
            .in2(N__19711),
            .in3(N__19739),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__20867),
            .ce(N__19493),
            .sr(N__20389));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_10_23_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_10_23_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_10_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_10_23_6  (
            .in0(_gnd_net_),
            .in1(N__19686),
            .in2(N__19736),
            .in3(N__19715),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__20867),
            .ce(N__19493),
            .sr(N__20389));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_10_23_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_10_23_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_10_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_10_23_7  (
            .in0(_gnd_net_),
            .in1(N__19665),
            .in2(N__19712),
            .in3(N__19691),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__20867),
            .ce(N__19493),
            .sr(N__20389));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_10_24_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_10_24_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_10_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_10_24_0  (
            .in0(_gnd_net_),
            .in1(N__19688),
            .in2(N__19633),
            .in3(N__19670),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_10_24_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__20865),
            .ce(N__19492),
            .sr(N__20394));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_10_24_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_10_24_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_10_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_10_24_1  (
            .in0(_gnd_net_),
            .in1(N__19667),
            .in2(N__19597),
            .in3(N__19649),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__20865),
            .ce(N__19492),
            .sr(N__20394));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_10_24_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_10_24_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_10_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_10_24_2  (
            .in0(_gnd_net_),
            .in1(N__19645),
            .in2(N__19634),
            .in3(N__19613),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__20865),
            .ce(N__19492),
            .sr(N__20394));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_10_24_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_10_24_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_10_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_10_24_3  (
            .in0(_gnd_net_),
            .in1(N__19609),
            .in2(N__19598),
            .in3(N__19577),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__20865),
            .ce(N__19492),
            .sr(N__20394));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_10_24_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_10_24_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_10_24_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_10_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19574),
            .lcout(\delay_measurement_inst.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20865),
            .ce(N__19492),
            .sr(N__20394));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_11_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_11_13_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_11_13_5 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_11_13_5  (
            .in0(N__20102),
            .in1(N__20090),
            .in2(_gnd_net_),
            .in3(N__20072),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20911),
            .ce(),
            .sr(N__20350));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_11_14_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_11_14_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(N__20089),
            .in2(_gnd_net_),
            .in3(N__20069),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_255_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.S2_LC_11_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_11_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_11_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_11_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19919),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20878),
            .ce(),
            .sr(N__20367));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_11_23_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_11_23_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_11_23_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_11_23_1  (
            .in0(N__19865),
            .in1(N__19859),
            .in2(N__19853),
            .in3(N__19844),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_7_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_11_23_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_11_23_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_11_23_2  (
            .in0(N__19838),
            .in1(N__19763),
            .in2(N__19832),
            .in3(N__19745),
            .lcout(\delay_measurement_inst.N_276 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_11_23_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_11_23_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_11_23_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_11_23_3  (
            .in0(N__19790),
            .in1(N__19784),
            .in2(N__19778),
            .in3(N__19769),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_6_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI23AG_29_LC_11_24_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI23AG_29_LC_11_24_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI23AG_29_LC_11_24_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI23AG_29_LC_11_24_0  (
            .in0(_gnd_net_),
            .in1(N__19757),
            .in2(_gnd_net_),
            .in3(N__19751),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_tr_LC_12_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_12_12_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.start_timer_tr_LC_12_12_2 .LUT_INIT=16'b1010101001100110;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_12_12_2  (
            .in0(N__19973),
            .in1(N__20009),
            .in2(_gnd_net_),
            .in3(N__19989),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20910),
            .ce(),
            .sr(N__20346));
    defparam \delay_measurement_inst.prev_tr_sig_LC_12_12_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.prev_tr_sig_LC_12_12_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.prev_tr_sig_LC_12_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.prev_tr_sig_LC_12_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20010),
            .lcout(\delay_measurement_inst.prev_tr_sigZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20910),
            .ce(),
            .sr(N__20346));
    defparam \delay_measurement_inst.stop_timer_tr_LC_12_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_12_13_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.stop_timer_tr_LC_12_13_3 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_12_13_3  (
            .in0(N__20012),
            .in1(N__19972),
            .in2(N__20467),
            .in3(N__19990),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20906),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_12_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_12_13_5 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_12_13_5  (
            .in0(N__20101),
            .in1(N__20088),
            .in2(_gnd_net_),
            .in3(N__20070),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_256_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_TR2_LC_13_12_1.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_TR2_LC_13_12_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_TR2_LC_13_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_TR2_LC_13_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20018),
            .lcout(delay_tr_d2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20918),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_TR1_LC_13_12_5.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_TR1_LC_13_12_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_TR1_LC_13_12_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_DELAY_TR1_LC_13_12_5 (
            .in0(N__20036),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(delay_tr_d1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20918),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.tr_state_0_LC_13_13_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.tr_state_0_LC_13_13_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.tr_state_0_LC_13_13_6 .LUT_INIT=16'b1100110001100110;
    LogicCell40 \delay_measurement_inst.tr_state_0_LC_13_13_6  (
            .in0(N__20011),
            .in1(N__19971),
            .in2(_gnd_net_),
            .in3(N__19991),
            .lcout(\delay_measurement_inst.tr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20912),
            .ce(N__20188),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_HC2_LC_13_17_3.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_HC2_LC_13_17_3.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_HC2_LC_13_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_HC2_LC_13_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19940),
            .lcout(delay_hc_d2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20893),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_HC1_LC_13_17_6.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_HC1_LC_13_17_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_HC1_LC_13_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_HC1_LC_13_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19955),
            .lcout(delay_hc_d1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20893),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.hc_state_0_LC_13_18_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.hc_state_0_LC_13_18_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.hc_state_0_LC_13_18_3 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \delay_measurement_inst.hc_state_0_LC_13_18_3  (
            .in0(N__21008),
            .in1(N__20982),
            .in2(_gnd_net_),
            .in3(N__20955),
            .lcout(\delay_measurement_inst.hc_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20886),
            .ce(N__20171),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_hc_LC_13_19_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_13_19_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.stop_timer_hc_LC_13_19_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_13_19_5  (
            .in0(N__21004),
            .in1(N__20983),
            .in2(N__20468),
            .in3(N__20964),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20879),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.prev_hc_sig_LC_13_20_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.prev_hc_sig_LC_13_20_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.prev_hc_sig_LC_13_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.prev_hc_sig_LC_13_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20966),
            .lcout(\delay_measurement_inst.prev_hc_sigZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20874),
            .ce(),
            .sr(N__20360));
    defparam \delay_measurement_inst.start_timer_hc_LC_13_20_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_13_20_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.start_timer_hc_LC_13_20_2 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_13_20_2  (
            .in0(N__21003),
            .in1(N__20987),
            .in2(_gnd_net_),
            .in3(N__20965),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20874),
            .ce(),
            .sr(N__20360));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_13_20_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_13_20_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_13_20_5 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_13_20_5  (
            .in0(N__20679),
            .in1(N__20693),
            .in2(_gnd_net_),
            .in3(N__20615),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20874),
            .ce(),
            .sr(N__20360));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_21_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_21_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_21_2  (
            .in0(_gnd_net_),
            .in1(N__20680),
            .in2(_gnd_net_),
            .in3(N__20612),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_253_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_13_21_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_13_21_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_13_21_6 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_13_21_6  (
            .in0(N__20692),
            .in1(N__20681),
            .in2(_gnd_net_),
            .in3(N__20614),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_254_i_g ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_13_21_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_13_21_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_13_21_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_13_21_7  (
            .in0(N__20613),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam reset_ibuf_gb_io_RNI79U7_LC_13_25_4.C_ON=1'b0;
    defparam reset_ibuf_gb_io_RNI79U7_LC_13_25_4.SEQ_MODE=4'b0000;
    defparam reset_ibuf_gb_io_RNI79U7_LC_13_25_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 reset_ibuf_gb_io_RNI79U7_LC_13_25_4 (
            .in0(N__20462),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(red_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // MAIN
