// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Apr 4 2025 00:09:05

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    start_stop,
    s2_phy,
    T23,
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    T45,
    T12,
    s4_phy,
    rgb_g,
    T01,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    input start_stop;
    output s2_phy;
    output T23;
    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output T45;
    output T12;
    output s4_phy;
    output rgb_g;
    output T01;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__48428;
    wire N__48427;
    wire N__48426;
    wire N__48417;
    wire N__48416;
    wire N__48415;
    wire N__48408;
    wire N__48407;
    wire N__48406;
    wire N__48399;
    wire N__48398;
    wire N__48397;
    wire N__48390;
    wire N__48389;
    wire N__48388;
    wire N__48381;
    wire N__48380;
    wire N__48379;
    wire N__48372;
    wire N__48371;
    wire N__48370;
    wire N__48363;
    wire N__48362;
    wire N__48361;
    wire N__48354;
    wire N__48353;
    wire N__48352;
    wire N__48345;
    wire N__48344;
    wire N__48343;
    wire N__48336;
    wire N__48335;
    wire N__48334;
    wire N__48327;
    wire N__48326;
    wire N__48325;
    wire N__48318;
    wire N__48317;
    wire N__48316;
    wire N__48309;
    wire N__48308;
    wire N__48307;
    wire N__48300;
    wire N__48299;
    wire N__48298;
    wire N__48291;
    wire N__48290;
    wire N__48289;
    wire N__48282;
    wire N__48281;
    wire N__48280;
    wire N__48263;
    wire N__48262;
    wire N__48257;
    wire N__48256;
    wire N__48253;
    wire N__48250;
    wire N__48247;
    wire N__48242;
    wire N__48239;
    wire N__48238;
    wire N__48237;
    wire N__48234;
    wire N__48231;
    wire N__48228;
    wire N__48225;
    wire N__48220;
    wire N__48219;
    wire N__48214;
    wire N__48211;
    wire N__48206;
    wire N__48203;
    wire N__48202;
    wire N__48199;
    wire N__48196;
    wire N__48193;
    wire N__48190;
    wire N__48189;
    wire N__48186;
    wire N__48183;
    wire N__48180;
    wire N__48177;
    wire N__48174;
    wire N__48167;
    wire N__48166;
    wire N__48163;
    wire N__48160;
    wire N__48159;
    wire N__48156;
    wire N__48153;
    wire N__48150;
    wire N__48147;
    wire N__48144;
    wire N__48141;
    wire N__48140;
    wire N__48133;
    wire N__48130;
    wire N__48125;
    wire N__48122;
    wire N__48121;
    wire N__48118;
    wire N__48115;
    wire N__48112;
    wire N__48109;
    wire N__48108;
    wire N__48105;
    wire N__48102;
    wire N__48099;
    wire N__48096;
    wire N__48093;
    wire N__48086;
    wire N__48085;
    wire N__48084;
    wire N__48079;
    wire N__48076;
    wire N__48073;
    wire N__48070;
    wire N__48067;
    wire N__48066;
    wire N__48063;
    wire N__48060;
    wire N__48057;
    wire N__48050;
    wire N__48047;
    wire N__48044;
    wire N__48043;
    wire N__48040;
    wire N__48037;
    wire N__48034;
    wire N__48029;
    wire N__48026;
    wire N__48025;
    wire N__48024;
    wire N__48021;
    wire N__48018;
    wire N__48015;
    wire N__48010;
    wire N__48005;
    wire N__48002;
    wire N__48001;
    wire N__47998;
    wire N__47995;
    wire N__47992;
    wire N__47991;
    wire N__47988;
    wire N__47985;
    wire N__47982;
    wire N__47981;
    wire N__47978;
    wire N__47973;
    wire N__47970;
    wire N__47963;
    wire N__47960;
    wire N__47957;
    wire N__47956;
    wire N__47953;
    wire N__47950;
    wire N__47947;
    wire N__47942;
    wire N__47939;
    wire N__47938;
    wire N__47935;
    wire N__47932;
    wire N__47931;
    wire N__47926;
    wire N__47923;
    wire N__47920;
    wire N__47915;
    wire N__47914;
    wire N__47911;
    wire N__47908;
    wire N__47907;
    wire N__47904;
    wire N__47901;
    wire N__47898;
    wire N__47897;
    wire N__47894;
    wire N__47889;
    wire N__47886;
    wire N__47879;
    wire N__47876;
    wire N__47875;
    wire N__47874;
    wire N__47873;
    wire N__47872;
    wire N__47871;
    wire N__47870;
    wire N__47869;
    wire N__47868;
    wire N__47867;
    wire N__47866;
    wire N__47865;
    wire N__47864;
    wire N__47863;
    wire N__47862;
    wire N__47861;
    wire N__47860;
    wire N__47859;
    wire N__47858;
    wire N__47857;
    wire N__47856;
    wire N__47855;
    wire N__47854;
    wire N__47853;
    wire N__47852;
    wire N__47851;
    wire N__47850;
    wire N__47849;
    wire N__47848;
    wire N__47847;
    wire N__47846;
    wire N__47845;
    wire N__47844;
    wire N__47843;
    wire N__47842;
    wire N__47841;
    wire N__47840;
    wire N__47839;
    wire N__47838;
    wire N__47837;
    wire N__47836;
    wire N__47835;
    wire N__47834;
    wire N__47833;
    wire N__47832;
    wire N__47831;
    wire N__47830;
    wire N__47829;
    wire N__47828;
    wire N__47827;
    wire N__47826;
    wire N__47825;
    wire N__47824;
    wire N__47823;
    wire N__47822;
    wire N__47821;
    wire N__47820;
    wire N__47819;
    wire N__47818;
    wire N__47817;
    wire N__47816;
    wire N__47815;
    wire N__47814;
    wire N__47813;
    wire N__47812;
    wire N__47811;
    wire N__47810;
    wire N__47809;
    wire N__47808;
    wire N__47807;
    wire N__47806;
    wire N__47805;
    wire N__47804;
    wire N__47803;
    wire N__47802;
    wire N__47801;
    wire N__47800;
    wire N__47799;
    wire N__47798;
    wire N__47797;
    wire N__47796;
    wire N__47795;
    wire N__47794;
    wire N__47793;
    wire N__47792;
    wire N__47791;
    wire N__47790;
    wire N__47789;
    wire N__47788;
    wire N__47787;
    wire N__47786;
    wire N__47785;
    wire N__47784;
    wire N__47783;
    wire N__47782;
    wire N__47781;
    wire N__47780;
    wire N__47779;
    wire N__47778;
    wire N__47777;
    wire N__47776;
    wire N__47775;
    wire N__47774;
    wire N__47773;
    wire N__47772;
    wire N__47771;
    wire N__47770;
    wire N__47769;
    wire N__47768;
    wire N__47767;
    wire N__47766;
    wire N__47765;
    wire N__47764;
    wire N__47763;
    wire N__47762;
    wire N__47761;
    wire N__47760;
    wire N__47759;
    wire N__47758;
    wire N__47519;
    wire N__47516;
    wire N__47515;
    wire N__47514;
    wire N__47513;
    wire N__47512;
    wire N__47511;
    wire N__47510;
    wire N__47509;
    wire N__47508;
    wire N__47489;
    wire N__47486;
    wire N__47483;
    wire N__47482;
    wire N__47481;
    wire N__47480;
    wire N__47479;
    wire N__47478;
    wire N__47477;
    wire N__47476;
    wire N__47475;
    wire N__47474;
    wire N__47473;
    wire N__47472;
    wire N__47471;
    wire N__47470;
    wire N__47469;
    wire N__47466;
    wire N__47463;
    wire N__47460;
    wire N__47457;
    wire N__47454;
    wire N__47449;
    wire N__47444;
    wire N__47439;
    wire N__47434;
    wire N__47431;
    wire N__47428;
    wire N__47425;
    wire N__47422;
    wire N__47419;
    wire N__47418;
    wire N__47417;
    wire N__47416;
    wire N__47415;
    wire N__47414;
    wire N__47411;
    wire N__47410;
    wire N__47409;
    wire N__47408;
    wire N__47407;
    wire N__47406;
    wire N__47405;
    wire N__47404;
    wire N__47403;
    wire N__47402;
    wire N__47401;
    wire N__47400;
    wire N__47399;
    wire N__47398;
    wire N__47397;
    wire N__47396;
    wire N__47395;
    wire N__47394;
    wire N__47393;
    wire N__47392;
    wire N__47391;
    wire N__47390;
    wire N__47389;
    wire N__47388;
    wire N__47387;
    wire N__47386;
    wire N__47385;
    wire N__47384;
    wire N__47383;
    wire N__47382;
    wire N__47381;
    wire N__47380;
    wire N__47379;
    wire N__47378;
    wire N__47377;
    wire N__47376;
    wire N__47375;
    wire N__47374;
    wire N__47373;
    wire N__47372;
    wire N__47371;
    wire N__47370;
    wire N__47369;
    wire N__47368;
    wire N__47367;
    wire N__47366;
    wire N__47365;
    wire N__47364;
    wire N__47363;
    wire N__47362;
    wire N__47361;
    wire N__47360;
    wire N__47359;
    wire N__47358;
    wire N__47355;
    wire N__47354;
    wire N__47353;
    wire N__47352;
    wire N__47351;
    wire N__47350;
    wire N__47349;
    wire N__47346;
    wire N__47343;
    wire N__47342;
    wire N__47341;
    wire N__47340;
    wire N__47339;
    wire N__47336;
    wire N__47335;
    wire N__47334;
    wire N__47333;
    wire N__47332;
    wire N__47331;
    wire N__47330;
    wire N__47329;
    wire N__47328;
    wire N__47327;
    wire N__47326;
    wire N__47325;
    wire N__47324;
    wire N__47323;
    wire N__47322;
    wire N__47321;
    wire N__47320;
    wire N__47319;
    wire N__47318;
    wire N__47317;
    wire N__47316;
    wire N__47315;
    wire N__47314;
    wire N__47313;
    wire N__47312;
    wire N__47311;
    wire N__47308;
    wire N__47307;
    wire N__47306;
    wire N__47305;
    wire N__47304;
    wire N__47303;
    wire N__47302;
    wire N__47301;
    wire N__47300;
    wire N__47299;
    wire N__47296;
    wire N__47295;
    wire N__47294;
    wire N__47293;
    wire N__47290;
    wire N__47289;
    wire N__47288;
    wire N__47287;
    wire N__47286;
    wire N__47285;
    wire N__47284;
    wire N__47283;
    wire N__47282;
    wire N__47281;
    wire N__47030;
    wire N__47027;
    wire N__47024;
    wire N__47021;
    wire N__47020;
    wire N__47019;
    wire N__47016;
    wire N__47013;
    wire N__47010;
    wire N__47007;
    wire N__47004;
    wire N__47001;
    wire N__46998;
    wire N__46995;
    wire N__46992;
    wire N__46987;
    wire N__46982;
    wire N__46981;
    wire N__46978;
    wire N__46975;
    wire N__46972;
    wire N__46969;
    wire N__46968;
    wire N__46965;
    wire N__46962;
    wire N__46959;
    wire N__46956;
    wire N__46953;
    wire N__46946;
    wire N__46945;
    wire N__46942;
    wire N__46939;
    wire N__46936;
    wire N__46935;
    wire N__46930;
    wire N__46929;
    wire N__46926;
    wire N__46923;
    wire N__46920;
    wire N__46913;
    wire N__46910;
    wire N__46909;
    wire N__46906;
    wire N__46903;
    wire N__46900;
    wire N__46897;
    wire N__46896;
    wire N__46893;
    wire N__46890;
    wire N__46887;
    wire N__46884;
    wire N__46881;
    wire N__46874;
    wire N__46873;
    wire N__46872;
    wire N__46869;
    wire N__46864;
    wire N__46859;
    wire N__46858;
    wire N__46855;
    wire N__46852;
    wire N__46847;
    wire N__46844;
    wire N__46841;
    wire N__46840;
    wire N__46839;
    wire N__46836;
    wire N__46833;
    wire N__46830;
    wire N__46825;
    wire N__46820;
    wire N__46817;
    wire N__46814;
    wire N__46813;
    wire N__46812;
    wire N__46809;
    wire N__46806;
    wire N__46805;
    wire N__46802;
    wire N__46797;
    wire N__46794;
    wire N__46791;
    wire N__46788;
    wire N__46785;
    wire N__46782;
    wire N__46775;
    wire N__46772;
    wire N__46771;
    wire N__46766;
    wire N__46765;
    wire N__46762;
    wire N__46759;
    wire N__46756;
    wire N__46751;
    wire N__46750;
    wire N__46749;
    wire N__46742;
    wire N__46739;
    wire N__46736;
    wire N__46735;
    wire N__46732;
    wire N__46729;
    wire N__46724;
    wire N__46721;
    wire N__46718;
    wire N__46717;
    wire N__46714;
    wire N__46711;
    wire N__46710;
    wire N__46705;
    wire N__46702;
    wire N__46699;
    wire N__46694;
    wire N__46693;
    wire N__46692;
    wire N__46689;
    wire N__46686;
    wire N__46683;
    wire N__46682;
    wire N__46677;
    wire N__46674;
    wire N__46671;
    wire N__46668;
    wire N__46663;
    wire N__46658;
    wire N__46655;
    wire N__46654;
    wire N__46651;
    wire N__46648;
    wire N__46643;
    wire N__46642;
    wire N__46639;
    wire N__46636;
    wire N__46633;
    wire N__46628;
    wire N__46627;
    wire N__46624;
    wire N__46621;
    wire N__46620;
    wire N__46617;
    wire N__46612;
    wire N__46609;
    wire N__46606;
    wire N__46605;
    wire N__46602;
    wire N__46599;
    wire N__46596;
    wire N__46589;
    wire N__46586;
    wire N__46585;
    wire N__46580;
    wire N__46579;
    wire N__46576;
    wire N__46573;
    wire N__46570;
    wire N__46565;
    wire N__46562;
    wire N__46559;
    wire N__46558;
    wire N__46557;
    wire N__46554;
    wire N__46551;
    wire N__46548;
    wire N__46543;
    wire N__46542;
    wire N__46539;
    wire N__46536;
    wire N__46533;
    wire N__46526;
    wire N__46523;
    wire N__46520;
    wire N__46519;
    wire N__46516;
    wire N__46513;
    wire N__46512;
    wire N__46509;
    wire N__46506;
    wire N__46503;
    wire N__46500;
    wire N__46497;
    wire N__46490;
    wire N__46487;
    wire N__46484;
    wire N__46483;
    wire N__46482;
    wire N__46479;
    wire N__46474;
    wire N__46473;
    wire N__46468;
    wire N__46465;
    wire N__46460;
    wire N__46457;
    wire N__46454;
    wire N__46453;
    wire N__46450;
    wire N__46447;
    wire N__46446;
    wire N__46443;
    wire N__46440;
    wire N__46437;
    wire N__46434;
    wire N__46431;
    wire N__46424;
    wire N__46423;
    wire N__46420;
    wire N__46419;
    wire N__46416;
    wire N__46413;
    wire N__46412;
    wire N__46409;
    wire N__46404;
    wire N__46401;
    wire N__46398;
    wire N__46391;
    wire N__46388;
    wire N__46385;
    wire N__46384;
    wire N__46383;
    wire N__46380;
    wire N__46377;
    wire N__46374;
    wire N__46369;
    wire N__46364;
    wire N__46361;
    wire N__46358;
    wire N__46355;
    wire N__46352;
    wire N__46351;
    wire N__46348;
    wire N__46345;
    wire N__46344;
    wire N__46343;
    wire N__46340;
    wire N__46337;
    wire N__46334;
    wire N__46331;
    wire N__46322;
    wire N__46319;
    wire N__46318;
    wire N__46313;
    wire N__46312;
    wire N__46309;
    wire N__46306;
    wire N__46303;
    wire N__46298;
    wire N__46295;
    wire N__46294;
    wire N__46293;
    wire N__46292;
    wire N__46289;
    wire N__46284;
    wire N__46281;
    wire N__46276;
    wire N__46271;
    wire N__46268;
    wire N__46265;
    wire N__46264;
    wire N__46261;
    wire N__46258;
    wire N__46257;
    wire N__46252;
    wire N__46249;
    wire N__46246;
    wire N__46241;
    wire N__46238;
    wire N__46235;
    wire N__46234;
    wire N__46231;
    wire N__46228;
    wire N__46227;
    wire N__46222;
    wire N__46219;
    wire N__46216;
    wire N__46215;
    wire N__46212;
    wire N__46209;
    wire N__46206;
    wire N__46199;
    wire N__46196;
    wire N__46195;
    wire N__46192;
    wire N__46189;
    wire N__46184;
    wire N__46183;
    wire N__46180;
    wire N__46177;
    wire N__46174;
    wire N__46169;
    wire N__46166;
    wire N__46165;
    wire N__46164;
    wire N__46161;
    wire N__46158;
    wire N__46155;
    wire N__46154;
    wire N__46151;
    wire N__46146;
    wire N__46143;
    wire N__46136;
    wire N__46133;
    wire N__46132;
    wire N__46127;
    wire N__46126;
    wire N__46123;
    wire N__46120;
    wire N__46117;
    wire N__46112;
    wire N__46111;
    wire N__46110;
    wire N__46107;
    wire N__46102;
    wire N__46099;
    wire N__46096;
    wire N__46095;
    wire N__46092;
    wire N__46089;
    wire N__46086;
    wire N__46079;
    wire N__46076;
    wire N__46075;
    wire N__46070;
    wire N__46069;
    wire N__46066;
    wire N__46063;
    wire N__46060;
    wire N__46055;
    wire N__46054;
    wire N__46051;
    wire N__46050;
    wire N__46047;
    wire N__46046;
    wire N__46043;
    wire N__46040;
    wire N__46037;
    wire N__46034;
    wire N__46029;
    wire N__46022;
    wire N__46019;
    wire N__46018;
    wire N__46015;
    wire N__46012;
    wire N__46009;
    wire N__46008;
    wire N__46005;
    wire N__46002;
    wire N__45999;
    wire N__45996;
    wire N__45989;
    wire N__45986;
    wire N__45985;
    wire N__45984;
    wire N__45979;
    wire N__45976;
    wire N__45975;
    wire N__45972;
    wire N__45969;
    wire N__45966;
    wire N__45963;
    wire N__45960;
    wire N__45957;
    wire N__45950;
    wire N__45947;
    wire N__45946;
    wire N__45943;
    wire N__45940;
    wire N__45937;
    wire N__45936;
    wire N__45933;
    wire N__45930;
    wire N__45927;
    wire N__45924;
    wire N__45917;
    wire N__45916;
    wire N__45915;
    wire N__45912;
    wire N__45909;
    wire N__45906;
    wire N__45903;
    wire N__45900;
    wire N__45899;
    wire N__45894;
    wire N__45891;
    wire N__45888;
    wire N__45885;
    wire N__45882;
    wire N__45879;
    wire N__45872;
    wire N__45869;
    wire N__45868;
    wire N__45865;
    wire N__45862;
    wire N__45861;
    wire N__45856;
    wire N__45853;
    wire N__45850;
    wire N__45845;
    wire N__45842;
    wire N__45839;
    wire N__45838;
    wire N__45837;
    wire N__45836;
    wire N__45833;
    wire N__45830;
    wire N__45827;
    wire N__45824;
    wire N__45821;
    wire N__45818;
    wire N__45813;
    wire N__45810;
    wire N__45807;
    wire N__45804;
    wire N__45797;
    wire N__45794;
    wire N__45793;
    wire N__45790;
    wire N__45787;
    wire N__45782;
    wire N__45781;
    wire N__45778;
    wire N__45775;
    wire N__45772;
    wire N__45767;
    wire N__45764;
    wire N__45763;
    wire N__45758;
    wire N__45757;
    wire N__45756;
    wire N__45753;
    wire N__45750;
    wire N__45747;
    wire N__45744;
    wire N__45741;
    wire N__45738;
    wire N__45735;
    wire N__45732;
    wire N__45729;
    wire N__45722;
    wire N__45719;
    wire N__45716;
    wire N__45715;
    wire N__45712;
    wire N__45709;
    wire N__45708;
    wire N__45703;
    wire N__45700;
    wire N__45697;
    wire N__45692;
    wire N__45691;
    wire N__45688;
    wire N__45683;
    wire N__45682;
    wire N__45679;
    wire N__45676;
    wire N__45673;
    wire N__45670;
    wire N__45669;
    wire N__45666;
    wire N__45663;
    wire N__45660;
    wire N__45653;
    wire N__45650;
    wire N__45647;
    wire N__45646;
    wire N__45643;
    wire N__45640;
    wire N__45639;
    wire N__45634;
    wire N__45631;
    wire N__45628;
    wire N__45623;
    wire N__45622;
    wire N__45619;
    wire N__45616;
    wire N__45611;
    wire N__45610;
    wire N__45607;
    wire N__45604;
    wire N__45603;
    wire N__45600;
    wire N__45597;
    wire N__45594;
    wire N__45591;
    wire N__45588;
    wire N__45585;
    wire N__45578;
    wire N__45575;
    wire N__45572;
    wire N__45571;
    wire N__45568;
    wire N__45565;
    wire N__45564;
    wire N__45559;
    wire N__45556;
    wire N__45553;
    wire N__45548;
    wire N__45545;
    wire N__45544;
    wire N__45543;
    wire N__45540;
    wire N__45535;
    wire N__45530;
    wire N__45529;
    wire N__45526;
    wire N__45523;
    wire N__45518;
    wire N__45515;
    wire N__45512;
    wire N__45511;
    wire N__45508;
    wire N__45505;
    wire N__45504;
    wire N__45499;
    wire N__45496;
    wire N__45493;
    wire N__45488;
    wire N__45485;
    wire N__45482;
    wire N__45479;
    wire N__45478;
    wire N__45477;
    wire N__45474;
    wire N__45471;
    wire N__45470;
    wire N__45467;
    wire N__45464;
    wire N__45461;
    wire N__45458;
    wire N__45449;
    wire N__45446;
    wire N__45443;
    wire N__45440;
    wire N__45437;
    wire N__45434;
    wire N__45431;
    wire N__45428;
    wire N__45425;
    wire N__45424;
    wire N__45421;
    wire N__45418;
    wire N__45417;
    wire N__45414;
    wire N__45411;
    wire N__45408;
    wire N__45401;
    wire N__45398;
    wire N__45395;
    wire N__45392;
    wire N__45389;
    wire N__45386;
    wire N__45383;
    wire N__45380;
    wire N__45377;
    wire N__45374;
    wire N__45371;
    wire N__45368;
    wire N__45367;
    wire N__45366;
    wire N__45363;
    wire N__45360;
    wire N__45357;
    wire N__45354;
    wire N__45347;
    wire N__45344;
    wire N__45341;
    wire N__45338;
    wire N__45335;
    wire N__45332;
    wire N__45329;
    wire N__45326;
    wire N__45323;
    wire N__45320;
    wire N__45317;
    wire N__45316;
    wire N__45315;
    wire N__45312;
    wire N__45309;
    wire N__45306;
    wire N__45303;
    wire N__45300;
    wire N__45293;
    wire N__45292;
    wire N__45291;
    wire N__45290;
    wire N__45289;
    wire N__45288;
    wire N__45287;
    wire N__45284;
    wire N__45281;
    wire N__45280;
    wire N__45279;
    wire N__45278;
    wire N__45275;
    wire N__45272;
    wire N__45271;
    wire N__45268;
    wire N__45267;
    wire N__45266;
    wire N__45265;
    wire N__45264;
    wire N__45263;
    wire N__45260;
    wire N__45259;
    wire N__45258;
    wire N__45257;
    wire N__45254;
    wire N__45253;
    wire N__45248;
    wire N__45245;
    wire N__45242;
    wire N__45241;
    wire N__45238;
    wire N__45237;
    wire N__45236;
    wire N__45235;
    wire N__45234;
    wire N__45233;
    wire N__45232;
    wire N__45227;
    wire N__45216;
    wire N__45215;
    wire N__45212;
    wire N__45211;
    wire N__45210;
    wire N__45209;
    wire N__45208;
    wire N__45207;
    wire N__45206;
    wire N__45203;
    wire N__45202;
    wire N__45201;
    wire N__45200;
    wire N__45199;
    wire N__45198;
    wire N__45195;
    wire N__45190;
    wire N__45185;
    wire N__45182;
    wire N__45181;
    wire N__45180;
    wire N__45179;
    wire N__45178;
    wire N__45177;
    wire N__45176;
    wire N__45173;
    wire N__45170;
    wire N__45163;
    wire N__45152;
    wire N__45149;
    wire N__45148;
    wire N__45147;
    wire N__45146;
    wire N__45145;
    wire N__45144;
    wire N__45143;
    wire N__45142;
    wire N__45141;
    wire N__45140;
    wire N__45139;
    wire N__45138;
    wire N__45137;
    wire N__45136;
    wire N__45135;
    wire N__45134;
    wire N__45133;
    wire N__45132;
    wire N__45131;
    wire N__45130;
    wire N__45129;
    wire N__45128;
    wire N__45127;
    wire N__45126;
    wire N__45125;
    wire N__45120;
    wire N__45113;
    wire N__45102;
    wire N__45099;
    wire N__45098;
    wire N__45095;
    wire N__45092;
    wire N__45085;
    wire N__45080;
    wire N__45077;
    wire N__45074;
    wire N__45071;
    wire N__45070;
    wire N__45067;
    wire N__45066;
    wire N__45065;
    wire N__45062;
    wire N__45061;
    wire N__45060;
    wire N__45059;
    wire N__45058;
    wire N__45055;
    wire N__45052;
    wire N__45051;
    wire N__45048;
    wire N__45047;
    wire N__45046;
    wire N__45045;
    wire N__45044;
    wire N__45043;
    wire N__45042;
    wire N__45041;
    wire N__45032;
    wire N__45023;
    wire N__45022;
    wire N__45019;
    wire N__45018;
    wire N__45015;
    wire N__45014;
    wire N__45011;
    wire N__45010;
    wire N__45009;
    wire N__45008;
    wire N__45005;
    wire N__45004;
    wire N__45001;
    wire N__45000;
    wire N__44997;
    wire N__44996;
    wire N__44995;
    wire N__44992;
    wire N__44991;
    wire N__44988;
    wire N__44987;
    wire N__44984;
    wire N__44983;
    wire N__44980;
    wire N__44977;
    wire N__44976;
    wire N__44973;
    wire N__44972;
    wire N__44969;
    wire N__44968;
    wire N__44965;
    wire N__44964;
    wire N__44961;
    wire N__44960;
    wire N__44957;
    wire N__44956;
    wire N__44953;
    wire N__44952;
    wire N__44949;
    wire N__44948;
    wire N__44945;
    wire N__44944;
    wire N__44941;
    wire N__44940;
    wire N__44937;
    wire N__44936;
    wire N__44931;
    wire N__44928;
    wire N__44925;
    wire N__44922;
    wire N__44917;
    wire N__44914;
    wire N__44905;
    wire N__44902;
    wire N__44893;
    wire N__44876;
    wire N__44875;
    wire N__44872;
    wire N__44871;
    wire N__44868;
    wire N__44867;
    wire N__44864;
    wire N__44863;
    wire N__44860;
    wire N__44857;
    wire N__44856;
    wire N__44853;
    wire N__44852;
    wire N__44849;
    wire N__44848;
    wire N__44843;
    wire N__44828;
    wire N__44811;
    wire N__44794;
    wire N__44777;
    wire N__44760;
    wire N__44747;
    wire N__44744;
    wire N__44735;
    wire N__44730;
    wire N__44727;
    wire N__44722;
    wire N__44705;
    wire N__44692;
    wire N__44677;
    wire N__44660;
    wire N__44659;
    wire N__44658;
    wire N__44657;
    wire N__44656;
    wire N__44655;
    wire N__44654;
    wire N__44653;
    wire N__44652;
    wire N__44651;
    wire N__44650;
    wire N__44649;
    wire N__44648;
    wire N__44647;
    wire N__44646;
    wire N__44645;
    wire N__44644;
    wire N__44639;
    wire N__44630;
    wire N__44629;
    wire N__44628;
    wire N__44627;
    wire N__44626;
    wire N__44625;
    wire N__44624;
    wire N__44623;
    wire N__44622;
    wire N__44621;
    wire N__44620;
    wire N__44619;
    wire N__44618;
    wire N__44615;
    wire N__44612;
    wire N__44611;
    wire N__44610;
    wire N__44609;
    wire N__44606;
    wire N__44595;
    wire N__44594;
    wire N__44593;
    wire N__44592;
    wire N__44591;
    wire N__44590;
    wire N__44587;
    wire N__44586;
    wire N__44583;
    wire N__44580;
    wire N__44579;
    wire N__44578;
    wire N__44577;
    wire N__44576;
    wire N__44575;
    wire N__44574;
    wire N__44573;
    wire N__44568;
    wire N__44557;
    wire N__44554;
    wire N__44547;
    wire N__44540;
    wire N__44535;
    wire N__44534;
    wire N__44531;
    wire N__44528;
    wire N__44525;
    wire N__44520;
    wire N__44509;
    wire N__44506;
    wire N__44503;
    wire N__44500;
    wire N__44497;
    wire N__44492;
    wire N__44481;
    wire N__44480;
    wire N__44479;
    wire N__44478;
    wire N__44477;
    wire N__44476;
    wire N__44471;
    wire N__44466;
    wire N__44465;
    wire N__44464;
    wire N__44463;
    wire N__44458;
    wire N__44457;
    wire N__44456;
    wire N__44453;
    wire N__44442;
    wire N__44437;
    wire N__44428;
    wire N__44427;
    wire N__44426;
    wire N__44425;
    wire N__44424;
    wire N__44423;
    wire N__44422;
    wire N__44421;
    wire N__44420;
    wire N__44419;
    wire N__44418;
    wire N__44417;
    wire N__44414;
    wire N__44413;
    wire N__44412;
    wire N__44409;
    wire N__44408;
    wire N__44401;
    wire N__44396;
    wire N__44389;
    wire N__44386;
    wire N__44381;
    wire N__44376;
    wire N__44371;
    wire N__44364;
    wire N__44353;
    wire N__44348;
    wire N__44345;
    wire N__44334;
    wire N__44327;
    wire N__44306;
    wire N__44303;
    wire N__44300;
    wire N__44297;
    wire N__44294;
    wire N__44291;
    wire N__44288;
    wire N__44285;
    wire N__44282;
    wire N__44279;
    wire N__44276;
    wire N__44273;
    wire N__44270;
    wire N__44267;
    wire N__44264;
    wire N__44261;
    wire N__44258;
    wire N__44255;
    wire N__44254;
    wire N__44249;
    wire N__44246;
    wire N__44243;
    wire N__44242;
    wire N__44239;
    wire N__44236;
    wire N__44233;
    wire N__44230;
    wire N__44227;
    wire N__44224;
    wire N__44219;
    wire N__44216;
    wire N__44213;
    wire N__44210;
    wire N__44207;
    wire N__44204;
    wire N__44201;
    wire N__44198;
    wire N__44197;
    wire N__44194;
    wire N__44193;
    wire N__44190;
    wire N__44187;
    wire N__44184;
    wire N__44177;
    wire N__44174;
    wire N__44171;
    wire N__44168;
    wire N__44165;
    wire N__44162;
    wire N__44159;
    wire N__44156;
    wire N__44155;
    wire N__44152;
    wire N__44149;
    wire N__44146;
    wire N__44145;
    wire N__44142;
    wire N__44139;
    wire N__44136;
    wire N__44129;
    wire N__44126;
    wire N__44123;
    wire N__44120;
    wire N__44117;
    wire N__44114;
    wire N__44111;
    wire N__44108;
    wire N__44105;
    wire N__44102;
    wire N__44099;
    wire N__44098;
    wire N__44095;
    wire N__44094;
    wire N__44093;
    wire N__44092;
    wire N__44089;
    wire N__44088;
    wire N__44087;
    wire N__44086;
    wire N__44085;
    wire N__44084;
    wire N__44083;
    wire N__44082;
    wire N__44081;
    wire N__44080;
    wire N__44079;
    wire N__44078;
    wire N__44077;
    wire N__44076;
    wire N__44075;
    wire N__44072;
    wire N__44067;
    wire N__44066;
    wire N__44065;
    wire N__44062;
    wire N__44055;
    wire N__44052;
    wire N__44037;
    wire N__44034;
    wire N__44031;
    wire N__44026;
    wire N__44025;
    wire N__44020;
    wire N__44015;
    wire N__44014;
    wire N__44007;
    wire N__44004;
    wire N__44001;
    wire N__43998;
    wire N__43997;
    wire N__43996;
    wire N__43993;
    wire N__43990;
    wire N__43987;
    wire N__43984;
    wire N__43981;
    wire N__43976;
    wire N__43973;
    wire N__43970;
    wire N__43967;
    wire N__43964;
    wire N__43961;
    wire N__43956;
    wire N__43947;
    wire N__43944;
    wire N__43931;
    wire N__43928;
    wire N__43927;
    wire N__43924;
    wire N__43923;
    wire N__43920;
    wire N__43917;
    wire N__43914;
    wire N__43907;
    wire N__43904;
    wire N__43901;
    wire N__43898;
    wire N__43895;
    wire N__43892;
    wire N__43889;
    wire N__43886;
    wire N__43883;
    wire N__43882;
    wire N__43879;
    wire N__43876;
    wire N__43873;
    wire N__43872;
    wire N__43869;
    wire N__43866;
    wire N__43863;
    wire N__43856;
    wire N__43853;
    wire N__43850;
    wire N__43847;
    wire N__43844;
    wire N__43841;
    wire N__43838;
    wire N__43835;
    wire N__43832;
    wire N__43829;
    wire N__43826;
    wire N__43823;
    wire N__43820;
    wire N__43817;
    wire N__43814;
    wire N__43811;
    wire N__43810;
    wire N__43807;
    wire N__43802;
    wire N__43801;
    wire N__43798;
    wire N__43797;
    wire N__43794;
    wire N__43791;
    wire N__43788;
    wire N__43785;
    wire N__43778;
    wire N__43775;
    wire N__43772;
    wire N__43769;
    wire N__43766;
    wire N__43763;
    wire N__43760;
    wire N__43759;
    wire N__43758;
    wire N__43751;
    wire N__43748;
    wire N__43747;
    wire N__43746;
    wire N__43745;
    wire N__43736;
    wire N__43733;
    wire N__43730;
    wire N__43727;
    wire N__43724;
    wire N__43721;
    wire N__43718;
    wire N__43715;
    wire N__43712;
    wire N__43709;
    wire N__43708;
    wire N__43705;
    wire N__43702;
    wire N__43701;
    wire N__43698;
    wire N__43693;
    wire N__43690;
    wire N__43687;
    wire N__43682;
    wire N__43679;
    wire N__43676;
    wire N__43673;
    wire N__43670;
    wire N__43667;
    wire N__43664;
    wire N__43663;
    wire N__43660;
    wire N__43657;
    wire N__43654;
    wire N__43651;
    wire N__43650;
    wire N__43647;
    wire N__43644;
    wire N__43641;
    wire N__43638;
    wire N__43635;
    wire N__43632;
    wire N__43625;
    wire N__43622;
    wire N__43619;
    wire N__43616;
    wire N__43613;
    wire N__43612;
    wire N__43611;
    wire N__43608;
    wire N__43605;
    wire N__43602;
    wire N__43599;
    wire N__43596;
    wire N__43593;
    wire N__43586;
    wire N__43583;
    wire N__43580;
    wire N__43577;
    wire N__43574;
    wire N__43571;
    wire N__43568;
    wire N__43565;
    wire N__43562;
    wire N__43559;
    wire N__43556;
    wire N__43553;
    wire N__43552;
    wire N__43549;
    wire N__43546;
    wire N__43545;
    wire N__43542;
    wire N__43539;
    wire N__43536;
    wire N__43533;
    wire N__43526;
    wire N__43523;
    wire N__43520;
    wire N__43517;
    wire N__43514;
    wire N__43511;
    wire N__43508;
    wire N__43505;
    wire N__43504;
    wire N__43501;
    wire N__43498;
    wire N__43497;
    wire N__43494;
    wire N__43491;
    wire N__43488;
    wire N__43483;
    wire N__43480;
    wire N__43475;
    wire N__43472;
    wire N__43469;
    wire N__43466;
    wire N__43463;
    wire N__43460;
    wire N__43457;
    wire N__43454;
    wire N__43451;
    wire N__43448;
    wire N__43447;
    wire N__43444;
    wire N__43441;
    wire N__43436;
    wire N__43433;
    wire N__43432;
    wire N__43429;
    wire N__43426;
    wire N__43421;
    wire N__43418;
    wire N__43417;
    wire N__43414;
    wire N__43411;
    wire N__43406;
    wire N__43403;
    wire N__43402;
    wire N__43399;
    wire N__43396;
    wire N__43391;
    wire N__43388;
    wire N__43387;
    wire N__43384;
    wire N__43381;
    wire N__43376;
    wire N__43373;
    wire N__43372;
    wire N__43371;
    wire N__43370;
    wire N__43369;
    wire N__43368;
    wire N__43367;
    wire N__43364;
    wire N__43355;
    wire N__43352;
    wire N__43351;
    wire N__43348;
    wire N__43345;
    wire N__43340;
    wire N__43339;
    wire N__43338;
    wire N__43337;
    wire N__43336;
    wire N__43335;
    wire N__43334;
    wire N__43333;
    wire N__43332;
    wire N__43331;
    wire N__43330;
    wire N__43329;
    wire N__43328;
    wire N__43327;
    wire N__43326;
    wire N__43323;
    wire N__43318;
    wire N__43315;
    wire N__43308;
    wire N__43299;
    wire N__43296;
    wire N__43291;
    wire N__43282;
    wire N__43265;
    wire N__43262;
    wire N__43261;
    wire N__43258;
    wire N__43255;
    wire N__43250;
    wire N__43249;
    wire N__43248;
    wire N__43245;
    wire N__43242;
    wire N__43239;
    wire N__43232;
    wire N__43229;
    wire N__43226;
    wire N__43223;
    wire N__43220;
    wire N__43217;
    wire N__43214;
    wire N__43211;
    wire N__43208;
    wire N__43205;
    wire N__43202;
    wire N__43199;
    wire N__43196;
    wire N__43193;
    wire N__43190;
    wire N__43187;
    wire N__43184;
    wire N__43181;
    wire N__43180;
    wire N__43177;
    wire N__43174;
    wire N__43169;
    wire N__43166;
    wire N__43165;
    wire N__43162;
    wire N__43159;
    wire N__43154;
    wire N__43151;
    wire N__43150;
    wire N__43147;
    wire N__43144;
    wire N__43139;
    wire N__43136;
    wire N__43135;
    wire N__43132;
    wire N__43129;
    wire N__43124;
    wire N__43121;
    wire N__43120;
    wire N__43117;
    wire N__43114;
    wire N__43109;
    wire N__43106;
    wire N__43105;
    wire N__43102;
    wire N__43099;
    wire N__43094;
    wire N__43091;
    wire N__43090;
    wire N__43087;
    wire N__43084;
    wire N__43079;
    wire N__43076;
    wire N__43075;
    wire N__43072;
    wire N__43069;
    wire N__43064;
    wire N__43061;
    wire N__43058;
    wire N__43055;
    wire N__43054;
    wire N__43051;
    wire N__43048;
    wire N__43043;
    wire N__43040;
    wire N__43037;
    wire N__43034;
    wire N__43031;
    wire N__43030;
    wire N__43025;
    wire N__43024;
    wire N__43023;
    wire N__43022;
    wire N__43021;
    wire N__43020;
    wire N__43017;
    wire N__43016;
    wire N__43013;
    wire N__43010;
    wire N__43005;
    wire N__43002;
    wire N__42999;
    wire N__42996;
    wire N__42989;
    wire N__42980;
    wire N__42979;
    wire N__42976;
    wire N__42975;
    wire N__42972;
    wire N__42971;
    wire N__42968;
    wire N__42965;
    wire N__42962;
    wire N__42959;
    wire N__42958;
    wire N__42955;
    wire N__42952;
    wire N__42949;
    wire N__42946;
    wire N__42945;
    wire N__42944;
    wire N__42941;
    wire N__42938;
    wire N__42931;
    wire N__42926;
    wire N__42923;
    wire N__42914;
    wire N__42911;
    wire N__42908;
    wire N__42907;
    wire N__42904;
    wire N__42901;
    wire N__42900;
    wire N__42897;
    wire N__42894;
    wire N__42891;
    wire N__42888;
    wire N__42885;
    wire N__42878;
    wire N__42875;
    wire N__42872;
    wire N__42869;
    wire N__42866;
    wire N__42865;
    wire N__42864;
    wire N__42861;
    wire N__42858;
    wire N__42855;
    wire N__42852;
    wire N__42845;
    wire N__42844;
    wire N__42841;
    wire N__42840;
    wire N__42839;
    wire N__42836;
    wire N__42833;
    wire N__42830;
    wire N__42827;
    wire N__42824;
    wire N__42821;
    wire N__42816;
    wire N__42813;
    wire N__42806;
    wire N__42803;
    wire N__42800;
    wire N__42797;
    wire N__42796;
    wire N__42795;
    wire N__42792;
    wire N__42789;
    wire N__42786;
    wire N__42783;
    wire N__42780;
    wire N__42777;
    wire N__42774;
    wire N__42771;
    wire N__42764;
    wire N__42763;
    wire N__42760;
    wire N__42757;
    wire N__42752;
    wire N__42749;
    wire N__42746;
    wire N__42743;
    wire N__42740;
    wire N__42739;
    wire N__42736;
    wire N__42733;
    wire N__42728;
    wire N__42725;
    wire N__42724;
    wire N__42721;
    wire N__42718;
    wire N__42713;
    wire N__42710;
    wire N__42709;
    wire N__42706;
    wire N__42703;
    wire N__42698;
    wire N__42695;
    wire N__42692;
    wire N__42691;
    wire N__42690;
    wire N__42687;
    wire N__42684;
    wire N__42681;
    wire N__42678;
    wire N__42671;
    wire N__42668;
    wire N__42665;
    wire N__42662;
    wire N__42661;
    wire N__42658;
    wire N__42655;
    wire N__42652;
    wire N__42647;
    wire N__42644;
    wire N__42641;
    wire N__42638;
    wire N__42635;
    wire N__42632;
    wire N__42629;
    wire N__42626;
    wire N__42625;
    wire N__42622;
    wire N__42621;
    wire N__42618;
    wire N__42615;
    wire N__42614;
    wire N__42611;
    wire N__42608;
    wire N__42605;
    wire N__42602;
    wire N__42593;
    wire N__42590;
    wire N__42587;
    wire N__42586;
    wire N__42583;
    wire N__42580;
    wire N__42577;
    wire N__42574;
    wire N__42571;
    wire N__42568;
    wire N__42567;
    wire N__42564;
    wire N__42561;
    wire N__42558;
    wire N__42551;
    wire N__42548;
    wire N__42545;
    wire N__42542;
    wire N__42539;
    wire N__42536;
    wire N__42535;
    wire N__42534;
    wire N__42533;
    wire N__42532;
    wire N__42531;
    wire N__42530;
    wire N__42529;
    wire N__42528;
    wire N__42527;
    wire N__42526;
    wire N__42525;
    wire N__42524;
    wire N__42523;
    wire N__42522;
    wire N__42521;
    wire N__42520;
    wire N__42519;
    wire N__42518;
    wire N__42517;
    wire N__42516;
    wire N__42515;
    wire N__42514;
    wire N__42513;
    wire N__42512;
    wire N__42511;
    wire N__42510;
    wire N__42499;
    wire N__42494;
    wire N__42479;
    wire N__42468;
    wire N__42467;
    wire N__42454;
    wire N__42453;
    wire N__42452;
    wire N__42451;
    wire N__42450;
    wire N__42445;
    wire N__42442;
    wire N__42439;
    wire N__42434;
    wire N__42433;
    wire N__42432;
    wire N__42431;
    wire N__42428;
    wire N__42425;
    wire N__42422;
    wire N__42419;
    wire N__42414;
    wire N__42409;
    wire N__42404;
    wire N__42397;
    wire N__42388;
    wire N__42377;
    wire N__42374;
    wire N__42373;
    wire N__42370;
    wire N__42367;
    wire N__42366;
    wire N__42361;
    wire N__42360;
    wire N__42357;
    wire N__42354;
    wire N__42351;
    wire N__42344;
    wire N__42341;
    wire N__42338;
    wire N__42335;
    wire N__42332;
    wire N__42331;
    wire N__42328;
    wire N__42325;
    wire N__42322;
    wire N__42319;
    wire N__42316;
    wire N__42313;
    wire N__42308;
    wire N__42307;
    wire N__42306;
    wire N__42305;
    wire N__42304;
    wire N__42303;
    wire N__42300;
    wire N__42297;
    wire N__42296;
    wire N__42295;
    wire N__42294;
    wire N__42293;
    wire N__42292;
    wire N__42291;
    wire N__42290;
    wire N__42289;
    wire N__42282;
    wire N__42279;
    wire N__42268;
    wire N__42261;
    wire N__42256;
    wire N__42253;
    wire N__42242;
    wire N__42241;
    wire N__42240;
    wire N__42239;
    wire N__42236;
    wire N__42233;
    wire N__42232;
    wire N__42231;
    wire N__42228;
    wire N__42225;
    wire N__42224;
    wire N__42223;
    wire N__42222;
    wire N__42221;
    wire N__42220;
    wire N__42217;
    wire N__42212;
    wire N__42209;
    wire N__42206;
    wire N__42203;
    wire N__42200;
    wire N__42191;
    wire N__42186;
    wire N__42183;
    wire N__42170;
    wire N__42169;
    wire N__42166;
    wire N__42165;
    wire N__42164;
    wire N__42161;
    wire N__42158;
    wire N__42155;
    wire N__42154;
    wire N__42151;
    wire N__42148;
    wire N__42145;
    wire N__42142;
    wire N__42139;
    wire N__42128;
    wire N__42125;
    wire N__42122;
    wire N__42119;
    wire N__42118;
    wire N__42117;
    wire N__42116;
    wire N__42115;
    wire N__42112;
    wire N__42109;
    wire N__42106;
    wire N__42103;
    wire N__42102;
    wire N__42099;
    wire N__42098;
    wire N__42097;
    wire N__42096;
    wire N__42095;
    wire N__42094;
    wire N__42093;
    wire N__42092;
    wire N__42091;
    wire N__42090;
    wire N__42089;
    wire N__42088;
    wire N__42087;
    wire N__42084;
    wire N__42083;
    wire N__42082;
    wire N__42081;
    wire N__42076;
    wire N__42073;
    wire N__42072;
    wire N__42071;
    wire N__42070;
    wire N__42069;
    wire N__42066;
    wire N__42063;
    wire N__42060;
    wire N__42051;
    wire N__42048;
    wire N__42039;
    wire N__42034;
    wire N__42031;
    wire N__42024;
    wire N__42019;
    wire N__42010;
    wire N__42007;
    wire N__42004;
    wire N__42001;
    wire N__41994;
    wire N__41991;
    wire N__41982;
    wire N__41979;
    wire N__41976;
    wire N__41973;
    wire N__41968;
    wire N__41965;
    wire N__41960;
    wire N__41951;
    wire N__41948;
    wire N__41945;
    wire N__41942;
    wire N__41939;
    wire N__41936;
    wire N__41933;
    wire N__41930;
    wire N__41927;
    wire N__41924;
    wire N__41921;
    wire N__41918;
    wire N__41915;
    wire N__41912;
    wire N__41909;
    wire N__41906;
    wire N__41903;
    wire N__41900;
    wire N__41897;
    wire N__41896;
    wire N__41893;
    wire N__41890;
    wire N__41885;
    wire N__41882;
    wire N__41879;
    wire N__41878;
    wire N__41877;
    wire N__41874;
    wire N__41869;
    wire N__41864;
    wire N__41861;
    wire N__41860;
    wire N__41857;
    wire N__41856;
    wire N__41853;
    wire N__41850;
    wire N__41847;
    wire N__41846;
    wire N__41845;
    wire N__41842;
    wire N__41837;
    wire N__41832;
    wire N__41825;
    wire N__41824;
    wire N__41823;
    wire N__41822;
    wire N__41821;
    wire N__41820;
    wire N__41817;
    wire N__41816;
    wire N__41815;
    wire N__41812;
    wire N__41811;
    wire N__41810;
    wire N__41809;
    wire N__41806;
    wire N__41805;
    wire N__41804;
    wire N__41803;
    wire N__41800;
    wire N__41797;
    wire N__41796;
    wire N__41793;
    wire N__41790;
    wire N__41787;
    wire N__41786;
    wire N__41783;
    wire N__41780;
    wire N__41777;
    wire N__41774;
    wire N__41771;
    wire N__41770;
    wire N__41769;
    wire N__41768;
    wire N__41765;
    wire N__41762;
    wire N__41755;
    wire N__41754;
    wire N__41753;
    wire N__41752;
    wire N__41751;
    wire N__41750;
    wire N__41747;
    wire N__41744;
    wire N__41743;
    wire N__41738;
    wire N__41731;
    wire N__41728;
    wire N__41725;
    wire N__41722;
    wire N__41721;
    wire N__41718;
    wire N__41715;
    wire N__41712;
    wire N__41709;
    wire N__41706;
    wire N__41701;
    wire N__41700;
    wire N__41697;
    wire N__41694;
    wire N__41691;
    wire N__41690;
    wire N__41689;
    wire N__41686;
    wire N__41685;
    wire N__41682;
    wire N__41679;
    wire N__41674;
    wire N__41669;
    wire N__41662;
    wire N__41659;
    wire N__41656;
    wire N__41653;
    wire N__41650;
    wire N__41647;
    wire N__41642;
    wire N__41635;
    wire N__41622;
    wire N__41617;
    wire N__41612;
    wire N__41609;
    wire N__41588;
    wire N__41587;
    wire N__41586;
    wire N__41585;
    wire N__41584;
    wire N__41583;
    wire N__41582;
    wire N__41579;
    wire N__41576;
    wire N__41573;
    wire N__41570;
    wire N__41565;
    wire N__41562;
    wire N__41561;
    wire N__41556;
    wire N__41555;
    wire N__41552;
    wire N__41547;
    wire N__41544;
    wire N__41541;
    wire N__41538;
    wire N__41535;
    wire N__41530;
    wire N__41525;
    wire N__41516;
    wire N__41513;
    wire N__41510;
    wire N__41507;
    wire N__41504;
    wire N__41503;
    wire N__41500;
    wire N__41499;
    wire N__41498;
    wire N__41497;
    wire N__41496;
    wire N__41493;
    wire N__41490;
    wire N__41487;
    wire N__41484;
    wire N__41481;
    wire N__41480;
    wire N__41479;
    wire N__41476;
    wire N__41469;
    wire N__41466;
    wire N__41461;
    wire N__41458;
    wire N__41453;
    wire N__41450;
    wire N__41441;
    wire N__41438;
    wire N__41435;
    wire N__41432;
    wire N__41431;
    wire N__41430;
    wire N__41427;
    wire N__41422;
    wire N__41419;
    wire N__41414;
    wire N__41413;
    wire N__41410;
    wire N__41407;
    wire N__41402;
    wire N__41399;
    wire N__41396;
    wire N__41393;
    wire N__41390;
    wire N__41387;
    wire N__41384;
    wire N__41381;
    wire N__41378;
    wire N__41375;
    wire N__41372;
    wire N__41369;
    wire N__41366;
    wire N__41363;
    wire N__41360;
    wire N__41357;
    wire N__41354;
    wire N__41351;
    wire N__41348;
    wire N__41345;
    wire N__41342;
    wire N__41339;
    wire N__41336;
    wire N__41333;
    wire N__41330;
    wire N__41327;
    wire N__41324;
    wire N__41321;
    wire N__41318;
    wire N__41315;
    wire N__41312;
    wire N__41309;
    wire N__41306;
    wire N__41303;
    wire N__41300;
    wire N__41297;
    wire N__41294;
    wire N__41291;
    wire N__41288;
    wire N__41285;
    wire N__41284;
    wire N__41281;
    wire N__41278;
    wire N__41273;
    wire N__41272;
    wire N__41269;
    wire N__41266;
    wire N__41261;
    wire N__41258;
    wire N__41255;
    wire N__41252;
    wire N__41249;
    wire N__41246;
    wire N__41243;
    wire N__41240;
    wire N__41237;
    wire N__41234;
    wire N__41231;
    wire N__41228;
    wire N__41225;
    wire N__41222;
    wire N__41219;
    wire N__41216;
    wire N__41215;
    wire N__41212;
    wire N__41209;
    wire N__41208;
    wire N__41205;
    wire N__41202;
    wire N__41199;
    wire N__41196;
    wire N__41193;
    wire N__41190;
    wire N__41185;
    wire N__41182;
    wire N__41177;
    wire N__41174;
    wire N__41171;
    wire N__41168;
    wire N__41165;
    wire N__41162;
    wire N__41159;
    wire N__41156;
    wire N__41155;
    wire N__41152;
    wire N__41149;
    wire N__41148;
    wire N__41145;
    wire N__41142;
    wire N__41139;
    wire N__41136;
    wire N__41129;
    wire N__41126;
    wire N__41123;
    wire N__41120;
    wire N__41117;
    wire N__41114;
    wire N__41111;
    wire N__41108;
    wire N__41107;
    wire N__41106;
    wire N__41103;
    wire N__41098;
    wire N__41095;
    wire N__41092;
    wire N__41087;
    wire N__41084;
    wire N__41081;
    wire N__41078;
    wire N__41075;
    wire N__41072;
    wire N__41071;
    wire N__41068;
    wire N__41065;
    wire N__41064;
    wire N__41061;
    wire N__41058;
    wire N__41055;
    wire N__41048;
    wire N__41045;
    wire N__41042;
    wire N__41039;
    wire N__41036;
    wire N__41033;
    wire N__41030;
    wire N__41027;
    wire N__41024;
    wire N__41021;
    wire N__41018;
    wire N__41015;
    wire N__41012;
    wire N__41009;
    wire N__41006;
    wire N__41003;
    wire N__41002;
    wire N__40999;
    wire N__40996;
    wire N__40995;
    wire N__40992;
    wire N__40987;
    wire N__40984;
    wire N__40981;
    wire N__40976;
    wire N__40973;
    wire N__40970;
    wire N__40969;
    wire N__40966;
    wire N__40965;
    wire N__40960;
    wire N__40957;
    wire N__40952;
    wire N__40949;
    wire N__40946;
    wire N__40943;
    wire N__40942;
    wire N__40941;
    wire N__40938;
    wire N__40935;
    wire N__40932;
    wire N__40929;
    wire N__40926;
    wire N__40921;
    wire N__40916;
    wire N__40913;
    wire N__40912;
    wire N__40911;
    wire N__40906;
    wire N__40903;
    wire N__40900;
    wire N__40897;
    wire N__40894;
    wire N__40889;
    wire N__40886;
    wire N__40883;
    wire N__40880;
    wire N__40879;
    wire N__40876;
    wire N__40875;
    wire N__40872;
    wire N__40867;
    wire N__40862;
    wire N__40859;
    wire N__40856;
    wire N__40853;
    wire N__40850;
    wire N__40847;
    wire N__40844;
    wire N__40841;
    wire N__40838;
    wire N__40835;
    wire N__40832;
    wire N__40829;
    wire N__40828;
    wire N__40827;
    wire N__40826;
    wire N__40823;
    wire N__40820;
    wire N__40817;
    wire N__40814;
    wire N__40811;
    wire N__40808;
    wire N__40799;
    wire N__40798;
    wire N__40793;
    wire N__40792;
    wire N__40789;
    wire N__40786;
    wire N__40781;
    wire N__40778;
    wire N__40775;
    wire N__40774;
    wire N__40771;
    wire N__40768;
    wire N__40763;
    wire N__40762;
    wire N__40759;
    wire N__40756;
    wire N__40751;
    wire N__40748;
    wire N__40745;
    wire N__40742;
    wire N__40739;
    wire N__40736;
    wire N__40733;
    wire N__40732;
    wire N__40731;
    wire N__40726;
    wire N__40723;
    wire N__40718;
    wire N__40715;
    wire N__40714;
    wire N__40713;
    wire N__40708;
    wire N__40705;
    wire N__40700;
    wire N__40697;
    wire N__40696;
    wire N__40695;
    wire N__40690;
    wire N__40687;
    wire N__40682;
    wire N__40679;
    wire N__40676;
    wire N__40673;
    wire N__40670;
    wire N__40667;
    wire N__40664;
    wire N__40661;
    wire N__40658;
    wire N__40655;
    wire N__40652;
    wire N__40649;
    wire N__40646;
    wire N__40643;
    wire N__40640;
    wire N__40637;
    wire N__40636;
    wire N__40633;
    wire N__40630;
    wire N__40627;
    wire N__40624;
    wire N__40619;
    wire N__40616;
    wire N__40613;
    wire N__40612;
    wire N__40609;
    wire N__40606;
    wire N__40605;
    wire N__40602;
    wire N__40601;
    wire N__40598;
    wire N__40595;
    wire N__40592;
    wire N__40589;
    wire N__40586;
    wire N__40583;
    wire N__40578;
    wire N__40575;
    wire N__40572;
    wire N__40565;
    wire N__40562;
    wire N__40559;
    wire N__40556;
    wire N__40553;
    wire N__40550;
    wire N__40547;
    wire N__40546;
    wire N__40543;
    wire N__40540;
    wire N__40537;
    wire N__40536;
    wire N__40533;
    wire N__40530;
    wire N__40527;
    wire N__40524;
    wire N__40521;
    wire N__40520;
    wire N__40519;
    wire N__40512;
    wire N__40507;
    wire N__40502;
    wire N__40499;
    wire N__40496;
    wire N__40493;
    wire N__40490;
    wire N__40487;
    wire N__40484;
    wire N__40481;
    wire N__40480;
    wire N__40479;
    wire N__40476;
    wire N__40475;
    wire N__40472;
    wire N__40469;
    wire N__40466;
    wire N__40463;
    wire N__40454;
    wire N__40451;
    wire N__40448;
    wire N__40445;
    wire N__40442;
    wire N__40439;
    wire N__40436;
    wire N__40433;
    wire N__40430;
    wire N__40427;
    wire N__40424;
    wire N__40421;
    wire N__40418;
    wire N__40415;
    wire N__40412;
    wire N__40409;
    wire N__40406;
    wire N__40403;
    wire N__40400;
    wire N__40397;
    wire N__40394;
    wire N__40391;
    wire N__40388;
    wire N__40385;
    wire N__40382;
    wire N__40379;
    wire N__40376;
    wire N__40373;
    wire N__40370;
    wire N__40367;
    wire N__40364;
    wire N__40361;
    wire N__40358;
    wire N__40355;
    wire N__40352;
    wire N__40349;
    wire N__40346;
    wire N__40343;
    wire N__40340;
    wire N__40337;
    wire N__40334;
    wire N__40331;
    wire N__40328;
    wire N__40325;
    wire N__40322;
    wire N__40319;
    wire N__40316;
    wire N__40313;
    wire N__40310;
    wire N__40307;
    wire N__40304;
    wire N__40301;
    wire N__40298;
    wire N__40295;
    wire N__40292;
    wire N__40289;
    wire N__40286;
    wire N__40283;
    wire N__40280;
    wire N__40277;
    wire N__40274;
    wire N__40271;
    wire N__40268;
    wire N__40265;
    wire N__40262;
    wire N__40259;
    wire N__40256;
    wire N__40253;
    wire N__40250;
    wire N__40247;
    wire N__40244;
    wire N__40241;
    wire N__40238;
    wire N__40235;
    wire N__40232;
    wire N__40229;
    wire N__40226;
    wire N__40223;
    wire N__40220;
    wire N__40217;
    wire N__40214;
    wire N__40211;
    wire N__40208;
    wire N__40205;
    wire N__40202;
    wire N__40199;
    wire N__40196;
    wire N__40193;
    wire N__40190;
    wire N__40187;
    wire N__40184;
    wire N__40181;
    wire N__40178;
    wire N__40175;
    wire N__40172;
    wire N__40169;
    wire N__40166;
    wire N__40163;
    wire N__40160;
    wire N__40157;
    wire N__40154;
    wire N__40151;
    wire N__40148;
    wire N__40145;
    wire N__40142;
    wire N__40139;
    wire N__40136;
    wire N__40133;
    wire N__40132;
    wire N__40131;
    wire N__40128;
    wire N__40127;
    wire N__40124;
    wire N__40121;
    wire N__40118;
    wire N__40115;
    wire N__40110;
    wire N__40103;
    wire N__40100;
    wire N__40097;
    wire N__40096;
    wire N__40095;
    wire N__40092;
    wire N__40089;
    wire N__40086;
    wire N__40079;
    wire N__40078;
    wire N__40077;
    wire N__40076;
    wire N__40075;
    wire N__40072;
    wire N__40069;
    wire N__40068;
    wire N__40063;
    wire N__40060;
    wire N__40059;
    wire N__40058;
    wire N__40057;
    wire N__40056;
    wire N__40053;
    wire N__40052;
    wire N__40049;
    wire N__40046;
    wire N__40045;
    wire N__40040;
    wire N__40039;
    wire N__40038;
    wire N__40037;
    wire N__40036;
    wire N__40035;
    wire N__40034;
    wire N__40033;
    wire N__40032;
    wire N__40031;
    wire N__40030;
    wire N__40023;
    wire N__40020;
    wire N__40017;
    wire N__40014;
    wire N__40011;
    wire N__40008;
    wire N__40005;
    wire N__40002;
    wire N__39995;
    wire N__39980;
    wire N__39975;
    wire N__39970;
    wire N__39953;
    wire N__39950;
    wire N__39947;
    wire N__39946;
    wire N__39943;
    wire N__39940;
    wire N__39935;
    wire N__39932;
    wire N__39929;
    wire N__39926;
    wire N__39925;
    wire N__39922;
    wire N__39919;
    wire N__39918;
    wire N__39917;
    wire N__39916;
    wire N__39913;
    wire N__39908;
    wire N__39903;
    wire N__39896;
    wire N__39893;
    wire N__39892;
    wire N__39891;
    wire N__39890;
    wire N__39889;
    wire N__39886;
    wire N__39883;
    wire N__39880;
    wire N__39875;
    wire N__39866;
    wire N__39863;
    wire N__39862;
    wire N__39861;
    wire N__39858;
    wire N__39855;
    wire N__39852;
    wire N__39845;
    wire N__39844;
    wire N__39841;
    wire N__39840;
    wire N__39839;
    wire N__39836;
    wire N__39833;
    wire N__39830;
    wire N__39827;
    wire N__39824;
    wire N__39815;
    wire N__39812;
    wire N__39811;
    wire N__39808;
    wire N__39807;
    wire N__39806;
    wire N__39803;
    wire N__39802;
    wire N__39801;
    wire N__39800;
    wire N__39797;
    wire N__39794;
    wire N__39791;
    wire N__39786;
    wire N__39781;
    wire N__39770;
    wire N__39767;
    wire N__39766;
    wire N__39765;
    wire N__39764;
    wire N__39763;
    wire N__39762;
    wire N__39761;
    wire N__39760;
    wire N__39759;
    wire N__39758;
    wire N__39757;
    wire N__39756;
    wire N__39755;
    wire N__39754;
    wire N__39753;
    wire N__39752;
    wire N__39749;
    wire N__39746;
    wire N__39745;
    wire N__39744;
    wire N__39743;
    wire N__39742;
    wire N__39739;
    wire N__39736;
    wire N__39735;
    wire N__39734;
    wire N__39733;
    wire N__39732;
    wire N__39725;
    wire N__39716;
    wire N__39715;
    wire N__39714;
    wire N__39713;
    wire N__39710;
    wire N__39707;
    wire N__39696;
    wire N__39689;
    wire N__39678;
    wire N__39673;
    wire N__39670;
    wire N__39667;
    wire N__39664;
    wire N__39659;
    wire N__39656;
    wire N__39635;
    wire N__39632;
    wire N__39629;
    wire N__39626;
    wire N__39623;
    wire N__39620;
    wire N__39617;
    wire N__39614;
    wire N__39611;
    wire N__39608;
    wire N__39605;
    wire N__39602;
    wire N__39599;
    wire N__39596;
    wire N__39593;
    wire N__39590;
    wire N__39587;
    wire N__39584;
    wire N__39581;
    wire N__39578;
    wire N__39575;
    wire N__39574;
    wire N__39571;
    wire N__39568;
    wire N__39565;
    wire N__39564;
    wire N__39559;
    wire N__39556;
    wire N__39551;
    wire N__39550;
    wire N__39549;
    wire N__39546;
    wire N__39541;
    wire N__39538;
    wire N__39533;
    wire N__39530;
    wire N__39527;
    wire N__39524;
    wire N__39521;
    wire N__39520;
    wire N__39517;
    wire N__39514;
    wire N__39513;
    wire N__39510;
    wire N__39509;
    wire N__39506;
    wire N__39503;
    wire N__39500;
    wire N__39497;
    wire N__39494;
    wire N__39485;
    wire N__39482;
    wire N__39479;
    wire N__39478;
    wire N__39477;
    wire N__39474;
    wire N__39471;
    wire N__39468;
    wire N__39461;
    wire N__39458;
    wire N__39455;
    wire N__39452;
    wire N__39449;
    wire N__39446;
    wire N__39443;
    wire N__39440;
    wire N__39437;
    wire N__39434;
    wire N__39431;
    wire N__39430;
    wire N__39429;
    wire N__39428;
    wire N__39427;
    wire N__39426;
    wire N__39425;
    wire N__39424;
    wire N__39423;
    wire N__39422;
    wire N__39421;
    wire N__39420;
    wire N__39419;
    wire N__39418;
    wire N__39417;
    wire N__39416;
    wire N__39415;
    wire N__39414;
    wire N__39413;
    wire N__39412;
    wire N__39411;
    wire N__39410;
    wire N__39409;
    wire N__39408;
    wire N__39407;
    wire N__39406;
    wire N__39405;
    wire N__39404;
    wire N__39403;
    wire N__39402;
    wire N__39393;
    wire N__39388;
    wire N__39379;
    wire N__39370;
    wire N__39361;
    wire N__39352;
    wire N__39343;
    wire N__39334;
    wire N__39321;
    wire N__39314;
    wire N__39311;
    wire N__39310;
    wire N__39307;
    wire N__39304;
    wire N__39303;
    wire N__39302;
    wire N__39299;
    wire N__39296;
    wire N__39293;
    wire N__39290;
    wire N__39285;
    wire N__39280;
    wire N__39275;
    wire N__39272;
    wire N__39271;
    wire N__39270;
    wire N__39269;
    wire N__39266;
    wire N__39263;
    wire N__39258;
    wire N__39251;
    wire N__39248;
    wire N__39245;
    wire N__39242;
    wire N__39239;
    wire N__39236;
    wire N__39233;
    wire N__39230;
    wire N__39227;
    wire N__39224;
    wire N__39221;
    wire N__39218;
    wire N__39215;
    wire N__39212;
    wire N__39209;
    wire N__39206;
    wire N__39203;
    wire N__39200;
    wire N__39197;
    wire N__39194;
    wire N__39191;
    wire N__39188;
    wire N__39185;
    wire N__39182;
    wire N__39179;
    wire N__39176;
    wire N__39173;
    wire N__39170;
    wire N__39167;
    wire N__39164;
    wire N__39161;
    wire N__39158;
    wire N__39155;
    wire N__39152;
    wire N__39149;
    wire N__39146;
    wire N__39143;
    wire N__39142;
    wire N__39141;
    wire N__39138;
    wire N__39135;
    wire N__39132;
    wire N__39127;
    wire N__39126;
    wire N__39121;
    wire N__39118;
    wire N__39115;
    wire N__39110;
    wire N__39107;
    wire N__39104;
    wire N__39101;
    wire N__39098;
    wire N__39095;
    wire N__39092;
    wire N__39089;
    wire N__39086;
    wire N__39083;
    wire N__39080;
    wire N__39077;
    wire N__39074;
    wire N__39071;
    wire N__39068;
    wire N__39067;
    wire N__39066;
    wire N__39065;
    wire N__39064;
    wire N__39063;
    wire N__39062;
    wire N__39061;
    wire N__39060;
    wire N__39059;
    wire N__39058;
    wire N__39057;
    wire N__39056;
    wire N__39055;
    wire N__39052;
    wire N__39049;
    wire N__39048;
    wire N__39047;
    wire N__39044;
    wire N__39043;
    wire N__39040;
    wire N__39039;
    wire N__39036;
    wire N__39035;
    wire N__39034;
    wire N__39033;
    wire N__39032;
    wire N__39031;
    wire N__39030;
    wire N__39029;
    wire N__39028;
    wire N__39027;
    wire N__39024;
    wire N__39023;
    wire N__39020;
    wire N__39019;
    wire N__39016;
    wire N__39015;
    wire N__39012;
    wire N__39011;
    wire N__39010;
    wire N__39009;
    wire N__39008;
    wire N__39007;
    wire N__38998;
    wire N__38997;
    wire N__38996;
    wire N__38995;
    wire N__38994;
    wire N__38993;
    wire N__38992;
    wire N__38991;
    wire N__38990;
    wire N__38989;
    wire N__38986;
    wire N__38985;
    wire N__38982;
    wire N__38979;
    wire N__38976;
    wire N__38975;
    wire N__38960;
    wire N__38951;
    wire N__38942;
    wire N__38925;
    wire N__38924;
    wire N__38923;
    wire N__38922;
    wire N__38919;
    wire N__38912;
    wire N__38909;
    wire N__38906;
    wire N__38899;
    wire N__38890;
    wire N__38883;
    wire N__38876;
    wire N__38873;
    wire N__38868;
    wire N__38863;
    wire N__38862;
    wire N__38859;
    wire N__38858;
    wire N__38855;
    wire N__38854;
    wire N__38851;
    wire N__38850;
    wire N__38845;
    wire N__38840;
    wire N__38835;
    wire N__38832;
    wire N__38829;
    wire N__38826;
    wire N__38821;
    wire N__38806;
    wire N__38803;
    wire N__38800;
    wire N__38799;
    wire N__38798;
    wire N__38795;
    wire N__38790;
    wire N__38783;
    wire N__38780;
    wire N__38777;
    wire N__38772;
    wire N__38769;
    wire N__38764;
    wire N__38757;
    wire N__38750;
    wire N__38747;
    wire N__38744;
    wire N__38741;
    wire N__38740;
    wire N__38737;
    wire N__38736;
    wire N__38735;
    wire N__38734;
    wire N__38733;
    wire N__38730;
    wire N__38729;
    wire N__38728;
    wire N__38727;
    wire N__38726;
    wire N__38725;
    wire N__38724;
    wire N__38723;
    wire N__38720;
    wire N__38711;
    wire N__38708;
    wire N__38693;
    wire N__38684;
    wire N__38681;
    wire N__38678;
    wire N__38675;
    wire N__38672;
    wire N__38669;
    wire N__38666;
    wire N__38663;
    wire N__38660;
    wire N__38657;
    wire N__38654;
    wire N__38651;
    wire N__38648;
    wire N__38645;
    wire N__38642;
    wire N__38639;
    wire N__38636;
    wire N__38633;
    wire N__38630;
    wire N__38627;
    wire N__38624;
    wire N__38621;
    wire N__38618;
    wire N__38615;
    wire N__38612;
    wire N__38609;
    wire N__38606;
    wire N__38603;
    wire N__38600;
    wire N__38597;
    wire N__38594;
    wire N__38591;
    wire N__38588;
    wire N__38585;
    wire N__38582;
    wire N__38579;
    wire N__38578;
    wire N__38577;
    wire N__38574;
    wire N__38569;
    wire N__38566;
    wire N__38563;
    wire N__38558;
    wire N__38557;
    wire N__38554;
    wire N__38551;
    wire N__38548;
    wire N__38545;
    wire N__38542;
    wire N__38537;
    wire N__38534;
    wire N__38531;
    wire N__38528;
    wire N__38525;
    wire N__38522;
    wire N__38519;
    wire N__38516;
    wire N__38513;
    wire N__38510;
    wire N__38507;
    wire N__38504;
    wire N__38501;
    wire N__38498;
    wire N__38495;
    wire N__38492;
    wire N__38489;
    wire N__38486;
    wire N__38483;
    wire N__38480;
    wire N__38477;
    wire N__38474;
    wire N__38471;
    wire N__38468;
    wire N__38465;
    wire N__38462;
    wire N__38459;
    wire N__38456;
    wire N__38453;
    wire N__38450;
    wire N__38447;
    wire N__38444;
    wire N__38441;
    wire N__38438;
    wire N__38435;
    wire N__38432;
    wire N__38429;
    wire N__38428;
    wire N__38427;
    wire N__38424;
    wire N__38421;
    wire N__38418;
    wire N__38417;
    wire N__38414;
    wire N__38411;
    wire N__38406;
    wire N__38399;
    wire N__38396;
    wire N__38395;
    wire N__38394;
    wire N__38391;
    wire N__38388;
    wire N__38385;
    wire N__38378;
    wire N__38375;
    wire N__38372;
    wire N__38369;
    wire N__38366;
    wire N__38365;
    wire N__38360;
    wire N__38357;
    wire N__38354;
    wire N__38353;
    wire N__38350;
    wire N__38347;
    wire N__38344;
    wire N__38341;
    wire N__38336;
    wire N__38335;
    wire N__38334;
    wire N__38327;
    wire N__38324;
    wire N__38321;
    wire N__38318;
    wire N__38315;
    wire N__38312;
    wire N__38309;
    wire N__38306;
    wire N__38303;
    wire N__38300;
    wire N__38297;
    wire N__38294;
    wire N__38291;
    wire N__38288;
    wire N__38285;
    wire N__38282;
    wire N__38279;
    wire N__38276;
    wire N__38273;
    wire N__38270;
    wire N__38267;
    wire N__38264;
    wire N__38261;
    wire N__38258;
    wire N__38255;
    wire N__38252;
    wire N__38249;
    wire N__38246;
    wire N__38245;
    wire N__38242;
    wire N__38239;
    wire N__38238;
    wire N__38237;
    wire N__38234;
    wire N__38231;
    wire N__38226;
    wire N__38221;
    wire N__38218;
    wire N__38213;
    wire N__38210;
    wire N__38207;
    wire N__38204;
    wire N__38203;
    wire N__38200;
    wire N__38197;
    wire N__38196;
    wire N__38195;
    wire N__38190;
    wire N__38185;
    wire N__38180;
    wire N__38177;
    wire N__38174;
    wire N__38171;
    wire N__38170;
    wire N__38169;
    wire N__38168;
    wire N__38167;
    wire N__38164;
    wire N__38161;
    wire N__38158;
    wire N__38153;
    wire N__38150;
    wire N__38147;
    wire N__38144;
    wire N__38139;
    wire N__38136;
    wire N__38131;
    wire N__38126;
    wire N__38123;
    wire N__38120;
    wire N__38117;
    wire N__38114;
    wire N__38111;
    wire N__38110;
    wire N__38109;
    wire N__38108;
    wire N__38105;
    wire N__38102;
    wire N__38099;
    wire N__38096;
    wire N__38095;
    wire N__38094;
    wire N__38093;
    wire N__38092;
    wire N__38091;
    wire N__38090;
    wire N__38089;
    wire N__38084;
    wire N__38079;
    wire N__38068;
    wire N__38063;
    wire N__38060;
    wire N__38051;
    wire N__38048;
    wire N__38045;
    wire N__38042;
    wire N__38039;
    wire N__38036;
    wire N__38033;
    wire N__38032;
    wire N__38029;
    wire N__38026;
    wire N__38021;
    wire N__38018;
    wire N__38015;
    wire N__38014;
    wire N__38011;
    wire N__38008;
    wire N__38003;
    wire N__38000;
    wire N__37997;
    wire N__37996;
    wire N__37993;
    wire N__37990;
    wire N__37987;
    wire N__37982;
    wire N__37981;
    wire N__37978;
    wire N__37975;
    wire N__37970;
    wire N__37967;
    wire N__37964;
    wire N__37963;
    wire N__37960;
    wire N__37957;
    wire N__37954;
    wire N__37949;
    wire N__37948;
    wire N__37943;
    wire N__37940;
    wire N__37937;
    wire N__37934;
    wire N__37931;
    wire N__37928;
    wire N__37925;
    wire N__37922;
    wire N__37919;
    wire N__37916;
    wire N__37913;
    wire N__37910;
    wire N__37907;
    wire N__37904;
    wire N__37903;
    wire N__37902;
    wire N__37899;
    wire N__37896;
    wire N__37893;
    wire N__37890;
    wire N__37889;
    wire N__37884;
    wire N__37881;
    wire N__37878;
    wire N__37875;
    wire N__37868;
    wire N__37865;
    wire N__37862;
    wire N__37859;
    wire N__37856;
    wire N__37853;
    wire N__37850;
    wire N__37847;
    wire N__37844;
    wire N__37841;
    wire N__37838;
    wire N__37835;
    wire N__37832;
    wire N__37829;
    wire N__37826;
    wire N__37823;
    wire N__37820;
    wire N__37817;
    wire N__37816;
    wire N__37815;
    wire N__37812;
    wire N__37809;
    wire N__37806;
    wire N__37799;
    wire N__37798;
    wire N__37797;
    wire N__37794;
    wire N__37793;
    wire N__37790;
    wire N__37787;
    wire N__37784;
    wire N__37781;
    wire N__37772;
    wire N__37771;
    wire N__37770;
    wire N__37769;
    wire N__37766;
    wire N__37763;
    wire N__37760;
    wire N__37757;
    wire N__37754;
    wire N__37745;
    wire N__37744;
    wire N__37743;
    wire N__37742;
    wire N__37739;
    wire N__37736;
    wire N__37733;
    wire N__37730;
    wire N__37721;
    wire N__37720;
    wire N__37717;
    wire N__37716;
    wire N__37713;
    wire N__37710;
    wire N__37707;
    wire N__37704;
    wire N__37697;
    wire N__37694;
    wire N__37691;
    wire N__37688;
    wire N__37687;
    wire N__37686;
    wire N__37683;
    wire N__37678;
    wire N__37673;
    wire N__37670;
    wire N__37667;
    wire N__37664;
    wire N__37661;
    wire N__37658;
    wire N__37657;
    wire N__37654;
    wire N__37651;
    wire N__37646;
    wire N__37643;
    wire N__37640;
    wire N__37637;
    wire N__37634;
    wire N__37631;
    wire N__37628;
    wire N__37625;
    wire N__37622;
    wire N__37619;
    wire N__37616;
    wire N__37613;
    wire N__37610;
    wire N__37607;
    wire N__37604;
    wire N__37601;
    wire N__37600;
    wire N__37599;
    wire N__37596;
    wire N__37591;
    wire N__37586;
    wire N__37585;
    wire N__37582;
    wire N__37579;
    wire N__37576;
    wire N__37573;
    wire N__37568;
    wire N__37565;
    wire N__37562;
    wire N__37559;
    wire N__37556;
    wire N__37553;
    wire N__37552;
    wire N__37551;
    wire N__37548;
    wire N__37547;
    wire N__37544;
    wire N__37543;
    wire N__37542;
    wire N__37539;
    wire N__37536;
    wire N__37527;
    wire N__37520;
    wire N__37519;
    wire N__37518;
    wire N__37515;
    wire N__37512;
    wire N__37509;
    wire N__37506;
    wire N__37501;
    wire N__37496;
    wire N__37493;
    wire N__37490;
    wire N__37487;
    wire N__37484;
    wire N__37481;
    wire N__37478;
    wire N__37475;
    wire N__37472;
    wire N__37469;
    wire N__37466;
    wire N__37463;
    wire N__37460;
    wire N__37459;
    wire N__37456;
    wire N__37453;
    wire N__37452;
    wire N__37451;
    wire N__37448;
    wire N__37443;
    wire N__37440;
    wire N__37433;
    wire N__37430;
    wire N__37427;
    wire N__37424;
    wire N__37423;
    wire N__37420;
    wire N__37419;
    wire N__37418;
    wire N__37415;
    wire N__37412;
    wire N__37409;
    wire N__37406;
    wire N__37397;
    wire N__37394;
    wire N__37393;
    wire N__37392;
    wire N__37389;
    wire N__37386;
    wire N__37383;
    wire N__37380;
    wire N__37377;
    wire N__37374;
    wire N__37367;
    wire N__37364;
    wire N__37361;
    wire N__37358;
    wire N__37355;
    wire N__37352;
    wire N__37349;
    wire N__37346;
    wire N__37343;
    wire N__37340;
    wire N__37337;
    wire N__37334;
    wire N__37331;
    wire N__37328;
    wire N__37325;
    wire N__37322;
    wire N__37319;
    wire N__37316;
    wire N__37313;
    wire N__37310;
    wire N__37307;
    wire N__37304;
    wire N__37301;
    wire N__37298;
    wire N__37295;
    wire N__37292;
    wire N__37289;
    wire N__37286;
    wire N__37283;
    wire N__37280;
    wire N__37277;
    wire N__37274;
    wire N__37271;
    wire N__37268;
    wire N__37265;
    wire N__37262;
    wire N__37259;
    wire N__37256;
    wire N__37253;
    wire N__37252;
    wire N__37247;
    wire N__37244;
    wire N__37243;
    wire N__37240;
    wire N__37237;
    wire N__37234;
    wire N__37229;
    wire N__37226;
    wire N__37225;
    wire N__37222;
    wire N__37219;
    wire N__37218;
    wire N__37215;
    wire N__37212;
    wire N__37209;
    wire N__37202;
    wire N__37201;
    wire N__37200;
    wire N__37195;
    wire N__37192;
    wire N__37189;
    wire N__37186;
    wire N__37183;
    wire N__37178;
    wire N__37177;
    wire N__37176;
    wire N__37175;
    wire N__37174;
    wire N__37163;
    wire N__37160;
    wire N__37157;
    wire N__37156;
    wire N__37155;
    wire N__37154;
    wire N__37153;
    wire N__37148;
    wire N__37147;
    wire N__37146;
    wire N__37145;
    wire N__37144;
    wire N__37143;
    wire N__37142;
    wire N__37141;
    wire N__37138;
    wire N__37135;
    wire N__37132;
    wire N__37131;
    wire N__37128;
    wire N__37125;
    wire N__37122;
    wire N__37119;
    wire N__37116;
    wire N__37107;
    wire N__37106;
    wire N__37105;
    wire N__37104;
    wire N__37103;
    wire N__37102;
    wire N__37099;
    wire N__37096;
    wire N__37093;
    wire N__37090;
    wire N__37079;
    wire N__37078;
    wire N__37077;
    wire N__37076;
    wire N__37075;
    wire N__37072;
    wire N__37069;
    wire N__37066;
    wire N__37061;
    wire N__37058;
    wire N__37049;
    wire N__37040;
    wire N__37025;
    wire N__37022;
    wire N__37019;
    wire N__37018;
    wire N__37015;
    wire N__37012;
    wire N__37009;
    wire N__37006;
    wire N__37001;
    wire N__37000;
    wire N__36999;
    wire N__36998;
    wire N__36997;
    wire N__36996;
    wire N__36995;
    wire N__36994;
    wire N__36991;
    wire N__36988;
    wire N__36985;
    wire N__36984;
    wire N__36983;
    wire N__36982;
    wire N__36981;
    wire N__36980;
    wire N__36975;
    wire N__36974;
    wire N__36971;
    wire N__36970;
    wire N__36969;
    wire N__36966;
    wire N__36963;
    wire N__36962;
    wire N__36961;
    wire N__36958;
    wire N__36953;
    wire N__36948;
    wire N__36945;
    wire N__36944;
    wire N__36941;
    wire N__36938;
    wire N__36935;
    wire N__36934;
    wire N__36929;
    wire N__36926;
    wire N__36921;
    wire N__36918;
    wire N__36913;
    wire N__36906;
    wire N__36903;
    wire N__36900;
    wire N__36899;
    wire N__36898;
    wire N__36897;
    wire N__36896;
    wire N__36895;
    wire N__36892;
    wire N__36887;
    wire N__36884;
    wire N__36869;
    wire N__36868;
    wire N__36867;
    wire N__36866;
    wire N__36865;
    wire N__36864;
    wire N__36861;
    wire N__36856;
    wire N__36849;
    wire N__36840;
    wire N__36829;
    wire N__36826;
    wire N__36815;
    wire N__36812;
    wire N__36809;
    wire N__36808;
    wire N__36805;
    wire N__36802;
    wire N__36799;
    wire N__36794;
    wire N__36791;
    wire N__36788;
    wire N__36785;
    wire N__36782;
    wire N__36779;
    wire N__36776;
    wire N__36773;
    wire N__36770;
    wire N__36767;
    wire N__36764;
    wire N__36761;
    wire N__36758;
    wire N__36755;
    wire N__36752;
    wire N__36749;
    wire N__36746;
    wire N__36743;
    wire N__36740;
    wire N__36737;
    wire N__36734;
    wire N__36731;
    wire N__36728;
    wire N__36725;
    wire N__36722;
    wire N__36719;
    wire N__36716;
    wire N__36713;
    wire N__36710;
    wire N__36707;
    wire N__36704;
    wire N__36701;
    wire N__36698;
    wire N__36695;
    wire N__36692;
    wire N__36689;
    wire N__36686;
    wire N__36683;
    wire N__36680;
    wire N__36677;
    wire N__36674;
    wire N__36671;
    wire N__36668;
    wire N__36665;
    wire N__36664;
    wire N__36661;
    wire N__36658;
    wire N__36653;
    wire N__36650;
    wire N__36647;
    wire N__36644;
    wire N__36641;
    wire N__36638;
    wire N__36637;
    wire N__36634;
    wire N__36631;
    wire N__36628;
    wire N__36623;
    wire N__36620;
    wire N__36617;
    wire N__36614;
    wire N__36611;
    wire N__36608;
    wire N__36605;
    wire N__36602;
    wire N__36599;
    wire N__36596;
    wire N__36593;
    wire N__36590;
    wire N__36587;
    wire N__36584;
    wire N__36581;
    wire N__36578;
    wire N__36575;
    wire N__36572;
    wire N__36569;
    wire N__36566;
    wire N__36563;
    wire N__36560;
    wire N__36557;
    wire N__36554;
    wire N__36551;
    wire N__36548;
    wire N__36545;
    wire N__36542;
    wire N__36539;
    wire N__36536;
    wire N__36533;
    wire N__36530;
    wire N__36527;
    wire N__36524;
    wire N__36521;
    wire N__36518;
    wire N__36515;
    wire N__36512;
    wire N__36509;
    wire N__36506;
    wire N__36503;
    wire N__36500;
    wire N__36497;
    wire N__36494;
    wire N__36491;
    wire N__36488;
    wire N__36485;
    wire N__36482;
    wire N__36479;
    wire N__36476;
    wire N__36473;
    wire N__36470;
    wire N__36467;
    wire N__36464;
    wire N__36461;
    wire N__36458;
    wire N__36455;
    wire N__36452;
    wire N__36449;
    wire N__36446;
    wire N__36443;
    wire N__36440;
    wire N__36437;
    wire N__36434;
    wire N__36431;
    wire N__36428;
    wire N__36425;
    wire N__36422;
    wire N__36419;
    wire N__36416;
    wire N__36413;
    wire N__36410;
    wire N__36407;
    wire N__36404;
    wire N__36401;
    wire N__36398;
    wire N__36395;
    wire N__36392;
    wire N__36391;
    wire N__36388;
    wire N__36385;
    wire N__36382;
    wire N__36377;
    wire N__36374;
    wire N__36373;
    wire N__36370;
    wire N__36367;
    wire N__36364;
    wire N__36359;
    wire N__36356;
    wire N__36355;
    wire N__36352;
    wire N__36349;
    wire N__36346;
    wire N__36341;
    wire N__36338;
    wire N__36335;
    wire N__36334;
    wire N__36331;
    wire N__36328;
    wire N__36325;
    wire N__36320;
    wire N__36317;
    wire N__36314;
    wire N__36311;
    wire N__36308;
    wire N__36305;
    wire N__36302;
    wire N__36301;
    wire N__36300;
    wire N__36297;
    wire N__36294;
    wire N__36293;
    wire N__36290;
    wire N__36285;
    wire N__36284;
    wire N__36281;
    wire N__36280;
    wire N__36279;
    wire N__36276;
    wire N__36273;
    wire N__36270;
    wire N__36263;
    wire N__36254;
    wire N__36253;
    wire N__36252;
    wire N__36251;
    wire N__36248;
    wire N__36245;
    wire N__36242;
    wire N__36241;
    wire N__36240;
    wire N__36239;
    wire N__36236;
    wire N__36233;
    wire N__36228;
    wire N__36221;
    wire N__36220;
    wire N__36217;
    wire N__36214;
    wire N__36209;
    wire N__36206;
    wire N__36203;
    wire N__36198;
    wire N__36191;
    wire N__36190;
    wire N__36189;
    wire N__36186;
    wire N__36181;
    wire N__36180;
    wire N__36177;
    wire N__36174;
    wire N__36171;
    wire N__36166;
    wire N__36161;
    wire N__36158;
    wire N__36157;
    wire N__36154;
    wire N__36151;
    wire N__36146;
    wire N__36143;
    wire N__36140;
    wire N__36137;
    wire N__36134;
    wire N__36131;
    wire N__36128;
    wire N__36125;
    wire N__36122;
    wire N__36119;
    wire N__36116;
    wire N__36113;
    wire N__36110;
    wire N__36109;
    wire N__36106;
    wire N__36103;
    wire N__36100;
    wire N__36095;
    wire N__36092;
    wire N__36091;
    wire N__36088;
    wire N__36085;
    wire N__36082;
    wire N__36077;
    wire N__36074;
    wire N__36073;
    wire N__36070;
    wire N__36067;
    wire N__36064;
    wire N__36059;
    wire N__36056;
    wire N__36055;
    wire N__36052;
    wire N__36049;
    wire N__36046;
    wire N__36041;
    wire N__36038;
    wire N__36037;
    wire N__36034;
    wire N__36031;
    wire N__36028;
    wire N__36023;
    wire N__36020;
    wire N__36019;
    wire N__36016;
    wire N__36013;
    wire N__36010;
    wire N__36005;
    wire N__36002;
    wire N__35999;
    wire N__35998;
    wire N__35995;
    wire N__35992;
    wire N__35989;
    wire N__35984;
    wire N__35981;
    wire N__35980;
    wire N__35977;
    wire N__35974;
    wire N__35971;
    wire N__35966;
    wire N__35963;
    wire N__35960;
    wire N__35959;
    wire N__35956;
    wire N__35953;
    wire N__35950;
    wire N__35945;
    wire N__35942;
    wire N__35939;
    wire N__35936;
    wire N__35933;
    wire N__35930;
    wire N__35929;
    wire N__35928;
    wire N__35927;
    wire N__35926;
    wire N__35923;
    wire N__35922;
    wire N__35919;
    wire N__35918;
    wire N__35917;
    wire N__35914;
    wire N__35911;
    wire N__35908;
    wire N__35905;
    wire N__35902;
    wire N__35899;
    wire N__35894;
    wire N__35891;
    wire N__35886;
    wire N__35883;
    wire N__35880;
    wire N__35877;
    wire N__35874;
    wire N__35867;
    wire N__35862;
    wire N__35855;
    wire N__35852;
    wire N__35849;
    wire N__35846;
    wire N__35845;
    wire N__35844;
    wire N__35843;
    wire N__35840;
    wire N__35837;
    wire N__35834;
    wire N__35831;
    wire N__35822;
    wire N__35821;
    wire N__35820;
    wire N__35817;
    wire N__35816;
    wire N__35815;
    wire N__35810;
    wire N__35807;
    wire N__35804;
    wire N__35801;
    wire N__35798;
    wire N__35795;
    wire N__35792;
    wire N__35785;
    wire N__35780;
    wire N__35777;
    wire N__35774;
    wire N__35771;
    wire N__35768;
    wire N__35765;
    wire N__35762;
    wire N__35759;
    wire N__35756;
    wire N__35755;
    wire N__35752;
    wire N__35749;
    wire N__35746;
    wire N__35743;
    wire N__35742;
    wire N__35739;
    wire N__35736;
    wire N__35733;
    wire N__35728;
    wire N__35725;
    wire N__35722;
    wire N__35717;
    wire N__35716;
    wire N__35713;
    wire N__35710;
    wire N__35707;
    wire N__35702;
    wire N__35699;
    wire N__35696;
    wire N__35693;
    wire N__35690;
    wire N__35687;
    wire N__35686;
    wire N__35683;
    wire N__35680;
    wire N__35677;
    wire N__35672;
    wire N__35669;
    wire N__35668;
    wire N__35665;
    wire N__35662;
    wire N__35659;
    wire N__35654;
    wire N__35651;
    wire N__35650;
    wire N__35647;
    wire N__35644;
    wire N__35641;
    wire N__35636;
    wire N__35633;
    wire N__35632;
    wire N__35629;
    wire N__35626;
    wire N__35623;
    wire N__35618;
    wire N__35615;
    wire N__35612;
    wire N__35609;
    wire N__35606;
    wire N__35603;
    wire N__35600;
    wire N__35597;
    wire N__35594;
    wire N__35591;
    wire N__35588;
    wire N__35585;
    wire N__35582;
    wire N__35579;
    wire N__35576;
    wire N__35573;
    wire N__35570;
    wire N__35567;
    wire N__35564;
    wire N__35561;
    wire N__35558;
    wire N__35555;
    wire N__35552;
    wire N__35549;
    wire N__35546;
    wire N__35543;
    wire N__35540;
    wire N__35539;
    wire N__35536;
    wire N__35533;
    wire N__35528;
    wire N__35525;
    wire N__35522;
    wire N__35519;
    wire N__35516;
    wire N__35513;
    wire N__35510;
    wire N__35507;
    wire N__35504;
    wire N__35501;
    wire N__35498;
    wire N__35495;
    wire N__35492;
    wire N__35489;
    wire N__35486;
    wire N__35483;
    wire N__35480;
    wire N__35477;
    wire N__35474;
    wire N__35471;
    wire N__35468;
    wire N__35465;
    wire N__35462;
    wire N__35459;
    wire N__35456;
    wire N__35453;
    wire N__35450;
    wire N__35447;
    wire N__35446;
    wire N__35443;
    wire N__35440;
    wire N__35435;
    wire N__35432;
    wire N__35429;
    wire N__35426;
    wire N__35425;
    wire N__35422;
    wire N__35419;
    wire N__35414;
    wire N__35413;
    wire N__35408;
    wire N__35405;
    wire N__35402;
    wire N__35399;
    wire N__35398;
    wire N__35395;
    wire N__35392;
    wire N__35387;
    wire N__35386;
    wire N__35383;
    wire N__35382;
    wire N__35379;
    wire N__35376;
    wire N__35373;
    wire N__35370;
    wire N__35363;
    wire N__35360;
    wire N__35357;
    wire N__35356;
    wire N__35353;
    wire N__35350;
    wire N__35347;
    wire N__35344;
    wire N__35339;
    wire N__35336;
    wire N__35335;
    wire N__35332;
    wire N__35329;
    wire N__35326;
    wire N__35323;
    wire N__35318;
    wire N__35315;
    wire N__35312;
    wire N__35309;
    wire N__35306;
    wire N__35303;
    wire N__35300;
    wire N__35297;
    wire N__35294;
    wire N__35291;
    wire N__35288;
    wire N__35285;
    wire N__35282;
    wire N__35279;
    wire N__35278;
    wire N__35275;
    wire N__35272;
    wire N__35267;
    wire N__35264;
    wire N__35261;
    wire N__35258;
    wire N__35257;
    wire N__35254;
    wire N__35251;
    wire N__35246;
    wire N__35243;
    wire N__35240;
    wire N__35239;
    wire N__35236;
    wire N__35233;
    wire N__35228;
    wire N__35225;
    wire N__35222;
    wire N__35221;
    wire N__35218;
    wire N__35215;
    wire N__35210;
    wire N__35207;
    wire N__35204;
    wire N__35201;
    wire N__35200;
    wire N__35197;
    wire N__35194;
    wire N__35193;
    wire N__35192;
    wire N__35189;
    wire N__35186;
    wire N__35181;
    wire N__35174;
    wire N__35171;
    wire N__35168;
    wire N__35165;
    wire N__35164;
    wire N__35161;
    wire N__35158;
    wire N__35153;
    wire N__35150;
    wire N__35147;
    wire N__35146;
    wire N__35143;
    wire N__35140;
    wire N__35135;
    wire N__35132;
    wire N__35129;
    wire N__35126;
    wire N__35123;
    wire N__35120;
    wire N__35119;
    wire N__35116;
    wire N__35113;
    wire N__35108;
    wire N__35107;
    wire N__35104;
    wire N__35103;
    wire N__35100;
    wire N__35097;
    wire N__35094;
    wire N__35091;
    wire N__35088;
    wire N__35083;
    wire N__35078;
    wire N__35075;
    wire N__35072;
    wire N__35069;
    wire N__35066;
    wire N__35063;
    wire N__35060;
    wire N__35057;
    wire N__35054;
    wire N__35051;
    wire N__35048;
    wire N__35045;
    wire N__35042;
    wire N__35039;
    wire N__35036;
    wire N__35033;
    wire N__35030;
    wire N__35027;
    wire N__35024;
    wire N__35021;
    wire N__35018;
    wire N__35015;
    wire N__35012;
    wire N__35009;
    wire N__35006;
    wire N__35003;
    wire N__35000;
    wire N__34997;
    wire N__34994;
    wire N__34991;
    wire N__34988;
    wire N__34985;
    wire N__34982;
    wire N__34979;
    wire N__34976;
    wire N__34973;
    wire N__34970;
    wire N__34967;
    wire N__34964;
    wire N__34963;
    wire N__34960;
    wire N__34957;
    wire N__34954;
    wire N__34951;
    wire N__34946;
    wire N__34943;
    wire N__34940;
    wire N__34937;
    wire N__34934;
    wire N__34931;
    wire N__34928;
    wire N__34925;
    wire N__34922;
    wire N__34919;
    wire N__34916;
    wire N__34913;
    wire N__34910;
    wire N__34907;
    wire N__34904;
    wire N__34901;
    wire N__34898;
    wire N__34895;
    wire N__34892;
    wire N__34889;
    wire N__34886;
    wire N__34883;
    wire N__34880;
    wire N__34877;
    wire N__34874;
    wire N__34871;
    wire N__34868;
    wire N__34865;
    wire N__34862;
    wire N__34859;
    wire N__34856;
    wire N__34853;
    wire N__34850;
    wire N__34847;
    wire N__34844;
    wire N__34841;
    wire N__34838;
    wire N__34835;
    wire N__34832;
    wire N__34829;
    wire N__34828;
    wire N__34827;
    wire N__34822;
    wire N__34819;
    wire N__34816;
    wire N__34813;
    wire N__34812;
    wire N__34809;
    wire N__34806;
    wire N__34803;
    wire N__34802;
    wire N__34801;
    wire N__34798;
    wire N__34793;
    wire N__34790;
    wire N__34787;
    wire N__34778;
    wire N__34775;
    wire N__34772;
    wire N__34769;
    wire N__34768;
    wire N__34765;
    wire N__34762;
    wire N__34761;
    wire N__34756;
    wire N__34753;
    wire N__34750;
    wire N__34745;
    wire N__34742;
    wire N__34739;
    wire N__34736;
    wire N__34735;
    wire N__34734;
    wire N__34731;
    wire N__34726;
    wire N__34721;
    wire N__34720;
    wire N__34719;
    wire N__34718;
    wire N__34717;
    wire N__34716;
    wire N__34709;
    wire N__34702;
    wire N__34697;
    wire N__34696;
    wire N__34693;
    wire N__34690;
    wire N__34687;
    wire N__34682;
    wire N__34681;
    wire N__34680;
    wire N__34679;
    wire N__34678;
    wire N__34677;
    wire N__34672;
    wire N__34669;
    wire N__34664;
    wire N__34661;
    wire N__34660;
    wire N__34657;
    wire N__34656;
    wire N__34651;
    wire N__34646;
    wire N__34643;
    wire N__34640;
    wire N__34637;
    wire N__34632;
    wire N__34625;
    wire N__34622;
    wire N__34619;
    wire N__34616;
    wire N__34613;
    wire N__34612;
    wire N__34609;
    wire N__34606;
    wire N__34601;
    wire N__34598;
    wire N__34595;
    wire N__34592;
    wire N__34589;
    wire N__34586;
    wire N__34585;
    wire N__34584;
    wire N__34581;
    wire N__34576;
    wire N__34571;
    wire N__34568;
    wire N__34565;
    wire N__34562;
    wire N__34561;
    wire N__34558;
    wire N__34555;
    wire N__34552;
    wire N__34547;
    wire N__34544;
    wire N__34541;
    wire N__34538;
    wire N__34535;
    wire N__34534;
    wire N__34531;
    wire N__34528;
    wire N__34523;
    wire N__34520;
    wire N__34517;
    wire N__34514;
    wire N__34511;
    wire N__34510;
    wire N__34509;
    wire N__34502;
    wire N__34499;
    wire N__34498;
    wire N__34495;
    wire N__34490;
    wire N__34487;
    wire N__34484;
    wire N__34483;
    wire N__34478;
    wire N__34475;
    wire N__34474;
    wire N__34473;
    wire N__34468;
    wire N__34465;
    wire N__34462;
    wire N__34457;
    wire N__34454;
    wire N__34451;
    wire N__34448;
    wire N__34447;
    wire N__34446;
    wire N__34443;
    wire N__34440;
    wire N__34435;
    wire N__34432;
    wire N__34429;
    wire N__34424;
    wire N__34423;
    wire N__34420;
    wire N__34417;
    wire N__34414;
    wire N__34411;
    wire N__34406;
    wire N__34405;
    wire N__34404;
    wire N__34401;
    wire N__34396;
    wire N__34393;
    wire N__34390;
    wire N__34385;
    wire N__34384;
    wire N__34381;
    wire N__34378;
    wire N__34373;
    wire N__34370;
    wire N__34367;
    wire N__34366;
    wire N__34363;
    wire N__34360;
    wire N__34357;
    wire N__34352;
    wire N__34351;
    wire N__34348;
    wire N__34345;
    wire N__34342;
    wire N__34339;
    wire N__34338;
    wire N__34335;
    wire N__34332;
    wire N__34329;
    wire N__34326;
    wire N__34319;
    wire N__34318;
    wire N__34317;
    wire N__34312;
    wire N__34309;
    wire N__34304;
    wire N__34303;
    wire N__34302;
    wire N__34301;
    wire N__34300;
    wire N__34299;
    wire N__34286;
    wire N__34283;
    wire N__34280;
    wire N__34277;
    wire N__34274;
    wire N__34271;
    wire N__34270;
    wire N__34267;
    wire N__34264;
    wire N__34259;
    wire N__34256;
    wire N__34253;
    wire N__34252;
    wire N__34249;
    wire N__34246;
    wire N__34243;
    wire N__34238;
    wire N__34235;
    wire N__34232;
    wire N__34231;
    wire N__34230;
    wire N__34225;
    wire N__34222;
    wire N__34217;
    wire N__34214;
    wire N__34211;
    wire N__34208;
    wire N__34207;
    wire N__34202;
    wire N__34201;
    wire N__34198;
    wire N__34195;
    wire N__34192;
    wire N__34187;
    wire N__34184;
    wire N__34181;
    wire N__34178;
    wire N__34175;
    wire N__34172;
    wire N__34169;
    wire N__34166;
    wire N__34163;
    wire N__34160;
    wire N__34159;
    wire N__34156;
    wire N__34153;
    wire N__34148;
    wire N__34147;
    wire N__34146;
    wire N__34143;
    wire N__34140;
    wire N__34137;
    wire N__34134;
    wire N__34131;
    wire N__34128;
    wire N__34125;
    wire N__34122;
    wire N__34119;
    wire N__34116;
    wire N__34113;
    wire N__34110;
    wire N__34107;
    wire N__34102;
    wire N__34099;
    wire N__34096;
    wire N__34091;
    wire N__34088;
    wire N__34085;
    wire N__34082;
    wire N__34079;
    wire N__34076;
    wire N__34073;
    wire N__34070;
    wire N__34067;
    wire N__34064;
    wire N__34063;
    wire N__34060;
    wire N__34059;
    wire N__34056;
    wire N__34053;
    wire N__34050;
    wire N__34043;
    wire N__34040;
    wire N__34037;
    wire N__34036;
    wire N__34033;
    wire N__34030;
    wire N__34029;
    wire N__34028;
    wire N__34027;
    wire N__34026;
    wire N__34021;
    wire N__34018;
    wire N__34013;
    wire N__34010;
    wire N__34001;
    wire N__34000;
    wire N__33997;
    wire N__33996;
    wire N__33993;
    wire N__33988;
    wire N__33985;
    wire N__33982;
    wire N__33979;
    wire N__33976;
    wire N__33973;
    wire N__33970;
    wire N__33967;
    wire N__33962;
    wire N__33959;
    wire N__33956;
    wire N__33953;
    wire N__33950;
    wire N__33947;
    wire N__33944;
    wire N__33941;
    wire N__33940;
    wire N__33939;
    wire N__33936;
    wire N__33933;
    wire N__33930;
    wire N__33929;
    wire N__33926;
    wire N__33923;
    wire N__33920;
    wire N__33917;
    wire N__33914;
    wire N__33905;
    wire N__33902;
    wire N__33899;
    wire N__33898;
    wire N__33895;
    wire N__33892;
    wire N__33891;
    wire N__33888;
    wire N__33883;
    wire N__33878;
    wire N__33875;
    wire N__33872;
    wire N__33869;
    wire N__33866;
    wire N__33863;
    wire N__33860;
    wire N__33857;
    wire N__33854;
    wire N__33851;
    wire N__33848;
    wire N__33847;
    wire N__33844;
    wire N__33841;
    wire N__33840;
    wire N__33837;
    wire N__33834;
    wire N__33831;
    wire N__33828;
    wire N__33821;
    wire N__33820;
    wire N__33819;
    wire N__33816;
    wire N__33815;
    wire N__33810;
    wire N__33807;
    wire N__33804;
    wire N__33797;
    wire N__33794;
    wire N__33791;
    wire N__33788;
    wire N__33785;
    wire N__33782;
    wire N__33779;
    wire N__33776;
    wire N__33775;
    wire N__33774;
    wire N__33773;
    wire N__33770;
    wire N__33767;
    wire N__33766;
    wire N__33765;
    wire N__33764;
    wire N__33763;
    wire N__33762;
    wire N__33761;
    wire N__33760;
    wire N__33759;
    wire N__33758;
    wire N__33757;
    wire N__33756;
    wire N__33755;
    wire N__33752;
    wire N__33749;
    wire N__33746;
    wire N__33745;
    wire N__33744;
    wire N__33743;
    wire N__33742;
    wire N__33741;
    wire N__33738;
    wire N__33735;
    wire N__33728;
    wire N__33727;
    wire N__33726;
    wire N__33725;
    wire N__33722;
    wire N__33719;
    wire N__33718;
    wire N__33717;
    wire N__33716;
    wire N__33713;
    wire N__33712;
    wire N__33709;
    wire N__33708;
    wire N__33707;
    wire N__33704;
    wire N__33703;
    wire N__33702;
    wire N__33699;
    wire N__33696;
    wire N__33695;
    wire N__33694;
    wire N__33693;
    wire N__33692;
    wire N__33691;
    wire N__33688;
    wire N__33685;
    wire N__33680;
    wire N__33679;
    wire N__33678;
    wire N__33677;
    wire N__33676;
    wire N__33673;
    wire N__33672;
    wire N__33671;
    wire N__33670;
    wire N__33669;
    wire N__33666;
    wire N__33661;
    wire N__33658;
    wire N__33651;
    wire N__33644;
    wire N__33631;
    wire N__33616;
    wire N__33603;
    wire N__33602;
    wire N__33601;
    wire N__33600;
    wire N__33599;
    wire N__33598;
    wire N__33597;
    wire N__33594;
    wire N__33587;
    wire N__33584;
    wire N__33579;
    wire N__33566;
    wire N__33561;
    wire N__33548;
    wire N__33545;
    wire N__33534;
    wire N__33529;
    wire N__33526;
    wire N__33523;
    wire N__33516;
    wire N__33503;
    wire N__33502;
    wire N__33501;
    wire N__33498;
    wire N__33495;
    wire N__33490;
    wire N__33485;
    wire N__33482;
    wire N__33479;
    wire N__33476;
    wire N__33473;
    wire N__33470;
    wire N__33467;
    wire N__33464;
    wire N__33463;
    wire N__33462;
    wire N__33457;
    wire N__33454;
    wire N__33451;
    wire N__33446;
    wire N__33443;
    wire N__33442;
    wire N__33439;
    wire N__33436;
    wire N__33433;
    wire N__33428;
    wire N__33425;
    wire N__33424;
    wire N__33421;
    wire N__33418;
    wire N__33415;
    wire N__33410;
    wire N__33407;
    wire N__33406;
    wire N__33403;
    wire N__33400;
    wire N__33399;
    wire N__33394;
    wire N__33391;
    wire N__33388;
    wire N__33383;
    wire N__33380;
    wire N__33377;
    wire N__33376;
    wire N__33373;
    wire N__33370;
    wire N__33367;
    wire N__33366;
    wire N__33361;
    wire N__33360;
    wire N__33357;
    wire N__33354;
    wire N__33351;
    wire N__33348;
    wire N__33345;
    wire N__33338;
    wire N__33337;
    wire N__33336;
    wire N__33335;
    wire N__33332;
    wire N__33329;
    wire N__33326;
    wire N__33323;
    wire N__33320;
    wire N__33317;
    wire N__33314;
    wire N__33311;
    wire N__33308;
    wire N__33305;
    wire N__33302;
    wire N__33293;
    wire N__33290;
    wire N__33287;
    wire N__33284;
    wire N__33281;
    wire N__33280;
    wire N__33279;
    wire N__33274;
    wire N__33271;
    wire N__33268;
    wire N__33263;
    wire N__33260;
    wire N__33259;
    wire N__33258;
    wire N__33253;
    wire N__33250;
    wire N__33247;
    wire N__33242;
    wire N__33239;
    wire N__33238;
    wire N__33235;
    wire N__33232;
    wire N__33231;
    wire N__33226;
    wire N__33223;
    wire N__33220;
    wire N__33215;
    wire N__33212;
    wire N__33211;
    wire N__33208;
    wire N__33205;
    wire N__33204;
    wire N__33199;
    wire N__33196;
    wire N__33193;
    wire N__33188;
    wire N__33185;
    wire N__33184;
    wire N__33179;
    wire N__33178;
    wire N__33175;
    wire N__33172;
    wire N__33169;
    wire N__33164;
    wire N__33161;
    wire N__33158;
    wire N__33157;
    wire N__33154;
    wire N__33151;
    wire N__33150;
    wire N__33145;
    wire N__33142;
    wire N__33139;
    wire N__33134;
    wire N__33131;
    wire N__33130;
    wire N__33127;
    wire N__33124;
    wire N__33121;
    wire N__33118;
    wire N__33117;
    wire N__33112;
    wire N__33109;
    wire N__33106;
    wire N__33101;
    wire N__33098;
    wire N__33095;
    wire N__33094;
    wire N__33093;
    wire N__33090;
    wire N__33087;
    wire N__33084;
    wire N__33079;
    wire N__33074;
    wire N__33071;
    wire N__33068;
    wire N__33067;
    wire N__33062;
    wire N__33061;
    wire N__33058;
    wire N__33055;
    wire N__33052;
    wire N__33047;
    wire N__33044;
    wire N__33043;
    wire N__33038;
    wire N__33037;
    wire N__33034;
    wire N__33031;
    wire N__33028;
    wire N__33023;
    wire N__33020;
    wire N__33019;
    wire N__33016;
    wire N__33013;
    wire N__33012;
    wire N__33007;
    wire N__33004;
    wire N__33001;
    wire N__32996;
    wire N__32993;
    wire N__32992;
    wire N__32989;
    wire N__32986;
    wire N__32985;
    wire N__32980;
    wire N__32977;
    wire N__32974;
    wire N__32969;
    wire N__32966;
    wire N__32965;
    wire N__32960;
    wire N__32959;
    wire N__32956;
    wire N__32953;
    wire N__32950;
    wire N__32945;
    wire N__32942;
    wire N__32939;
    wire N__32938;
    wire N__32935;
    wire N__32932;
    wire N__32931;
    wire N__32926;
    wire N__32923;
    wire N__32920;
    wire N__32915;
    wire N__32912;
    wire N__32909;
    wire N__32908;
    wire N__32905;
    wire N__32902;
    wire N__32901;
    wire N__32898;
    wire N__32895;
    wire N__32892;
    wire N__32887;
    wire N__32882;
    wire N__32879;
    wire N__32876;
    wire N__32873;
    wire N__32872;
    wire N__32871;
    wire N__32868;
    wire N__32865;
    wire N__32862;
    wire N__32857;
    wire N__32852;
    wire N__32849;
    wire N__32846;
    wire N__32845;
    wire N__32842;
    wire N__32839;
    wire N__32836;
    wire N__32835;
    wire N__32830;
    wire N__32827;
    wire N__32824;
    wire N__32819;
    wire N__32816;
    wire N__32815;
    wire N__32810;
    wire N__32809;
    wire N__32806;
    wire N__32803;
    wire N__32800;
    wire N__32795;
    wire N__32792;
    wire N__32791;
    wire N__32788;
    wire N__32785;
    wire N__32784;
    wire N__32779;
    wire N__32776;
    wire N__32773;
    wire N__32768;
    wire N__32765;
    wire N__32764;
    wire N__32761;
    wire N__32760;
    wire N__32757;
    wire N__32754;
    wire N__32751;
    wire N__32746;
    wire N__32741;
    wire N__32738;
    wire N__32737;
    wire N__32732;
    wire N__32731;
    wire N__32728;
    wire N__32725;
    wire N__32722;
    wire N__32717;
    wire N__32714;
    wire N__32713;
    wire N__32710;
    wire N__32707;
    wire N__32702;
    wire N__32701;
    wire N__32698;
    wire N__32695;
    wire N__32692;
    wire N__32687;
    wire N__32684;
    wire N__32681;
    wire N__32680;
    wire N__32677;
    wire N__32674;
    wire N__32673;
    wire N__32670;
    wire N__32667;
    wire N__32664;
    wire N__32659;
    wire N__32654;
    wire N__32651;
    wire N__32648;
    wire N__32645;
    wire N__32644;
    wire N__32643;
    wire N__32640;
    wire N__32637;
    wire N__32634;
    wire N__32629;
    wire N__32624;
    wire N__32621;
    wire N__32618;
    wire N__32615;
    wire N__32612;
    wire N__32609;
    wire N__32606;
    wire N__32603;
    wire N__32602;
    wire N__32601;
    wire N__32600;
    wire N__32599;
    wire N__32598;
    wire N__32597;
    wire N__32596;
    wire N__32595;
    wire N__32594;
    wire N__32593;
    wire N__32592;
    wire N__32591;
    wire N__32590;
    wire N__32589;
    wire N__32588;
    wire N__32579;
    wire N__32570;
    wire N__32569;
    wire N__32568;
    wire N__32567;
    wire N__32566;
    wire N__32565;
    wire N__32564;
    wire N__32563;
    wire N__32562;
    wire N__32561;
    wire N__32560;
    wire N__32559;
    wire N__32558;
    wire N__32557;
    wire N__32556;
    wire N__32547;
    wire N__32538;
    wire N__32535;
    wire N__32532;
    wire N__32527;
    wire N__32518;
    wire N__32509;
    wire N__32500;
    wire N__32495;
    wire N__32490;
    wire N__32477;
    wire N__32474;
    wire N__32471;
    wire N__32468;
    wire N__32465;
    wire N__32462;
    wire N__32459;
    wire N__32456;
    wire N__32453;
    wire N__32450;
    wire N__32447;
    wire N__32444;
    wire N__32441;
    wire N__32438;
    wire N__32435;
    wire N__32432;
    wire N__32429;
    wire N__32426;
    wire N__32423;
    wire N__32420;
    wire N__32419;
    wire N__32418;
    wire N__32415;
    wire N__32412;
    wire N__32409;
    wire N__32408;
    wire N__32403;
    wire N__32400;
    wire N__32399;
    wire N__32398;
    wire N__32395;
    wire N__32392;
    wire N__32389;
    wire N__32386;
    wire N__32383;
    wire N__32378;
    wire N__32369;
    wire N__32368;
    wire N__32363;
    wire N__32362;
    wire N__32361;
    wire N__32358;
    wire N__32353;
    wire N__32348;
    wire N__32345;
    wire N__32342;
    wire N__32339;
    wire N__32336;
    wire N__32335;
    wire N__32332;
    wire N__32329;
    wire N__32324;
    wire N__32321;
    wire N__32318;
    wire N__32315;
    wire N__32312;
    wire N__32311;
    wire N__32308;
    wire N__32307;
    wire N__32304;
    wire N__32301;
    wire N__32298;
    wire N__32295;
    wire N__32294;
    wire N__32289;
    wire N__32286;
    wire N__32283;
    wire N__32276;
    wire N__32275;
    wire N__32272;
    wire N__32269;
    wire N__32268;
    wire N__32267;
    wire N__32262;
    wire N__32259;
    wire N__32256;
    wire N__32253;
    wire N__32246;
    wire N__32245;
    wire N__32244;
    wire N__32241;
    wire N__32238;
    wire N__32235;
    wire N__32232;
    wire N__32225;
    wire N__32222;
    wire N__32219;
    wire N__32218;
    wire N__32217;
    wire N__32216;
    wire N__32213;
    wire N__32210;
    wire N__32207;
    wire N__32204;
    wire N__32195;
    wire N__32192;
    wire N__32189;
    wire N__32186;
    wire N__32183;
    wire N__32180;
    wire N__32177;
    wire N__32174;
    wire N__32171;
    wire N__32168;
    wire N__32167;
    wire N__32164;
    wire N__32161;
    wire N__32156;
    wire N__32153;
    wire N__32150;
    wire N__32149;
    wire N__32148;
    wire N__32145;
    wire N__32140;
    wire N__32139;
    wire N__32138;
    wire N__32133;
    wire N__32128;
    wire N__32123;
    wire N__32120;
    wire N__32117;
    wire N__32114;
    wire N__32113;
    wire N__32112;
    wire N__32111;
    wire N__32108;
    wire N__32105;
    wire N__32102;
    wire N__32099;
    wire N__32096;
    wire N__32091;
    wire N__32084;
    wire N__32081;
    wire N__32078;
    wire N__32075;
    wire N__32074;
    wire N__32071;
    wire N__32068;
    wire N__32067;
    wire N__32064;
    wire N__32059;
    wire N__32054;
    wire N__32051;
    wire N__32048;
    wire N__32045;
    wire N__32042;
    wire N__32039;
    wire N__32036;
    wire N__32033;
    wire N__32030;
    wire N__32027;
    wire N__32024;
    wire N__32023;
    wire N__32020;
    wire N__32017;
    wire N__32012;
    wire N__32009;
    wire N__32006;
    wire N__32003;
    wire N__32002;
    wire N__32001;
    wire N__31998;
    wire N__31993;
    wire N__31988;
    wire N__31985;
    wire N__31982;
    wire N__31979;
    wire N__31976;
    wire N__31973;
    wire N__31972;
    wire N__31971;
    wire N__31968;
    wire N__31963;
    wire N__31958;
    wire N__31955;
    wire N__31952;
    wire N__31951;
    wire N__31950;
    wire N__31947;
    wire N__31944;
    wire N__31941;
    wire N__31934;
    wire N__31933;
    wire N__31930;
    wire N__31927;
    wire N__31926;
    wire N__31923;
    wire N__31920;
    wire N__31917;
    wire N__31914;
    wire N__31911;
    wire N__31904;
    wire N__31901;
    wire N__31898;
    wire N__31895;
    wire N__31894;
    wire N__31891;
    wire N__31888;
    wire N__31887;
    wire N__31886;
    wire N__31881;
    wire N__31876;
    wire N__31871;
    wire N__31868;
    wire N__31865;
    wire N__31862;
    wire N__31861;
    wire N__31860;
    wire N__31857;
    wire N__31852;
    wire N__31847;
    wire N__31844;
    wire N__31841;
    wire N__31838;
    wire N__31837;
    wire N__31834;
    wire N__31833;
    wire N__31830;
    wire N__31827;
    wire N__31824;
    wire N__31817;
    wire N__31814;
    wire N__31813;
    wire N__31812;
    wire N__31809;
    wire N__31806;
    wire N__31803;
    wire N__31796;
    wire N__31793;
    wire N__31792;
    wire N__31791;
    wire N__31788;
    wire N__31787;
    wire N__31786;
    wire N__31783;
    wire N__31780;
    wire N__31777;
    wire N__31772;
    wire N__31771;
    wire N__31768;
    wire N__31765;
    wire N__31762;
    wire N__31759;
    wire N__31756;
    wire N__31753;
    wire N__31750;
    wire N__31747;
    wire N__31740;
    wire N__31733;
    wire N__31732;
    wire N__31729;
    wire N__31726;
    wire N__31721;
    wire N__31718;
    wire N__31715;
    wire N__31714;
    wire N__31711;
    wire N__31708;
    wire N__31703;
    wire N__31700;
    wire N__31697;
    wire N__31694;
    wire N__31693;
    wire N__31690;
    wire N__31687;
    wire N__31682;
    wire N__31681;
    wire N__31676;
    wire N__31675;
    wire N__31672;
    wire N__31669;
    wire N__31666;
    wire N__31663;
    wire N__31658;
    wire N__31655;
    wire N__31652;
    wire N__31649;
    wire N__31646;
    wire N__31643;
    wire N__31642;
    wire N__31639;
    wire N__31636;
    wire N__31631;
    wire N__31628;
    wire N__31625;
    wire N__31622;
    wire N__31619;
    wire N__31616;
    wire N__31613;
    wire N__31610;
    wire N__31607;
    wire N__31604;
    wire N__31603;
    wire N__31600;
    wire N__31597;
    wire N__31592;
    wire N__31591;
    wire N__31588;
    wire N__31585;
    wire N__31580;
    wire N__31577;
    wire N__31574;
    wire N__31573;
    wire N__31570;
    wire N__31567;
    wire N__31564;
    wire N__31561;
    wire N__31558;
    wire N__31555;
    wire N__31550;
    wire N__31547;
    wire N__31544;
    wire N__31541;
    wire N__31540;
    wire N__31539;
    wire N__31536;
    wire N__31531;
    wire N__31526;
    wire N__31523;
    wire N__31520;
    wire N__31519;
    wire N__31516;
    wire N__31513;
    wire N__31508;
    wire N__31505;
    wire N__31502;
    wire N__31499;
    wire N__31496;
    wire N__31495;
    wire N__31492;
    wire N__31489;
    wire N__31484;
    wire N__31481;
    wire N__31480;
    wire N__31477;
    wire N__31474;
    wire N__31469;
    wire N__31466;
    wire N__31463;
    wire N__31462;
    wire N__31459;
    wire N__31456;
    wire N__31453;
    wire N__31450;
    wire N__31445;
    wire N__31442;
    wire N__31439;
    wire N__31438;
    wire N__31435;
    wire N__31432;
    wire N__31427;
    wire N__31424;
    wire N__31423;
    wire N__31420;
    wire N__31417;
    wire N__31414;
    wire N__31409;
    wire N__31406;
    wire N__31403;
    wire N__31400;
    wire N__31397;
    wire N__31394;
    wire N__31391;
    wire N__31388;
    wire N__31385;
    wire N__31384;
    wire N__31383;
    wire N__31380;
    wire N__31377;
    wire N__31374;
    wire N__31371;
    wire N__31368;
    wire N__31361;
    wire N__31358;
    wire N__31357;
    wire N__31354;
    wire N__31353;
    wire N__31350;
    wire N__31347;
    wire N__31344;
    wire N__31337;
    wire N__31334;
    wire N__31333;
    wire N__31330;
    wire N__31329;
    wire N__31326;
    wire N__31323;
    wire N__31320;
    wire N__31313;
    wire N__31310;
    wire N__31309;
    wire N__31306;
    wire N__31305;
    wire N__31302;
    wire N__31299;
    wire N__31296;
    wire N__31289;
    wire N__31286;
    wire N__31285;
    wire N__31282;
    wire N__31281;
    wire N__31278;
    wire N__31275;
    wire N__31272;
    wire N__31265;
    wire N__31262;
    wire N__31259;
    wire N__31256;
    wire N__31253;
    wire N__31250;
    wire N__31247;
    wire N__31246;
    wire N__31245;
    wire N__31242;
    wire N__31239;
    wire N__31236;
    wire N__31235;
    wire N__31232;
    wire N__31227;
    wire N__31224;
    wire N__31221;
    wire N__31218;
    wire N__31211;
    wire N__31210;
    wire N__31209;
    wire N__31206;
    wire N__31203;
    wire N__31200;
    wire N__31197;
    wire N__31192;
    wire N__31187;
    wire N__31184;
    wire N__31183;
    wire N__31182;
    wire N__31179;
    wire N__31176;
    wire N__31173;
    wire N__31166;
    wire N__31163;
    wire N__31162;
    wire N__31161;
    wire N__31158;
    wire N__31155;
    wire N__31152;
    wire N__31145;
    wire N__31142;
    wire N__31139;
    wire N__31136;
    wire N__31133;
    wire N__31132;
    wire N__31129;
    wire N__31126;
    wire N__31123;
    wire N__31120;
    wire N__31119;
    wire N__31114;
    wire N__31111;
    wire N__31108;
    wire N__31105;
    wire N__31100;
    wire N__31097;
    wire N__31094;
    wire N__31091;
    wire N__31090;
    wire N__31087;
    wire N__31084;
    wire N__31079;
    wire N__31078;
    wire N__31075;
    wire N__31072;
    wire N__31067;
    wire N__31064;
    wire N__31061;
    wire N__31058;
    wire N__31057;
    wire N__31054;
    wire N__31051;
    wire N__31046;
    wire N__31045;
    wire N__31042;
    wire N__31039;
    wire N__31034;
    wire N__31031;
    wire N__31028;
    wire N__31025;
    wire N__31024;
    wire N__31021;
    wire N__31018;
    wire N__31013;
    wire N__31012;
    wire N__31009;
    wire N__31006;
    wire N__31001;
    wire N__30998;
    wire N__30995;
    wire N__30992;
    wire N__30989;
    wire N__30986;
    wire N__30983;
    wire N__30980;
    wire N__30979;
    wire N__30976;
    wire N__30973;
    wire N__30968;
    wire N__30965;
    wire N__30962;
    wire N__30961;
    wire N__30958;
    wire N__30955;
    wire N__30950;
    wire N__30947;
    wire N__30944;
    wire N__30941;
    wire N__30938;
    wire N__30937;
    wire N__30934;
    wire N__30931;
    wire N__30926;
    wire N__30923;
    wire N__30922;
    wire N__30919;
    wire N__30916;
    wire N__30913;
    wire N__30908;
    wire N__30907;
    wire N__30904;
    wire N__30901;
    wire N__30896;
    wire N__30893;
    wire N__30892;
    wire N__30889;
    wire N__30886;
    wire N__30885;
    wire N__30880;
    wire N__30877;
    wire N__30872;
    wire N__30869;
    wire N__30868;
    wire N__30865;
    wire N__30862;
    wire N__30859;
    wire N__30856;
    wire N__30853;
    wire N__30850;
    wire N__30849;
    wire N__30846;
    wire N__30843;
    wire N__30840;
    wire N__30833;
    wire N__30830;
    wire N__30829;
    wire N__30826;
    wire N__30823;
    wire N__30820;
    wire N__30815;
    wire N__30814;
    wire N__30811;
    wire N__30808;
    wire N__30803;
    wire N__30800;
    wire N__30797;
    wire N__30794;
    wire N__30791;
    wire N__30788;
    wire N__30785;
    wire N__30782;
    wire N__30781;
    wire N__30778;
    wire N__30775;
    wire N__30772;
    wire N__30769;
    wire N__30768;
    wire N__30767;
    wire N__30764;
    wire N__30761;
    wire N__30758;
    wire N__30755;
    wire N__30752;
    wire N__30747;
    wire N__30746;
    wire N__30741;
    wire N__30738;
    wire N__30735;
    wire N__30728;
    wire N__30725;
    wire N__30722;
    wire N__30719;
    wire N__30716;
    wire N__30713;
    wire N__30710;
    wire N__30707;
    wire N__30704;
    wire N__30701;
    wire N__30698;
    wire N__30697;
    wire N__30696;
    wire N__30693;
    wire N__30690;
    wire N__30687;
    wire N__30684;
    wire N__30681;
    wire N__30680;
    wire N__30679;
    wire N__30676;
    wire N__30671;
    wire N__30668;
    wire N__30665;
    wire N__30662;
    wire N__30653;
    wire N__30650;
    wire N__30647;
    wire N__30644;
    wire N__30641;
    wire N__30640;
    wire N__30639;
    wire N__30636;
    wire N__30633;
    wire N__30630;
    wire N__30627;
    wire N__30624;
    wire N__30617;
    wire N__30614;
    wire N__30611;
    wire N__30608;
    wire N__30605;
    wire N__30602;
    wire N__30599;
    wire N__30596;
    wire N__30593;
    wire N__30590;
    wire N__30587;
    wire N__30584;
    wire N__30581;
    wire N__30580;
    wire N__30575;
    wire N__30572;
    wire N__30569;
    wire N__30568;
    wire N__30565;
    wire N__30562;
    wire N__30559;
    wire N__30558;
    wire N__30557;
    wire N__30554;
    wire N__30551;
    wire N__30548;
    wire N__30545;
    wire N__30542;
    wire N__30539;
    wire N__30534;
    wire N__30527;
    wire N__30524;
    wire N__30521;
    wire N__30518;
    wire N__30515;
    wire N__30514;
    wire N__30511;
    wire N__30508;
    wire N__30503;
    wire N__30500;
    wire N__30499;
    wire N__30496;
    wire N__30495;
    wire N__30492;
    wire N__30489;
    wire N__30486;
    wire N__30483;
    wire N__30480;
    wire N__30477;
    wire N__30476;
    wire N__30475;
    wire N__30472;
    wire N__30469;
    wire N__30466;
    wire N__30463;
    wire N__30460;
    wire N__30449;
    wire N__30446;
    wire N__30443;
    wire N__30440;
    wire N__30437;
    wire N__30436;
    wire N__30433;
    wire N__30430;
    wire N__30429;
    wire N__30424;
    wire N__30421;
    wire N__30418;
    wire N__30413;
    wire N__30410;
    wire N__30409;
    wire N__30406;
    wire N__30403;
    wire N__30402;
    wire N__30397;
    wire N__30394;
    wire N__30391;
    wire N__30386;
    wire N__30383;
    wire N__30380;
    wire N__30379;
    wire N__30378;
    wire N__30375;
    wire N__30372;
    wire N__30369;
    wire N__30364;
    wire N__30359;
    wire N__30356;
    wire N__30355;
    wire N__30352;
    wire N__30349;
    wire N__30348;
    wire N__30343;
    wire N__30340;
    wire N__30337;
    wire N__30332;
    wire N__30329;
    wire N__30326;
    wire N__30325;
    wire N__30322;
    wire N__30319;
    wire N__30318;
    wire N__30313;
    wire N__30310;
    wire N__30307;
    wire N__30302;
    wire N__30299;
    wire N__30298;
    wire N__30295;
    wire N__30292;
    wire N__30291;
    wire N__30286;
    wire N__30283;
    wire N__30280;
    wire N__30275;
    wire N__30272;
    wire N__30271;
    wire N__30268;
    wire N__30265;
    wire N__30262;
    wire N__30257;
    wire N__30254;
    wire N__30251;
    wire N__30250;
    wire N__30247;
    wire N__30244;
    wire N__30241;
    wire N__30236;
    wire N__30235;
    wire N__30234;
    wire N__30233;
    wire N__30232;
    wire N__30231;
    wire N__30230;
    wire N__30229;
    wire N__30228;
    wire N__30227;
    wire N__30226;
    wire N__30225;
    wire N__30224;
    wire N__30223;
    wire N__30222;
    wire N__30221;
    wire N__30220;
    wire N__30219;
    wire N__30218;
    wire N__30217;
    wire N__30216;
    wire N__30215;
    wire N__30214;
    wire N__30213;
    wire N__30204;
    wire N__30195;
    wire N__30194;
    wire N__30193;
    wire N__30192;
    wire N__30191;
    wire N__30190;
    wire N__30189;
    wire N__30180;
    wire N__30171;
    wire N__30162;
    wire N__30153;
    wire N__30150;
    wire N__30147;
    wire N__30142;
    wire N__30133;
    wire N__30130;
    wire N__30119;
    wire N__30110;
    wire N__30107;
    wire N__30106;
    wire N__30103;
    wire N__30100;
    wire N__30099;
    wire N__30094;
    wire N__30091;
    wire N__30088;
    wire N__30083;
    wire N__30080;
    wire N__30079;
    wire N__30074;
    wire N__30073;
    wire N__30070;
    wire N__30067;
    wire N__30064;
    wire N__30059;
    wire N__30056;
    wire N__30053;
    wire N__30052;
    wire N__30049;
    wire N__30046;
    wire N__30045;
    wire N__30042;
    wire N__30039;
    wire N__30036;
    wire N__30031;
    wire N__30026;
    wire N__30023;
    wire N__30022;
    wire N__30019;
    wire N__30016;
    wire N__30013;
    wire N__30010;
    wire N__30009;
    wire N__30004;
    wire N__30001;
    wire N__29998;
    wire N__29993;
    wire N__29990;
    wire N__29987;
    wire N__29986;
    wire N__29983;
    wire N__29980;
    wire N__29979;
    wire N__29974;
    wire N__29971;
    wire N__29968;
    wire N__29963;
    wire N__29960;
    wire N__29959;
    wire N__29958;
    wire N__29953;
    wire N__29950;
    wire N__29947;
    wire N__29942;
    wire N__29939;
    wire N__29938;
    wire N__29937;
    wire N__29932;
    wire N__29929;
    wire N__29926;
    wire N__29921;
    wire N__29918;
    wire N__29917;
    wire N__29914;
    wire N__29913;
    wire N__29910;
    wire N__29907;
    wire N__29904;
    wire N__29899;
    wire N__29894;
    wire N__29891;
    wire N__29888;
    wire N__29885;
    wire N__29884;
    wire N__29881;
    wire N__29878;
    wire N__29877;
    wire N__29872;
    wire N__29869;
    wire N__29866;
    wire N__29861;
    wire N__29858;
    wire N__29857;
    wire N__29852;
    wire N__29851;
    wire N__29848;
    wire N__29845;
    wire N__29842;
    wire N__29837;
    wire N__29834;
    wire N__29831;
    wire N__29828;
    wire N__29827;
    wire N__29826;
    wire N__29823;
    wire N__29820;
    wire N__29817;
    wire N__29814;
    wire N__29811;
    wire N__29804;
    wire N__29801;
    wire N__29800;
    wire N__29797;
    wire N__29794;
    wire N__29793;
    wire N__29790;
    wire N__29787;
    wire N__29784;
    wire N__29781;
    wire N__29778;
    wire N__29771;
    wire N__29768;
    wire N__29767;
    wire N__29762;
    wire N__29761;
    wire N__29758;
    wire N__29755;
    wire N__29752;
    wire N__29747;
    wire N__29744;
    wire N__29743;
    wire N__29740;
    wire N__29737;
    wire N__29736;
    wire N__29731;
    wire N__29728;
    wire N__29725;
    wire N__29720;
    wire N__29717;
    wire N__29716;
    wire N__29713;
    wire N__29710;
    wire N__29709;
    wire N__29704;
    wire N__29701;
    wire N__29698;
    wire N__29693;
    wire N__29690;
    wire N__29687;
    wire N__29686;
    wire N__29683;
    wire N__29680;
    wire N__29679;
    wire N__29674;
    wire N__29671;
    wire N__29668;
    wire N__29663;
    wire N__29660;
    wire N__29657;
    wire N__29654;
    wire N__29653;
    wire N__29650;
    wire N__29647;
    wire N__29642;
    wire N__29639;
    wire N__29636;
    wire N__29635;
    wire N__29632;
    wire N__29631;
    wire N__29628;
    wire N__29625;
    wire N__29622;
    wire N__29615;
    wire N__29612;
    wire N__29609;
    wire N__29608;
    wire N__29605;
    wire N__29602;
    wire N__29601;
    wire N__29598;
    wire N__29595;
    wire N__29592;
    wire N__29589;
    wire N__29586;
    wire N__29579;
    wire N__29576;
    wire N__29575;
    wire N__29572;
    wire N__29569;
    wire N__29566;
    wire N__29565;
    wire N__29560;
    wire N__29557;
    wire N__29554;
    wire N__29549;
    wire N__29546;
    wire N__29545;
    wire N__29542;
    wire N__29539;
    wire N__29538;
    wire N__29533;
    wire N__29530;
    wire N__29527;
    wire N__29522;
    wire N__29519;
    wire N__29518;
    wire N__29515;
    wire N__29512;
    wire N__29507;
    wire N__29506;
    wire N__29503;
    wire N__29500;
    wire N__29497;
    wire N__29492;
    wire N__29489;
    wire N__29486;
    wire N__29483;
    wire N__29482;
    wire N__29479;
    wire N__29476;
    wire N__29471;
    wire N__29468;
    wire N__29465;
    wire N__29464;
    wire N__29461;
    wire N__29458;
    wire N__29453;
    wire N__29450;
    wire N__29447;
    wire N__29446;
    wire N__29443;
    wire N__29440;
    wire N__29437;
    wire N__29434;
    wire N__29429;
    wire N__29426;
    wire N__29423;
    wire N__29420;
    wire N__29417;
    wire N__29416;
    wire N__29413;
    wire N__29410;
    wire N__29405;
    wire N__29402;
    wire N__29399;
    wire N__29396;
    wire N__29393;
    wire N__29390;
    wire N__29389;
    wire N__29386;
    wire N__29383;
    wire N__29378;
    wire N__29375;
    wire N__29372;
    wire N__29369;
    wire N__29368;
    wire N__29365;
    wire N__29362;
    wire N__29359;
    wire N__29356;
    wire N__29351;
    wire N__29348;
    wire N__29345;
    wire N__29342;
    wire N__29339;
    wire N__29338;
    wire N__29335;
    wire N__29332;
    wire N__29327;
    wire N__29324;
    wire N__29321;
    wire N__29318;
    wire N__29315;
    wire N__29312;
    wire N__29309;
    wire N__29306;
    wire N__29303;
    wire N__29300;
    wire N__29297;
    wire N__29294;
    wire N__29291;
    wire N__29288;
    wire N__29285;
    wire N__29282;
    wire N__29279;
    wire N__29276;
    wire N__29273;
    wire N__29272;
    wire N__29271;
    wire N__29268;
    wire N__29265;
    wire N__29264;
    wire N__29263;
    wire N__29260;
    wire N__29257;
    wire N__29254;
    wire N__29247;
    wire N__29244;
    wire N__29239;
    wire N__29234;
    wire N__29231;
    wire N__29228;
    wire N__29225;
    wire N__29222;
    wire N__29219;
    wire N__29216;
    wire N__29213;
    wire N__29212;
    wire N__29209;
    wire N__29206;
    wire N__29201;
    wire N__29198;
    wire N__29195;
    wire N__29192;
    wire N__29189;
    wire N__29188;
    wire N__29185;
    wire N__29184;
    wire N__29177;
    wire N__29174;
    wire N__29171;
    wire N__29168;
    wire N__29165;
    wire N__29164;
    wire N__29161;
    wire N__29158;
    wire N__29153;
    wire N__29150;
    wire N__29147;
    wire N__29144;
    wire N__29141;
    wire N__29138;
    wire N__29135;
    wire N__29132;
    wire N__29129;
    wire N__29126;
    wire N__29123;
    wire N__29120;
    wire N__29117;
    wire N__29114;
    wire N__29111;
    wire N__29108;
    wire N__29107;
    wire N__29106;
    wire N__29103;
    wire N__29100;
    wire N__29097;
    wire N__29092;
    wire N__29087;
    wire N__29084;
    wire N__29081;
    wire N__29078;
    wire N__29075;
    wire N__29072;
    wire N__29069;
    wire N__29066;
    wire N__29063;
    wire N__29060;
    wire N__29057;
    wire N__29056;
    wire N__29053;
    wire N__29050;
    wire N__29045;
    wire N__29042;
    wire N__29039;
    wire N__29036;
    wire N__29035;
    wire N__29032;
    wire N__29029;
    wire N__29024;
    wire N__29021;
    wire N__29018;
    wire N__29015;
    wire N__29014;
    wire N__29013;
    wire N__29010;
    wire N__29007;
    wire N__29004;
    wire N__29001;
    wire N__28998;
    wire N__28991;
    wire N__28988;
    wire N__28985;
    wire N__28982;
    wire N__28979;
    wire N__28976;
    wire N__28975;
    wire N__28974;
    wire N__28971;
    wire N__28968;
    wire N__28965;
    wire N__28962;
    wire N__28959;
    wire N__28952;
    wire N__28949;
    wire N__28946;
    wire N__28943;
    wire N__28940;
    wire N__28937;
    wire N__28934;
    wire N__28933;
    wire N__28930;
    wire N__28929;
    wire N__28926;
    wire N__28923;
    wire N__28920;
    wire N__28913;
    wire N__28910;
    wire N__28907;
    wire N__28904;
    wire N__28901;
    wire N__28898;
    wire N__28897;
    wire N__28896;
    wire N__28893;
    wire N__28890;
    wire N__28887;
    wire N__28884;
    wire N__28881;
    wire N__28876;
    wire N__28871;
    wire N__28868;
    wire N__28865;
    wire N__28862;
    wire N__28859;
    wire N__28856;
    wire N__28853;
    wire N__28850;
    wire N__28847;
    wire N__28844;
    wire N__28841;
    wire N__28840;
    wire N__28839;
    wire N__28836;
    wire N__28833;
    wire N__28830;
    wire N__28827;
    wire N__28824;
    wire N__28817;
    wire N__28814;
    wire N__28811;
    wire N__28808;
    wire N__28805;
    wire N__28802;
    wire N__28801;
    wire N__28800;
    wire N__28797;
    wire N__28794;
    wire N__28791;
    wire N__28788;
    wire N__28785;
    wire N__28778;
    wire N__28775;
    wire N__28772;
    wire N__28769;
    wire N__28766;
    wire N__28763;
    wire N__28760;
    wire N__28757;
    wire N__28754;
    wire N__28751;
    wire N__28748;
    wire N__28745;
    wire N__28742;
    wire N__28739;
    wire N__28736;
    wire N__28733;
    wire N__28730;
    wire N__28727;
    wire N__28724;
    wire N__28721;
    wire N__28718;
    wire N__28715;
    wire N__28712;
    wire N__28709;
    wire N__28706;
    wire N__28703;
    wire N__28700;
    wire N__28697;
    wire N__28696;
    wire N__28695;
    wire N__28692;
    wire N__28689;
    wire N__28686;
    wire N__28679;
    wire N__28676;
    wire N__28673;
    wire N__28670;
    wire N__28667;
    wire N__28664;
    wire N__28663;
    wire N__28662;
    wire N__28659;
    wire N__28656;
    wire N__28653;
    wire N__28646;
    wire N__28643;
    wire N__28640;
    wire N__28637;
    wire N__28636;
    wire N__28635;
    wire N__28632;
    wire N__28629;
    wire N__28626;
    wire N__28623;
    wire N__28616;
    wire N__28613;
    wire N__28610;
    wire N__28607;
    wire N__28604;
    wire N__28601;
    wire N__28598;
    wire N__28595;
    wire N__28592;
    wire N__28589;
    wire N__28586;
    wire N__28583;
    wire N__28580;
    wire N__28577;
    wire N__28574;
    wire N__28573;
    wire N__28570;
    wire N__28567;
    wire N__28562;
    wire N__28559;
    wire N__28556;
    wire N__28553;
    wire N__28550;
    wire N__28547;
    wire N__28544;
    wire N__28541;
    wire N__28538;
    wire N__28535;
    wire N__28532;
    wire N__28529;
    wire N__28526;
    wire N__28523;
    wire N__28520;
    wire N__28517;
    wire N__28514;
    wire N__28511;
    wire N__28508;
    wire N__28505;
    wire N__28502;
    wire N__28499;
    wire N__28496;
    wire N__28493;
    wire N__28490;
    wire N__28487;
    wire N__28484;
    wire N__28483;
    wire N__28480;
    wire N__28479;
    wire N__28478;
    wire N__28475;
    wire N__28472;
    wire N__28469;
    wire N__28466;
    wire N__28465;
    wire N__28462;
    wire N__28459;
    wire N__28454;
    wire N__28451;
    wire N__28442;
    wire N__28439;
    wire N__28436;
    wire N__28433;
    wire N__28430;
    wire N__28427;
    wire N__28426;
    wire N__28423;
    wire N__28420;
    wire N__28419;
    wire N__28416;
    wire N__28415;
    wire N__28412;
    wire N__28409;
    wire N__28408;
    wire N__28405;
    wire N__28402;
    wire N__28399;
    wire N__28396;
    wire N__28393;
    wire N__28382;
    wire N__28379;
    wire N__28376;
    wire N__28373;
    wire N__28370;
    wire N__28367;
    wire N__28364;
    wire N__28361;
    wire N__28358;
    wire N__28355;
    wire N__28352;
    wire N__28349;
    wire N__28346;
    wire N__28343;
    wire N__28340;
    wire N__28337;
    wire N__28334;
    wire N__28331;
    wire N__28328;
    wire N__28325;
    wire N__28322;
    wire N__28319;
    wire N__28318;
    wire N__28317;
    wire N__28316;
    wire N__28315;
    wire N__28314;
    wire N__28313;
    wire N__28310;
    wire N__28309;
    wire N__28308;
    wire N__28307;
    wire N__28306;
    wire N__28305;
    wire N__28304;
    wire N__28303;
    wire N__28302;
    wire N__28301;
    wire N__28300;
    wire N__28299;
    wire N__28298;
    wire N__28297;
    wire N__28296;
    wire N__28293;
    wire N__28290;
    wire N__28281;
    wire N__28270;
    wire N__28269;
    wire N__28268;
    wire N__28267;
    wire N__28266;
    wire N__28265;
    wire N__28264;
    wire N__28263;
    wire N__28262;
    wire N__28261;
    wire N__28260;
    wire N__28257;
    wire N__28246;
    wire N__28237;
    wire N__28234;
    wire N__28233;
    wire N__28230;
    wire N__28225;
    wire N__28222;
    wire N__28211;
    wire N__28202;
    wire N__28199;
    wire N__28194;
    wire N__28191;
    wire N__28188;
    wire N__28183;
    wire N__28166;
    wire N__28165;
    wire N__28164;
    wire N__28163;
    wire N__28162;
    wire N__28161;
    wire N__28160;
    wire N__28159;
    wire N__28158;
    wire N__28157;
    wire N__28156;
    wire N__28153;
    wire N__28152;
    wire N__28151;
    wire N__28150;
    wire N__28149;
    wire N__28148;
    wire N__28147;
    wire N__28146;
    wire N__28145;
    wire N__28144;
    wire N__28143;
    wire N__28140;
    wire N__28139;
    wire N__28136;
    wire N__28133;
    wire N__28130;
    wire N__28129;
    wire N__28126;
    wire N__28123;
    wire N__28114;
    wire N__28111;
    wire N__28108;
    wire N__28105;
    wire N__28102;
    wire N__28101;
    wire N__28100;
    wire N__28099;
    wire N__28098;
    wire N__28095;
    wire N__28092;
    wire N__28089;
    wire N__28086;
    wire N__28077;
    wire N__28068;
    wire N__28061;
    wire N__28056;
    wire N__28053;
    wire N__28046;
    wire N__28035;
    wire N__28030;
    wire N__28027;
    wire N__28024;
    wire N__28019;
    wire N__28004;
    wire N__28003;
    wire N__28002;
    wire N__28001;
    wire N__28000;
    wire N__27999;
    wire N__27998;
    wire N__27997;
    wire N__27996;
    wire N__27985;
    wire N__27984;
    wire N__27983;
    wire N__27982;
    wire N__27981;
    wire N__27980;
    wire N__27979;
    wire N__27978;
    wire N__27977;
    wire N__27976;
    wire N__27975;
    wire N__27974;
    wire N__27971;
    wire N__27968;
    wire N__27967;
    wire N__27966;
    wire N__27965;
    wire N__27962;
    wire N__27961;
    wire N__27960;
    wire N__27957;
    wire N__27956;
    wire N__27955;
    wire N__27954;
    wire N__27953;
    wire N__27952;
    wire N__27951;
    wire N__27948;
    wire N__27939;
    wire N__27936;
    wire N__27935;
    wire N__27932;
    wire N__27929;
    wire N__27926;
    wire N__27921;
    wire N__27912;
    wire N__27907;
    wire N__27904;
    wire N__27901;
    wire N__27892;
    wire N__27883;
    wire N__27878;
    wire N__27875;
    wire N__27868;
    wire N__27865;
    wire N__27856;
    wire N__27847;
    wire N__27836;
    wire N__27833;
    wire N__27832;
    wire N__27831;
    wire N__27828;
    wire N__27825;
    wire N__27822;
    wire N__27821;
    wire N__27820;
    wire N__27819;
    wire N__27818;
    wire N__27817;
    wire N__27810;
    wire N__27805;
    wire N__27802;
    wire N__27799;
    wire N__27796;
    wire N__27793;
    wire N__27782;
    wire N__27781;
    wire N__27778;
    wire N__27775;
    wire N__27772;
    wire N__27769;
    wire N__27766;
    wire N__27761;
    wire N__27758;
    wire N__27755;
    wire N__27752;
    wire N__27751;
    wire N__27750;
    wire N__27749;
    wire N__27744;
    wire N__27743;
    wire N__27740;
    wire N__27739;
    wire N__27738;
    wire N__27735;
    wire N__27732;
    wire N__27725;
    wire N__27722;
    wire N__27719;
    wire N__27714;
    wire N__27707;
    wire N__27706;
    wire N__27705;
    wire N__27700;
    wire N__27699;
    wire N__27698;
    wire N__27697;
    wire N__27696;
    wire N__27693;
    wire N__27690;
    wire N__27681;
    wire N__27674;
    wire N__27671;
    wire N__27668;
    wire N__27667;
    wire N__27666;
    wire N__27663;
    wire N__27658;
    wire N__27653;
    wire N__27650;
    wire N__27647;
    wire N__27644;
    wire N__27641;
    wire N__27638;
    wire N__27635;
    wire N__27632;
    wire N__27629;
    wire N__27626;
    wire N__27623;
    wire N__27620;
    wire N__27617;
    wire N__27614;
    wire N__27611;
    wire N__27608;
    wire N__27605;
    wire N__27602;
    wire N__27599;
    wire N__27598;
    wire N__27597;
    wire N__27596;
    wire N__27595;
    wire N__27592;
    wire N__27589;
    wire N__27586;
    wire N__27583;
    wire N__27580;
    wire N__27577;
    wire N__27574;
    wire N__27571;
    wire N__27568;
    wire N__27565;
    wire N__27562;
    wire N__27555;
    wire N__27552;
    wire N__27545;
    wire N__27542;
    wire N__27539;
    wire N__27536;
    wire N__27533;
    wire N__27530;
    wire N__27529;
    wire N__27526;
    wire N__27525;
    wire N__27522;
    wire N__27519;
    wire N__27516;
    wire N__27509;
    wire N__27506;
    wire N__27505;
    wire N__27504;
    wire N__27503;
    wire N__27500;
    wire N__27497;
    wire N__27494;
    wire N__27491;
    wire N__27488;
    wire N__27485;
    wire N__27482;
    wire N__27473;
    wire N__27470;
    wire N__27469;
    wire N__27466;
    wire N__27463;
    wire N__27460;
    wire N__27457;
    wire N__27454;
    wire N__27449;
    wire N__27448;
    wire N__27447;
    wire N__27444;
    wire N__27439;
    wire N__27434;
    wire N__27431;
    wire N__27428;
    wire N__27427;
    wire N__27426;
    wire N__27423;
    wire N__27420;
    wire N__27417;
    wire N__27416;
    wire N__27413;
    wire N__27408;
    wire N__27405;
    wire N__27404;
    wire N__27403;
    wire N__27400;
    wire N__27395;
    wire N__27390;
    wire N__27383;
    wire N__27380;
    wire N__27377;
    wire N__27376;
    wire N__27373;
    wire N__27370;
    wire N__27365;
    wire N__27362;
    wire N__27359;
    wire N__27358;
    wire N__27357;
    wire N__27356;
    wire N__27355;
    wire N__27354;
    wire N__27351;
    wire N__27350;
    wire N__27349;
    wire N__27348;
    wire N__27347;
    wire N__27346;
    wire N__27345;
    wire N__27344;
    wire N__27343;
    wire N__27342;
    wire N__27341;
    wire N__27340;
    wire N__27339;
    wire N__27338;
    wire N__27337;
    wire N__27336;
    wire N__27333;
    wire N__27326;
    wire N__27315;
    wire N__27306;
    wire N__27305;
    wire N__27304;
    wire N__27301;
    wire N__27300;
    wire N__27299;
    wire N__27298;
    wire N__27297;
    wire N__27296;
    wire N__27295;
    wire N__27294;
    wire N__27293;
    wire N__27292;
    wire N__27277;
    wire N__27270;
    wire N__27267;
    wire N__27266;
    wire N__27263;
    wire N__27256;
    wire N__27255;
    wire N__27252;
    wire N__27251;
    wire N__27248;
    wire N__27235;
    wire N__27232;
    wire N__27227;
    wire N__27224;
    wire N__27219;
    wire N__27212;
    wire N__27197;
    wire N__27196;
    wire N__27193;
    wire N__27192;
    wire N__27189;
    wire N__27188;
    wire N__27185;
    wire N__27182;
    wire N__27179;
    wire N__27176;
    wire N__27171;
    wire N__27164;
    wire N__27163;
    wire N__27162;
    wire N__27161;
    wire N__27160;
    wire N__27151;
    wire N__27150;
    wire N__27149;
    wire N__27148;
    wire N__27147;
    wire N__27146;
    wire N__27143;
    wire N__27142;
    wire N__27139;
    wire N__27136;
    wire N__27133;
    wire N__27126;
    wire N__27123;
    wire N__27122;
    wire N__27121;
    wire N__27120;
    wire N__27119;
    wire N__27118;
    wire N__27117;
    wire N__27116;
    wire N__27115;
    wire N__27114;
    wire N__27113;
    wire N__27112;
    wire N__27111;
    wire N__27110;
    wire N__27107;
    wire N__27106;
    wire N__27105;
    wire N__27102;
    wire N__27093;
    wire N__27090;
    wire N__27085;
    wire N__27076;
    wire N__27063;
    wire N__27060;
    wire N__27055;
    wire N__27050;
    wire N__27035;
    wire N__27032;
    wire N__27029;
    wire N__27026;
    wire N__27023;
    wire N__27022;
    wire N__27021;
    wire N__27020;
    wire N__27017;
    wire N__27016;
    wire N__27015;
    wire N__27014;
    wire N__27013;
    wire N__27010;
    wire N__27009;
    wire N__27008;
    wire N__27007;
    wire N__27006;
    wire N__27003;
    wire N__27000;
    wire N__26997;
    wire N__26994;
    wire N__26991;
    wire N__26988;
    wire N__26985;
    wire N__26982;
    wire N__26973;
    wire N__26970;
    wire N__26967;
    wire N__26966;
    wire N__26965;
    wire N__26964;
    wire N__26963;
    wire N__26962;
    wire N__26961;
    wire N__26960;
    wire N__26959;
    wire N__26958;
    wire N__26957;
    wire N__26956;
    wire N__26955;
    wire N__26954;
    wire N__26953;
    wire N__26950;
    wire N__26947;
    wire N__26942;
    wire N__26939;
    wire N__26936;
    wire N__26929;
    wire N__26922;
    wire N__26913;
    wire N__26910;
    wire N__26905;
    wire N__26896;
    wire N__26893;
    wire N__26888;
    wire N__26885;
    wire N__26864;
    wire N__26861;
    wire N__26860;
    wire N__26857;
    wire N__26854;
    wire N__26853;
    wire N__26848;
    wire N__26847;
    wire N__26844;
    wire N__26841;
    wire N__26838;
    wire N__26831;
    wire N__26828;
    wire N__26827;
    wire N__26826;
    wire N__26823;
    wire N__26820;
    wire N__26819;
    wire N__26816;
    wire N__26813;
    wire N__26810;
    wire N__26807;
    wire N__26798;
    wire N__26797;
    wire N__26794;
    wire N__26791;
    wire N__26788;
    wire N__26787;
    wire N__26786;
    wire N__26783;
    wire N__26780;
    wire N__26777;
    wire N__26774;
    wire N__26771;
    wire N__26768;
    wire N__26765;
    wire N__26756;
    wire N__26753;
    wire N__26752;
    wire N__26751;
    wire N__26750;
    wire N__26749;
    wire N__26748;
    wire N__26745;
    wire N__26742;
    wire N__26739;
    wire N__26736;
    wire N__26735;
    wire N__26734;
    wire N__26731;
    wire N__26728;
    wire N__26719;
    wire N__26714;
    wire N__26705;
    wire N__26702;
    wire N__26699;
    wire N__26698;
    wire N__26695;
    wire N__26692;
    wire N__26691;
    wire N__26688;
    wire N__26685;
    wire N__26682;
    wire N__26675;
    wire N__26674;
    wire N__26673;
    wire N__26672;
    wire N__26671;
    wire N__26668;
    wire N__26663;
    wire N__26658;
    wire N__26651;
    wire N__26648;
    wire N__26647;
    wire N__26646;
    wire N__26643;
    wire N__26640;
    wire N__26639;
    wire N__26638;
    wire N__26635;
    wire N__26630;
    wire N__26625;
    wire N__26618;
    wire N__26617;
    wire N__26614;
    wire N__26613;
    wire N__26612;
    wire N__26609;
    wire N__26604;
    wire N__26601;
    wire N__26594;
    wire N__26591;
    wire N__26590;
    wire N__26587;
    wire N__26584;
    wire N__26579;
    wire N__26576;
    wire N__26575;
    wire N__26574;
    wire N__26571;
    wire N__26564;
    wire N__26561;
    wire N__26558;
    wire N__26555;
    wire N__26554;
    wire N__26551;
    wire N__26550;
    wire N__26547;
    wire N__26544;
    wire N__26541;
    wire N__26538;
    wire N__26537;
    wire N__26536;
    wire N__26533;
    wire N__26528;
    wire N__26523;
    wire N__26516;
    wire N__26513;
    wire N__26510;
    wire N__26507;
    wire N__26506;
    wire N__26503;
    wire N__26500;
    wire N__26497;
    wire N__26492;
    wire N__26491;
    wire N__26488;
    wire N__26485;
    wire N__26480;
    wire N__26477;
    wire N__26474;
    wire N__26471;
    wire N__26468;
    wire N__26465;
    wire N__26462;
    wire N__26459;
    wire N__26456;
    wire N__26453;
    wire N__26450;
    wire N__26449;
    wire N__26444;
    wire N__26441;
    wire N__26438;
    wire N__26437;
    wire N__26432;
    wire N__26429;
    wire N__26426;
    wire N__26423;
    wire N__26420;
    wire N__26417;
    wire N__26414;
    wire N__26411;
    wire N__26408;
    wire N__26405;
    wire N__26402;
    wire N__26401;
    wire N__26396;
    wire N__26393;
    wire N__26392;
    wire N__26389;
    wire N__26386;
    wire N__26381;
    wire N__26378;
    wire N__26377;
    wire N__26374;
    wire N__26371;
    wire N__26366;
    wire N__26365;
    wire N__26364;
    wire N__26363;
    wire N__26360;
    wire N__26359;
    wire N__26352;
    wire N__26349;
    wire N__26346;
    wire N__26343;
    wire N__26340;
    wire N__26337;
    wire N__26334;
    wire N__26327;
    wire N__26324;
    wire N__26321;
    wire N__26318;
    wire N__26315;
    wire N__26312;
    wire N__26309;
    wire N__26306;
    wire N__26303;
    wire N__26300;
    wire N__26299;
    wire N__26298;
    wire N__26295;
    wire N__26292;
    wire N__26289;
    wire N__26286;
    wire N__26283;
    wire N__26280;
    wire N__26279;
    wire N__26278;
    wire N__26275;
    wire N__26270;
    wire N__26265;
    wire N__26258;
    wire N__26255;
    wire N__26252;
    wire N__26249;
    wire N__26246;
    wire N__26243;
    wire N__26240;
    wire N__26237;
    wire N__26236;
    wire N__26233;
    wire N__26230;
    wire N__26227;
    wire N__26226;
    wire N__26225;
    wire N__26222;
    wire N__26219;
    wire N__26216;
    wire N__26215;
    wire N__26212;
    wire N__26207;
    wire N__26204;
    wire N__26201;
    wire N__26198;
    wire N__26189;
    wire N__26186;
    wire N__26183;
    wire N__26180;
    wire N__26177;
    wire N__26176;
    wire N__26175;
    wire N__26172;
    wire N__26169;
    wire N__26166;
    wire N__26165;
    wire N__26162;
    wire N__26159;
    wire N__26156;
    wire N__26153;
    wire N__26150;
    wire N__26145;
    wire N__26138;
    wire N__26135;
    wire N__26132;
    wire N__26129;
    wire N__26126;
    wire N__26125;
    wire N__26122;
    wire N__26121;
    wire N__26118;
    wire N__26115;
    wire N__26112;
    wire N__26109;
    wire N__26106;
    wire N__26103;
    wire N__26102;
    wire N__26101;
    wire N__26096;
    wire N__26093;
    wire N__26088;
    wire N__26081;
    wire N__26078;
    wire N__26075;
    wire N__26072;
    wire N__26071;
    wire N__26068;
    wire N__26065;
    wire N__26062;
    wire N__26061;
    wire N__26058;
    wire N__26055;
    wire N__26054;
    wire N__26053;
    wire N__26050;
    wire N__26045;
    wire N__26042;
    wire N__26039;
    wire N__26036;
    wire N__26027;
    wire N__26024;
    wire N__26021;
    wire N__26018;
    wire N__26015;
    wire N__26014;
    wire N__26013;
    wire N__26010;
    wire N__26007;
    wire N__26006;
    wire N__26005;
    wire N__26002;
    wire N__25999;
    wire N__25994;
    wire N__25991;
    wire N__25988;
    wire N__25985;
    wire N__25980;
    wire N__25973;
    wire N__25970;
    wire N__25967;
    wire N__25964;
    wire N__25961;
    wire N__25958;
    wire N__25955;
    wire N__25952;
    wire N__25949;
    wire N__25948;
    wire N__25945;
    wire N__25942;
    wire N__25937;
    wire N__25936;
    wire N__25935;
    wire N__25934;
    wire N__25931;
    wire N__25928;
    wire N__25923;
    wire N__25916;
    wire N__25913;
    wire N__25910;
    wire N__25907;
    wire N__25906;
    wire N__25903;
    wire N__25900;
    wire N__25897;
    wire N__25894;
    wire N__25891;
    wire N__25890;
    wire N__25889;
    wire N__25888;
    wire N__25883;
    wire N__25880;
    wire N__25877;
    wire N__25874;
    wire N__25865;
    wire N__25862;
    wire N__25859;
    wire N__25856;
    wire N__25855;
    wire N__25852;
    wire N__25849;
    wire N__25846;
    wire N__25843;
    wire N__25842;
    wire N__25841;
    wire N__25840;
    wire N__25835;
    wire N__25832;
    wire N__25829;
    wire N__25826;
    wire N__25817;
    wire N__25814;
    wire N__25811;
    wire N__25808;
    wire N__25805;
    wire N__25802;
    wire N__25799;
    wire N__25796;
    wire N__25795;
    wire N__25792;
    wire N__25789;
    wire N__25786;
    wire N__25785;
    wire N__25782;
    wire N__25779;
    wire N__25776;
    wire N__25775;
    wire N__25774;
    wire N__25769;
    wire N__25766;
    wire N__25761;
    wire N__25754;
    wire N__25751;
    wire N__25750;
    wire N__25747;
    wire N__25746;
    wire N__25743;
    wire N__25740;
    wire N__25737;
    wire N__25736;
    wire N__25735;
    wire N__25732;
    wire N__25727;
    wire N__25722;
    wire N__25715;
    wire N__25714;
    wire N__25713;
    wire N__25710;
    wire N__25707;
    wire N__25704;
    wire N__25701;
    wire N__25698;
    wire N__25697;
    wire N__25694;
    wire N__25691;
    wire N__25688;
    wire N__25687;
    wire N__25684;
    wire N__25681;
    wire N__25676;
    wire N__25673;
    wire N__25664;
    wire N__25661;
    wire N__25658;
    wire N__25655;
    wire N__25654;
    wire N__25651;
    wire N__25648;
    wire N__25645;
    wire N__25642;
    wire N__25639;
    wire N__25636;
    wire N__25633;
    wire N__25628;
    wire N__25625;
    wire N__25622;
    wire N__25619;
    wire N__25616;
    wire N__25615;
    wire N__25612;
    wire N__25609;
    wire N__25606;
    wire N__25603;
    wire N__25600;
    wire N__25597;
    wire N__25592;
    wire N__25589;
    wire N__25586;
    wire N__25583;
    wire N__25580;
    wire N__25577;
    wire N__25574;
    wire N__25571;
    wire N__25568;
    wire N__25565;
    wire N__25562;
    wire N__25559;
    wire N__25558;
    wire N__25555;
    wire N__25552;
    wire N__25549;
    wire N__25548;
    wire N__25547;
    wire N__25546;
    wire N__25541;
    wire N__25536;
    wire N__25533;
    wire N__25526;
    wire N__25523;
    wire N__25520;
    wire N__25517;
    wire N__25514;
    wire N__25511;
    wire N__25510;
    wire N__25509;
    wire N__25506;
    wire N__25505;
    wire N__25502;
    wire N__25497;
    wire N__25494;
    wire N__25491;
    wire N__25490;
    wire N__25489;
    wire N__25486;
    wire N__25481;
    wire N__25476;
    wire N__25469;
    wire N__25466;
    wire N__25463;
    wire N__25460;
    wire N__25457;
    wire N__25454;
    wire N__25451;
    wire N__25448;
    wire N__25445;
    wire N__25442;
    wire N__25439;
    wire N__25436;
    wire N__25433;
    wire N__25430;
    wire N__25427;
    wire N__25424;
    wire N__25421;
    wire N__25418;
    wire N__25415;
    wire N__25412;
    wire N__25409;
    wire N__25406;
    wire N__25403;
    wire N__25400;
    wire N__25397;
    wire N__25394;
    wire N__25391;
    wire N__25388;
    wire N__25385;
    wire N__25382;
    wire N__25381;
    wire N__25380;
    wire N__25379;
    wire N__25378;
    wire N__25375;
    wire N__25372;
    wire N__25367;
    wire N__25364;
    wire N__25361;
    wire N__25358;
    wire N__25355;
    wire N__25352;
    wire N__25349;
    wire N__25346;
    wire N__25341;
    wire N__25334;
    wire N__25331;
    wire N__25328;
    wire N__25325;
    wire N__25324;
    wire N__25321;
    wire N__25318;
    wire N__25313;
    wire N__25310;
    wire N__25307;
    wire N__25304;
    wire N__25301;
    wire N__25298;
    wire N__25297;
    wire N__25294;
    wire N__25291;
    wire N__25286;
    wire N__25283;
    wire N__25280;
    wire N__25277;
    wire N__25276;
    wire N__25273;
    wire N__25270;
    wire N__25265;
    wire N__25262;
    wire N__25259;
    wire N__25256;
    wire N__25253;
    wire N__25250;
    wire N__25247;
    wire N__25244;
    wire N__25243;
    wire N__25240;
    wire N__25237;
    wire N__25232;
    wire N__25229;
    wire N__25226;
    wire N__25223;
    wire N__25222;
    wire N__25219;
    wire N__25216;
    wire N__25211;
    wire N__25208;
    wire N__25205;
    wire N__25202;
    wire N__25199;
    wire N__25196;
    wire N__25193;
    wire N__25190;
    wire N__25187;
    wire N__25184;
    wire N__25181;
    wire N__25178;
    wire N__25175;
    wire N__25172;
    wire N__25169;
    wire N__25166;
    wire N__25163;
    wire N__25160;
    wire N__25159;
    wire N__25156;
    wire N__25153;
    wire N__25150;
    wire N__25145;
    wire N__25142;
    wire N__25139;
    wire N__25136;
    wire N__25133;
    wire N__25130;
    wire N__25127;
    wire N__25126;
    wire N__25123;
    wire N__25120;
    wire N__25115;
    wire N__25112;
    wire N__25109;
    wire N__25106;
    wire N__25103;
    wire N__25100;
    wire N__25099;
    wire N__25096;
    wire N__25093;
    wire N__25088;
    wire N__25085;
    wire N__25082;
    wire N__25079;
    wire N__25076;
    wire N__25073;
    wire N__25070;
    wire N__25067;
    wire N__25066;
    wire N__25063;
    wire N__25060;
    wire N__25055;
    wire N__25052;
    wire N__25049;
    wire N__25046;
    wire N__25043;
    wire N__25040;
    wire N__25037;
    wire N__25034;
    wire N__25033;
    wire N__25030;
    wire N__25027;
    wire N__25022;
    wire N__25019;
    wire N__25016;
    wire N__25013;
    wire N__25010;
    wire N__25007;
    wire N__25006;
    wire N__25003;
    wire N__25000;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24986;
    wire N__24983;
    wire N__24980;
    wire N__24977;
    wire N__24974;
    wire N__24973;
    wire N__24970;
    wire N__24967;
    wire N__24962;
    wire N__24959;
    wire N__24956;
    wire N__24953;
    wire N__24952;
    wire N__24951;
    wire N__24950;
    wire N__24949;
    wire N__24946;
    wire N__24945;
    wire N__24944;
    wire N__24943;
    wire N__24942;
    wire N__24941;
    wire N__24940;
    wire N__24939;
    wire N__24938;
    wire N__24935;
    wire N__24932;
    wire N__24929;
    wire N__24926;
    wire N__24925;
    wire N__24922;
    wire N__24919;
    wire N__24910;
    wire N__24897;
    wire N__24892;
    wire N__24889;
    wire N__24886;
    wire N__24875;
    wire N__24872;
    wire N__24871;
    wire N__24870;
    wire N__24869;
    wire N__24868;
    wire N__24867;
    wire N__24866;
    wire N__24865;
    wire N__24864;
    wire N__24863;
    wire N__24862;
    wire N__24861;
    wire N__24856;
    wire N__24853;
    wire N__24846;
    wire N__24839;
    wire N__24836;
    wire N__24831;
    wire N__24818;
    wire N__24815;
    wire N__24812;
    wire N__24809;
    wire N__24806;
    wire N__24805;
    wire N__24802;
    wire N__24801;
    wire N__24798;
    wire N__24795;
    wire N__24792;
    wire N__24789;
    wire N__24786;
    wire N__24779;
    wire N__24776;
    wire N__24773;
    wire N__24770;
    wire N__24767;
    wire N__24764;
    wire N__24763;
    wire N__24760;
    wire N__24757;
    wire N__24752;
    wire N__24749;
    wire N__24746;
    wire N__24743;
    wire N__24742;
    wire N__24739;
    wire N__24736;
    wire N__24731;
    wire N__24728;
    wire N__24725;
    wire N__24722;
    wire N__24719;
    wire N__24716;
    wire N__24713;
    wire N__24710;
    wire N__24707;
    wire N__24706;
    wire N__24703;
    wire N__24700;
    wire N__24697;
    wire N__24692;
    wire N__24689;
    wire N__24686;
    wire N__24683;
    wire N__24680;
    wire N__24677;
    wire N__24674;
    wire N__24671;
    wire N__24668;
    wire N__24665;
    wire N__24664;
    wire N__24661;
    wire N__24658;
    wire N__24653;
    wire N__24650;
    wire N__24647;
    wire N__24644;
    wire N__24643;
    wire N__24640;
    wire N__24637;
    wire N__24632;
    wire N__24629;
    wire N__24626;
    wire N__24623;
    wire N__24620;
    wire N__24617;
    wire N__24614;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24602;
    wire N__24601;
    wire N__24598;
    wire N__24595;
    wire N__24590;
    wire N__24587;
    wire N__24584;
    wire N__24581;
    wire N__24580;
    wire N__24577;
    wire N__24576;
    wire N__24573;
    wire N__24570;
    wire N__24567;
    wire N__24560;
    wire N__24557;
    wire N__24556;
    wire N__24555;
    wire N__24552;
    wire N__24547;
    wire N__24542;
    wire N__24539;
    wire N__24536;
    wire N__24535;
    wire N__24532;
    wire N__24529;
    wire N__24526;
    wire N__24521;
    wire N__24518;
    wire N__24517;
    wire N__24516;
    wire N__24515;
    wire N__24512;
    wire N__24509;
    wire N__24504;
    wire N__24497;
    wire N__24496;
    wire N__24493;
    wire N__24490;
    wire N__24485;
    wire N__24482;
    wire N__24479;
    wire N__24476;
    wire N__24473;
    wire N__24470;
    wire N__24469;
    wire N__24468;
    wire N__24467;
    wire N__24462;
    wire N__24461;
    wire N__24460;
    wire N__24459;
    wire N__24458;
    wire N__24457;
    wire N__24454;
    wire N__24451;
    wire N__24450;
    wire N__24449;
    wire N__24446;
    wire N__24441;
    wire N__24438;
    wire N__24431;
    wire N__24428;
    wire N__24423;
    wire N__24418;
    wire N__24407;
    wire N__24406;
    wire N__24403;
    wire N__24400;
    wire N__24397;
    wire N__24392;
    wire N__24389;
    wire N__24388;
    wire N__24385;
    wire N__24382;
    wire N__24377;
    wire N__24374;
    wire N__24371;
    wire N__24368;
    wire N__24365;
    wire N__24364;
    wire N__24363;
    wire N__24362;
    wire N__24361;
    wire N__24360;
    wire N__24357;
    wire N__24356;
    wire N__24355;
    wire N__24354;
    wire N__24353;
    wire N__24352;
    wire N__24343;
    wire N__24340;
    wire N__24337;
    wire N__24336;
    wire N__24333;
    wire N__24332;
    wire N__24331;
    wire N__24330;
    wire N__24329;
    wire N__24328;
    wire N__24327;
    wire N__24326;
    wire N__24325;
    wire N__24324;
    wire N__24323;
    wire N__24314;
    wire N__24309;
    wire N__24306;
    wire N__24303;
    wire N__24300;
    wire N__24293;
    wire N__24284;
    wire N__24277;
    wire N__24270;
    wire N__24263;
    wire N__24254;
    wire N__24251;
    wire N__24248;
    wire N__24245;
    wire N__24242;
    wire N__24239;
    wire N__24236;
    wire N__24233;
    wire N__24230;
    wire N__24227;
    wire N__24224;
    wire N__24221;
    wire N__24218;
    wire N__24215;
    wire N__24212;
    wire N__24209;
    wire N__24206;
    wire N__24203;
    wire N__24200;
    wire N__24197;
    wire N__24194;
    wire N__24191;
    wire N__24188;
    wire N__24185;
    wire N__24182;
    wire N__24179;
    wire N__24176;
    wire N__24173;
    wire N__24170;
    wire N__24167;
    wire N__24164;
    wire N__24161;
    wire N__24158;
    wire N__24155;
    wire N__24152;
    wire N__24149;
    wire N__24146;
    wire N__24143;
    wire N__24140;
    wire N__24137;
    wire N__24136;
    wire N__24135;
    wire N__24130;
    wire N__24127;
    wire N__24126;
    wire N__24123;
    wire N__24120;
    wire N__24117;
    wire N__24114;
    wire N__24107;
    wire N__24104;
    wire N__24101;
    wire N__24098;
    wire N__24097;
    wire N__24096;
    wire N__24093;
    wire N__24088;
    wire N__24085;
    wire N__24084;
    wire N__24081;
    wire N__24078;
    wire N__24075;
    wire N__24072;
    wire N__24065;
    wire N__24062;
    wire N__24059;
    wire N__24056;
    wire N__24053;
    wire N__24050;
    wire N__24047;
    wire N__24046;
    wire N__24045;
    wire N__24042;
    wire N__24041;
    wire N__24040;
    wire N__24035;
    wire N__24032;
    wire N__24029;
    wire N__24026;
    wire N__24023;
    wire N__24020;
    wire N__24017;
    wire N__24014;
    wire N__24011;
    wire N__24002;
    wire N__23999;
    wire N__23996;
    wire N__23993;
    wire N__23990;
    wire N__23987;
    wire N__23984;
    wire N__23981;
    wire N__23978;
    wire N__23975;
    wire N__23972;
    wire N__23969;
    wire N__23966;
    wire N__23963;
    wire N__23960;
    wire N__23957;
    wire N__23954;
    wire N__23951;
    wire N__23948;
    wire N__23945;
    wire N__23942;
    wire N__23939;
    wire N__23936;
    wire N__23933;
    wire N__23930;
    wire N__23927;
    wire N__23924;
    wire N__23921;
    wire N__23918;
    wire N__23915;
    wire N__23912;
    wire N__23909;
    wire N__23906;
    wire N__23903;
    wire N__23900;
    wire N__23897;
    wire N__23894;
    wire N__23891;
    wire N__23888;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23876;
    wire N__23873;
    wire N__23870;
    wire N__23867;
    wire N__23864;
    wire N__23861;
    wire N__23858;
    wire N__23855;
    wire N__23852;
    wire N__23849;
    wire N__23846;
    wire N__23843;
    wire N__23840;
    wire N__23837;
    wire N__23834;
    wire N__23831;
    wire N__23828;
    wire N__23825;
    wire N__23822;
    wire N__23819;
    wire N__23816;
    wire N__23813;
    wire N__23810;
    wire N__23807;
    wire N__23804;
    wire N__23801;
    wire N__23798;
    wire N__23795;
    wire N__23792;
    wire N__23789;
    wire N__23786;
    wire N__23783;
    wire N__23780;
    wire N__23777;
    wire N__23774;
    wire N__23771;
    wire N__23768;
    wire N__23765;
    wire N__23762;
    wire N__23759;
    wire N__23756;
    wire N__23753;
    wire N__23750;
    wire N__23747;
    wire N__23744;
    wire N__23741;
    wire N__23738;
    wire N__23735;
    wire N__23732;
    wire N__23729;
    wire N__23726;
    wire N__23723;
    wire N__23720;
    wire N__23717;
    wire N__23714;
    wire N__23711;
    wire N__23708;
    wire N__23705;
    wire N__23702;
    wire N__23699;
    wire N__23696;
    wire N__23693;
    wire N__23690;
    wire N__23687;
    wire N__23684;
    wire N__23681;
    wire N__23678;
    wire N__23675;
    wire N__23672;
    wire N__23669;
    wire N__23666;
    wire N__23663;
    wire N__23660;
    wire N__23657;
    wire N__23654;
    wire N__23651;
    wire N__23648;
    wire N__23645;
    wire N__23642;
    wire N__23639;
    wire N__23636;
    wire N__23633;
    wire N__23630;
    wire N__23627;
    wire N__23624;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23603;
    wire N__23600;
    wire N__23597;
    wire N__23594;
    wire N__23591;
    wire N__23588;
    wire N__23585;
    wire N__23582;
    wire N__23579;
    wire N__23576;
    wire N__23573;
    wire N__23572;
    wire N__23571;
    wire N__23568;
    wire N__23565;
    wire N__23562;
    wire N__23557;
    wire N__23554;
    wire N__23551;
    wire N__23548;
    wire N__23545;
    wire N__23540;
    wire N__23537;
    wire N__23534;
    wire N__23531;
    wire N__23528;
    wire N__23525;
    wire N__23522;
    wire N__23519;
    wire N__23516;
    wire N__23513;
    wire N__23510;
    wire N__23507;
    wire N__23504;
    wire N__23501;
    wire N__23498;
    wire N__23495;
    wire N__23492;
    wire N__23489;
    wire N__23486;
    wire N__23483;
    wire N__23480;
    wire N__23477;
    wire N__23474;
    wire N__23471;
    wire N__23468;
    wire N__23465;
    wire N__23462;
    wire N__23459;
    wire N__23456;
    wire N__23453;
    wire N__23450;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23435;
    wire N__23432;
    wire N__23429;
    wire N__23426;
    wire N__23423;
    wire N__23420;
    wire N__23417;
    wire N__23414;
    wire N__23411;
    wire N__23408;
    wire N__23405;
    wire N__23402;
    wire N__23399;
    wire N__23396;
    wire N__23393;
    wire N__23390;
    wire N__23387;
    wire N__23384;
    wire N__23381;
    wire N__23378;
    wire N__23375;
    wire N__23372;
    wire N__23369;
    wire N__23366;
    wire N__23363;
    wire N__23360;
    wire N__23359;
    wire N__23356;
    wire N__23353;
    wire N__23348;
    wire N__23347;
    wire N__23344;
    wire N__23343;
    wire N__23340;
    wire N__23337;
    wire N__23334;
    wire N__23331;
    wire N__23326;
    wire N__23321;
    wire N__23320;
    wire N__23317;
    wire N__23314;
    wire N__23309;
    wire N__23306;
    wire N__23303;
    wire N__23300;
    wire N__23299;
    wire N__23296;
    wire N__23293;
    wire N__23288;
    wire N__23287;
    wire N__23284;
    wire N__23281;
    wire N__23276;
    wire N__23273;
    wire N__23270;
    wire N__23267;
    wire N__23264;
    wire N__23263;
    wire N__23262;
    wire N__23259;
    wire N__23254;
    wire N__23249;
    wire N__23248;
    wire N__23247;
    wire N__23246;
    wire N__23243;
    wire N__23240;
    wire N__23235;
    wire N__23228;
    wire N__23227;
    wire N__23224;
    wire N__23221;
    wire N__23216;
    wire N__23213;
    wire N__23212;
    wire N__23209;
    wire N__23206;
    wire N__23201;
    wire N__23198;
    wire N__23197;
    wire N__23194;
    wire N__23191;
    wire N__23186;
    wire N__23183;
    wire N__23182;
    wire N__23179;
    wire N__23176;
    wire N__23171;
    wire N__23168;
    wire N__23167;
    wire N__23164;
    wire N__23161;
    wire N__23156;
    wire N__23153;
    wire N__23152;
    wire N__23149;
    wire N__23146;
    wire N__23141;
    wire N__23138;
    wire N__23137;
    wire N__23134;
    wire N__23131;
    wire N__23126;
    wire N__23123;
    wire N__23122;
    wire N__23119;
    wire N__23116;
    wire N__23111;
    wire N__23108;
    wire N__23107;
    wire N__23104;
    wire N__23101;
    wire N__23096;
    wire N__23093;
    wire N__23092;
    wire N__23089;
    wire N__23086;
    wire N__23081;
    wire N__23078;
    wire N__23075;
    wire N__23074;
    wire N__23071;
    wire N__23068;
    wire N__23063;
    wire N__23060;
    wire N__23059;
    wire N__23056;
    wire N__23053;
    wire N__23048;
    wire N__23045;
    wire N__23044;
    wire N__23041;
    wire N__23038;
    wire N__23033;
    wire N__23030;
    wire N__23029;
    wire N__23026;
    wire N__23023;
    wire N__23018;
    wire N__23015;
    wire N__23014;
    wire N__23011;
    wire N__23008;
    wire N__23003;
    wire N__23000;
    wire N__22999;
    wire N__22996;
    wire N__22993;
    wire N__22988;
    wire N__22985;
    wire N__22982;
    wire N__22981;
    wire N__22978;
    wire N__22975;
    wire N__22970;
    wire N__22967;
    wire N__22964;
    wire N__22961;
    wire N__22958;
    wire N__22955;
    wire N__22954;
    wire N__22953;
    wire N__22952;
    wire N__22951;
    wire N__22950;
    wire N__22949;
    wire N__22946;
    wire N__22945;
    wire N__22942;
    wire N__22941;
    wire N__22938;
    wire N__22937;
    wire N__22936;
    wire N__22935;
    wire N__22934;
    wire N__22933;
    wire N__22930;
    wire N__22929;
    wire N__22926;
    wire N__22925;
    wire N__22908;
    wire N__22905;
    wire N__22904;
    wire N__22901;
    wire N__22900;
    wire N__22897;
    wire N__22896;
    wire N__22893;
    wire N__22892;
    wire N__22883;
    wire N__22880;
    wire N__22863;
    wire N__22860;
    wire N__22855;
    wire N__22852;
    wire N__22847;
    wire N__22846;
    wire N__22843;
    wire N__22840;
    wire N__22835;
    wire N__22832;
    wire N__22831;
    wire N__22828;
    wire N__22825;
    wire N__22822;
    wire N__22817;
    wire N__22814;
    wire N__22811;
    wire N__22808;
    wire N__22805;
    wire N__22804;
    wire N__22799;
    wire N__22796;
    wire N__22793;
    wire N__22792;
    wire N__22791;
    wire N__22786;
    wire N__22783;
    wire N__22778;
    wire N__22775;
    wire N__22772;
    wire N__22769;
    wire N__22766;
    wire N__22763;
    wire N__22762;
    wire N__22761;
    wire N__22758;
    wire N__22753;
    wire N__22752;
    wire N__22751;
    wire N__22748;
    wire N__22745;
    wire N__22740;
    wire N__22733;
    wire N__22730;
    wire N__22727;
    wire N__22724;
    wire N__22721;
    wire N__22718;
    wire N__22715;
    wire N__22712;
    wire N__22709;
    wire N__22706;
    wire N__22703;
    wire N__22700;
    wire N__22697;
    wire N__22694;
    wire N__22691;
    wire N__22688;
    wire N__22685;
    wire N__22682;
    wire N__22679;
    wire N__22676;
    wire N__22673;
    wire N__22670;
    wire N__22667;
    wire N__22664;
    wire N__22661;
    wire N__22658;
    wire N__22655;
    wire N__22652;
    wire N__22649;
    wire N__22646;
    wire N__22643;
    wire N__22640;
    wire N__22637;
    wire N__22634;
    wire N__22631;
    wire N__22628;
    wire N__22625;
    wire N__22622;
    wire N__22619;
    wire N__22616;
    wire N__22613;
    wire N__22610;
    wire N__22607;
    wire N__22604;
    wire N__22601;
    wire N__22598;
    wire N__22595;
    wire N__22592;
    wire N__22589;
    wire N__22586;
    wire N__22583;
    wire N__22580;
    wire N__22577;
    wire N__22574;
    wire N__22571;
    wire N__22568;
    wire N__22565;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22553;
    wire N__22550;
    wire N__22547;
    wire N__22544;
    wire N__22541;
    wire N__22538;
    wire N__22535;
    wire N__22532;
    wire N__22529;
    wire N__22526;
    wire N__22523;
    wire N__22520;
    wire N__22517;
    wire N__22514;
    wire N__22511;
    wire N__22508;
    wire N__22505;
    wire N__22502;
    wire N__22499;
    wire N__22496;
    wire N__22493;
    wire N__22490;
    wire N__22487;
    wire N__22484;
    wire N__22481;
    wire N__22478;
    wire N__22475;
    wire N__22472;
    wire N__22469;
    wire N__22466;
    wire N__22463;
    wire N__22460;
    wire N__22457;
    wire N__22454;
    wire N__22451;
    wire N__22448;
    wire N__22445;
    wire N__22442;
    wire N__22439;
    wire N__22436;
    wire N__22433;
    wire N__22430;
    wire N__22427;
    wire N__22424;
    wire N__22421;
    wire N__22418;
    wire N__22415;
    wire N__22412;
    wire N__22409;
    wire N__22406;
    wire N__22403;
    wire N__22400;
    wire N__22397;
    wire N__22394;
    wire N__22391;
    wire N__22388;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22376;
    wire N__22373;
    wire N__22370;
    wire N__22367;
    wire N__22364;
    wire N__22361;
    wire N__22360;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22346;
    wire N__22345;
    wire N__22340;
    wire N__22337;
    wire N__22334;
    wire N__22331;
    wire N__22330;
    wire N__22327;
    wire N__22324;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22312;
    wire N__22307;
    wire N__22304;
    wire N__22301;
    wire N__22298;
    wire N__22295;
    wire N__22294;
    wire N__22291;
    wire N__22288;
    wire N__22283;
    wire N__22280;
    wire N__22277;
    wire N__22276;
    wire N__22273;
    wire N__22270;
    wire N__22267;
    wire N__22264;
    wire N__22259;
    wire N__22256;
    wire N__22253;
    wire N__22252;
    wire N__22249;
    wire N__22248;
    wire N__22245;
    wire N__22244;
    wire N__22243;
    wire N__22242;
    wire N__22241;
    wire N__22240;
    wire N__22239;
    wire N__22236;
    wire N__22227;
    wire N__22224;
    wire N__22221;
    wire N__22216;
    wire N__22215;
    wire N__22204;
    wire N__22201;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22175;
    wire N__22174;
    wire N__22171;
    wire N__22168;
    wire N__22163;
    wire N__22160;
    wire N__22157;
    wire N__22156;
    wire N__22153;
    wire N__22150;
    wire N__22145;
    wire N__22142;
    wire N__22139;
    wire N__22138;
    wire N__22135;
    wire N__22132;
    wire N__22127;
    wire N__22124;
    wire N__22123;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22111;
    wire N__22108;
    wire N__22103;
    wire N__22100;
    wire N__22097;
    wire N__22096;
    wire N__22093;
    wire N__22088;
    wire N__22085;
    wire N__22082;
    wire N__22079;
    wire N__22078;
    wire N__22073;
    wire N__22070;
    wire N__22067;
    wire N__22066;
    wire N__22063;
    wire N__22060;
    wire N__22055;
    wire N__22052;
    wire N__22049;
    wire N__22046;
    wire N__22045;
    wire N__22042;
    wire N__22039;
    wire N__22034;
    wire N__22031;
    wire N__22030;
    wire N__22029;
    wire N__22026;
    wire N__22023;
    wire N__22020;
    wire N__22017;
    wire N__22012;
    wire N__22009;
    wire N__22004;
    wire N__22001;
    wire N__21998;
    wire N__21997;
    wire N__21996;
    wire N__21993;
    wire N__21990;
    wire N__21987;
    wire N__21984;
    wire N__21979;
    wire N__21974;
    wire N__21971;
    wire N__21970;
    wire N__21965;
    wire N__21962;
    wire N__21959;
    wire N__21956;
    wire N__21955;
    wire N__21952;
    wire N__21949;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21934;
    wire N__21931;
    wire N__21928;
    wire N__21923;
    wire N__21920;
    wire N__21919;
    wire N__21916;
    wire N__21913;
    wire N__21908;
    wire N__21905;
    wire N__21904;
    wire N__21901;
    wire N__21898;
    wire N__21893;
    wire N__21890;
    wire N__21889;
    wire N__21886;
    wire N__21883;
    wire N__21878;
    wire N__21875;
    wire N__21872;
    wire N__21869;
    wire N__21866;
    wire N__21863;
    wire N__21860;
    wire N__21857;
    wire N__21854;
    wire N__21851;
    wire N__21848;
    wire N__21845;
    wire N__21842;
    wire N__21839;
    wire N__21836;
    wire N__21833;
    wire N__21832;
    wire N__21831;
    wire N__21828;
    wire N__21825;
    wire N__21822;
    wire N__21817;
    wire N__21812;
    wire N__21809;
    wire N__21806;
    wire N__21805;
    wire N__21802;
    wire N__21801;
    wire N__21798;
    wire N__21797;
    wire N__21794;
    wire N__21791;
    wire N__21788;
    wire N__21785;
    wire N__21780;
    wire N__21777;
    wire N__21774;
    wire N__21771;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21757;
    wire N__21756;
    wire N__21753;
    wire N__21750;
    wire N__21747;
    wire N__21740;
    wire N__21737;
    wire N__21734;
    wire N__21731;
    wire N__21730;
    wire N__21729;
    wire N__21726;
    wire N__21723;
    wire N__21720;
    wire N__21715;
    wire N__21712;
    wire N__21709;
    wire N__21706;
    wire N__21701;
    wire N__21698;
    wire N__21697;
    wire N__21696;
    wire N__21693;
    wire N__21690;
    wire N__21687;
    wire N__21684;
    wire N__21679;
    wire N__21676;
    wire N__21673;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21653;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21641;
    wire N__21638;
    wire N__21635;
    wire N__21632;
    wire N__21629;
    wire N__21626;
    wire N__21623;
    wire N__21620;
    wire N__21617;
    wire N__21614;
    wire N__21611;
    wire N__21608;
    wire N__21605;
    wire N__21602;
    wire N__21599;
    wire N__21596;
    wire N__21593;
    wire N__21590;
    wire N__21589;
    wire N__21588;
    wire N__21587;
    wire N__21586;
    wire N__21585;
    wire N__21584;
    wire N__21583;
    wire N__21582;
    wire N__21577;
    wire N__21572;
    wire N__21561;
    wire N__21558;
    wire N__21555;
    wire N__21554;
    wire N__21551;
    wire N__21546;
    wire N__21543;
    wire N__21540;
    wire N__21537;
    wire N__21530;
    wire N__21529;
    wire N__21528;
    wire N__21527;
    wire N__21522;
    wire N__21517;
    wire N__21516;
    wire N__21515;
    wire N__21514;
    wire N__21513;
    wire N__21512;
    wire N__21509;
    wire N__21506;
    wire N__21495;
    wire N__21490;
    wire N__21487;
    wire N__21486;
    wire N__21483;
    wire N__21480;
    wire N__21477;
    wire N__21470;
    wire N__21469;
    wire N__21468;
    wire N__21465;
    wire N__21464;
    wire N__21461;
    wire N__21458;
    wire N__21453;
    wire N__21448;
    wire N__21445;
    wire N__21442;
    wire N__21441;
    wire N__21440;
    wire N__21439;
    wire N__21438;
    wire N__21437;
    wire N__21436;
    wire N__21435;
    wire N__21434;
    wire N__21431;
    wire N__21428;
    wire N__21423;
    wire N__21420;
    wire N__21417;
    wire N__21414;
    wire N__21411;
    wire N__21408;
    wire N__21405;
    wire N__21398;
    wire N__21397;
    wire N__21396;
    wire N__21395;
    wire N__21392;
    wire N__21385;
    wire N__21380;
    wire N__21379;
    wire N__21376;
    wire N__21369;
    wire N__21362;
    wire N__21359;
    wire N__21358;
    wire N__21357;
    wire N__21356;
    wire N__21355;
    wire N__21354;
    wire N__21353;
    wire N__21352;
    wire N__21351;
    wire N__21350;
    wire N__21349;
    wire N__21348;
    wire N__21347;
    wire N__21346;
    wire N__21345;
    wire N__21344;
    wire N__21343;
    wire N__21338;
    wire N__21335;
    wire N__21332;
    wire N__21329;
    wire N__21312;
    wire N__21297;
    wire N__21294;
    wire N__21281;
    wire N__21278;
    wire N__21275;
    wire N__21272;
    wire N__21269;
    wire N__21266;
    wire N__21263;
    wire N__21260;
    wire N__21257;
    wire N__21254;
    wire N__21253;
    wire N__21250;
    wire N__21247;
    wire N__21246;
    wire N__21241;
    wire N__21238;
    wire N__21235;
    wire N__21230;
    wire N__21227;
    wire N__21224;
    wire N__21221;
    wire N__21220;
    wire N__21217;
    wire N__21214;
    wire N__21209;
    wire N__21208;
    wire N__21205;
    wire N__21204;
    wire N__21203;
    wire N__21202;
    wire N__21201;
    wire N__21198;
    wire N__21197;
    wire N__21194;
    wire N__21191;
    wire N__21186;
    wire N__21183;
    wire N__21180;
    wire N__21177;
    wire N__21176;
    wire N__21173;
    wire N__21170;
    wire N__21169;
    wire N__21168;
    wire N__21167;
    wire N__21164;
    wire N__21157;
    wire N__21154;
    wire N__21151;
    wire N__21148;
    wire N__21145;
    wire N__21142;
    wire N__21139;
    wire N__21132;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21112;
    wire N__21111;
    wire N__21108;
    wire N__21105;
    wire N__21102;
    wire N__21095;
    wire N__21092;
    wire N__21091;
    wire N__21090;
    wire N__21087;
    wire N__21084;
    wire N__21081;
    wire N__21074;
    wire N__21071;
    wire N__21070;
    wire N__21069;
    wire N__21066;
    wire N__21063;
    wire N__21060;
    wire N__21053;
    wire N__21050;
    wire N__21049;
    wire N__21048;
    wire N__21045;
    wire N__21042;
    wire N__21039;
    wire N__21032;
    wire N__21029;
    wire N__21028;
    wire N__21027;
    wire N__21024;
    wire N__21021;
    wire N__21018;
    wire N__21011;
    wire N__21008;
    wire N__21007;
    wire N__21006;
    wire N__21003;
    wire N__21000;
    wire N__20997;
    wire N__20994;
    wire N__20987;
    wire N__20984;
    wire N__20983;
    wire N__20982;
    wire N__20981;
    wire N__20980;
    wire N__20979;
    wire N__20970;
    wire N__20969;
    wire N__20968;
    wire N__20967;
    wire N__20966;
    wire N__20961;
    wire N__20958;
    wire N__20949;
    wire N__20946;
    wire N__20939;
    wire N__20936;
    wire N__20935;
    wire N__20934;
    wire N__20931;
    wire N__20928;
    wire N__20925;
    wire N__20922;
    wire N__20915;
    wire N__20912;
    wire N__20909;
    wire N__20906;
    wire N__20903;
    wire N__20900;
    wire N__20897;
    wire N__20894;
    wire N__20891;
    wire N__20888;
    wire N__20885;
    wire N__20882;
    wire N__20879;
    wire N__20878;
    wire N__20877;
    wire N__20874;
    wire N__20871;
    wire N__20868;
    wire N__20861;
    wire N__20858;
    wire N__20857;
    wire N__20856;
    wire N__20853;
    wire N__20850;
    wire N__20847;
    wire N__20840;
    wire N__20837;
    wire N__20836;
    wire N__20835;
    wire N__20832;
    wire N__20829;
    wire N__20826;
    wire N__20819;
    wire N__20816;
    wire N__20813;
    wire N__20810;
    wire N__20807;
    wire N__20804;
    wire N__20801;
    wire N__20798;
    wire N__20795;
    wire N__20792;
    wire N__20789;
    wire N__20786;
    wire N__20783;
    wire N__20780;
    wire N__20777;
    wire N__20774;
    wire N__20771;
    wire N__20768;
    wire N__20765;
    wire N__20762;
    wire N__20759;
    wire N__20756;
    wire N__20753;
    wire N__20750;
    wire N__20747;
    wire N__20744;
    wire N__20741;
    wire N__20738;
    wire N__20735;
    wire N__20732;
    wire N__20729;
    wire N__20726;
    wire N__20723;
    wire N__20720;
    wire N__20717;
    wire N__20714;
    wire N__20711;
    wire N__20708;
    wire N__20705;
    wire N__20702;
    wire N__20699;
    wire N__20696;
    wire N__20693;
    wire N__20690;
    wire N__20687;
    wire N__20684;
    wire N__20681;
    wire N__20678;
    wire N__20675;
    wire N__20674;
    wire N__20671;
    wire N__20668;
    wire N__20663;
    wire N__20662;
    wire N__20659;
    wire N__20658;
    wire N__20655;
    wire N__20652;
    wire N__20649;
    wire N__20644;
    wire N__20639;
    wire N__20636;
    wire N__20633;
    wire N__20630;
    wire N__20627;
    wire N__20624;
    wire N__20621;
    wire N__20618;
    wire N__20615;
    wire N__20612;
    wire N__20609;
    wire N__20606;
    wire N__20603;
    wire N__20600;
    wire N__20597;
    wire N__20594;
    wire N__20591;
    wire N__20588;
    wire N__20585;
    wire N__20582;
    wire N__20579;
    wire N__20576;
    wire N__20573;
    wire N__20570;
    wire N__20567;
    wire N__20564;
    wire N__20561;
    wire N__20558;
    wire N__20555;
    wire N__20552;
    wire N__20549;
    wire N__20546;
    wire N__20543;
    wire N__20540;
    wire N__20537;
    wire N__20534;
    wire N__20531;
    wire N__20528;
    wire N__20525;
    wire N__20522;
    wire N__20519;
    wire N__20516;
    wire N__20513;
    wire N__20510;
    wire N__20507;
    wire N__20504;
    wire N__20501;
    wire N__20498;
    wire N__20495;
    wire N__20492;
    wire N__20489;
    wire N__20486;
    wire N__20483;
    wire N__20480;
    wire N__20477;
    wire N__20476;
    wire N__20473;
    wire N__20470;
    wire N__20467;
    wire N__20464;
    wire N__20461;
    wire N__20458;
    wire N__20453;
    wire N__20450;
    wire N__20449;
    wire N__20446;
    wire N__20445;
    wire N__20442;
    wire N__20439;
    wire N__20436;
    wire N__20429;
    wire N__20426;
    wire N__20423;
    wire N__20420;
    wire N__20417;
    wire N__20414;
    wire N__20411;
    wire N__20408;
    wire N__20405;
    wire N__20402;
    wire N__20399;
    wire N__20396;
    wire N__20393;
    wire N__20390;
    wire N__20387;
    wire N__20384;
    wire N__20381;
    wire N__20378;
    wire N__20375;
    wire N__20372;
    wire N__20369;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20330;
    wire N__20327;
    wire N__20324;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20312;
    wire N__20309;
    wire N__20306;
    wire N__20303;
    wire N__20300;
    wire N__20297;
    wire N__20294;
    wire N__20291;
    wire N__20290;
    wire N__20287;
    wire N__20286;
    wire N__20283;
    wire N__20280;
    wire N__20277;
    wire N__20270;
    wire N__20267;
    wire N__20264;
    wire N__20261;
    wire N__20260;
    wire N__20259;
    wire N__20258;
    wire N__20257;
    wire N__20254;
    wire N__20253;
    wire N__20250;
    wire N__20239;
    wire N__20236;
    wire N__20235;
    wire N__20234;
    wire N__20233;
    wire N__20228;
    wire N__20225;
    wire N__20220;
    wire N__20213;
    wire N__20210;
    wire N__20207;
    wire N__20206;
    wire N__20205;
    wire N__20204;
    wire N__20201;
    wire N__20198;
    wire N__20195;
    wire N__20192;
    wire N__20191;
    wire N__20190;
    wire N__20179;
    wire N__20176;
    wire N__20173;
    wire N__20172;
    wire N__20169;
    wire N__20166;
    wire N__20163;
    wire N__20156;
    wire N__20153;
    wire N__20150;
    wire N__20147;
    wire N__20144;
    wire N__20141;
    wire N__20138;
    wire N__20135;
    wire N__20132;
    wire N__20129;
    wire N__20126;
    wire N__20123;
    wire N__20120;
    wire N__20119;
    wire N__20116;
    wire N__20113;
    wire N__20110;
    wire N__20105;
    wire N__20102;
    wire N__20099;
    wire N__20096;
    wire N__20093;
    wire N__20092;
    wire N__20089;
    wire N__20086;
    wire N__20081;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20071;
    wire N__20068;
    wire N__20065;
    wire N__20060;
    wire N__20057;
    wire N__20054;
    wire N__20051;
    wire N__20048;
    wire N__20045;
    wire N__20042;
    wire N__20039;
    wire N__20036;
    wire N__20033;
    wire N__20030;
    wire N__20027;
    wire N__20026;
    wire N__20025;
    wire N__20022;
    wire N__20019;
    wire N__20016;
    wire N__20013;
    wire N__20010;
    wire N__20007;
    wire N__20000;
    wire N__19999;
    wire N__19998;
    wire N__19995;
    wire N__19992;
    wire N__19989;
    wire N__19986;
    wire N__19983;
    wire N__19980;
    wire N__19977;
    wire N__19974;
    wire N__19971;
    wire N__19964;
    wire N__19963;
    wire N__19960;
    wire N__19957;
    wire N__19956;
    wire N__19953;
    wire N__19950;
    wire N__19947;
    wire N__19942;
    wire N__19939;
    wire N__19936;
    wire N__19933;
    wire N__19928;
    wire N__19925;
    wire N__19922;
    wire N__19921;
    wire N__19918;
    wire N__19917;
    wire N__19914;
    wire N__19911;
    wire N__19908;
    wire N__19905;
    wire N__19900;
    wire N__19895;
    wire N__19892;
    wire N__19889;
    wire N__19886;
    wire N__19883;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19868;
    wire N__19865;
    wire N__19862;
    wire N__19859;
    wire N__19856;
    wire N__19853;
    wire N__19850;
    wire N__19847;
    wire N__19844;
    wire N__19841;
    wire N__19838;
    wire N__19835;
    wire N__19832;
    wire N__19829;
    wire N__19826;
    wire N__19823;
    wire N__19822;
    wire N__19819;
    wire N__19816;
    wire N__19813;
    wire N__19810;
    wire N__19805;
    wire N__19802;
    wire N__19801;
    wire N__19800;
    wire N__19797;
    wire N__19794;
    wire N__19791;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19769;
    wire N__19768;
    wire N__19765;
    wire N__19762;
    wire N__19759;
    wire N__19754;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19738;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19712;
    wire N__19709;
    wire N__19706;
    wire N__19703;
    wire N__19700;
    wire N__19697;
    wire N__19694;
    wire N__19691;
    wire N__19688;
    wire N__19685;
    wire N__19682;
    wire N__19679;
    wire N__19676;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19598;
    wire N__19595;
    wire N__19592;
    wire N__19589;
    wire N__19586;
    wire N__19583;
    wire N__19580;
    wire N__19577;
    wire N__19574;
    wire N__19571;
    wire N__19568;
    wire N__19565;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19553;
    wire N__19550;
    wire N__19547;
    wire N__19544;
    wire N__19541;
    wire N__19540;
    wire N__19539;
    wire N__19538;
    wire N__19537;
    wire N__19536;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19525;
    wire N__19522;
    wire N__19519;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19507;
    wire N__19498;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19482;
    wire N__19479;
    wire N__19476;
    wire N__19473;
    wire N__19466;
    wire N__19463;
    wire N__19460;
    wire N__19457;
    wire N__19454;
    wire N__19451;
    wire N__19448;
    wire N__19445;
    wire N__19442;
    wire N__19439;
    wire N__19436;
    wire N__19433;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19423;
    wire N__19420;
    wire N__19417;
    wire N__19414;
    wire N__19409;
    wire N__19406;
    wire N__19405;
    wire N__19400;
    wire N__19397;
    wire N__19394;
    wire N__19391;
    wire N__19388;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19349;
    wire N__19346;
    wire N__19343;
    wire N__19340;
    wire N__19337;
    wire N__19334;
    wire N__19331;
    wire N__19328;
    wire N__19325;
    wire N__19322;
    wire N__19319;
    wire N__19316;
    wire N__19313;
    wire N__19310;
    wire N__19307;
    wire N__19304;
    wire N__19301;
    wire N__19298;
    wire N__19295;
    wire N__19292;
    wire N__19289;
    wire N__19286;
    wire N__19283;
    wire N__19280;
    wire N__19277;
    wire N__19274;
    wire N__19271;
    wire N__19268;
    wire N__19265;
    wire N__19262;
    wire N__19259;
    wire N__19256;
    wire N__19253;
    wire N__19250;
    wire N__19247;
    wire N__19244;
    wire N__19241;
    wire N__19238;
    wire N__19235;
    wire N__19232;
    wire N__19229;
    wire N__19226;
    wire N__19223;
    wire N__19220;
    wire N__19217;
    wire N__19214;
    wire N__19211;
    wire N__19208;
    wire N__19205;
    wire N__19202;
    wire N__19199;
    wire N__19196;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire N__19178;
    wire N__19175;
    wire N__19172;
    wire N__19169;
    wire N__19166;
    wire N__19163;
    wire N__19160;
    wire N__19157;
    wire N__19154;
    wire N__19151;
    wire N__19148;
    wire N__19145;
    wire N__19142;
    wire N__19139;
    wire N__19136;
    wire N__19133;
    wire N__19130;
    wire N__19129;
    wire N__19128;
    wire N__19125;
    wire N__19124;
    wire N__19123;
    wire N__19116;
    wire N__19113;
    wire N__19110;
    wire N__19105;
    wire N__19100;
    wire N__19097;
    wire N__19094;
    wire N__19091;
    wire N__19088;
    wire N__19085;
    wire N__19082;
    wire N__19079;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19058;
    wire N__19055;
    wire N__19052;
    wire N__19049;
    wire N__19046;
    wire N__19043;
    wire N__19040;
    wire N__19037;
    wire N__19034;
    wire N__19031;
    wire N__19028;
    wire N__19025;
    wire N__19022;
    wire N__19019;
    wire N__19016;
    wire N__19013;
    wire N__19010;
    wire N__19007;
    wire N__19004;
    wire N__19001;
    wire N__18998;
    wire N__18995;
    wire N__18992;
    wire N__18989;
    wire N__18986;
    wire N__18983;
    wire N__18980;
    wire N__18977;
    wire N__18974;
    wire N__18971;
    wire N__18968;
    wire N__18965;
    wire N__18962;
    wire N__18959;
    wire N__18956;
    wire N__18953;
    wire N__18950;
    wire N__18947;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18935;
    wire N__18932;
    wire N__18929;
    wire N__18926;
    wire N__18923;
    wire N__18920;
    wire N__18917;
    wire N__18914;
    wire N__18911;
    wire N__18908;
    wire N__18905;
    wire N__18902;
    wire N__18899;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18866;
    wire N__18863;
    wire N__18860;
    wire N__18857;
    wire N__18854;
    wire N__18851;
    wire N__18848;
    wire N__18845;
    wire N__18844;
    wire N__18843;
    wire N__18840;
    wire N__18835;
    wire N__18832;
    wire N__18827;
    wire N__18826;
    wire N__18825;
    wire N__18822;
    wire N__18819;
    wire N__18816;
    wire N__18811;
    wire N__18808;
    wire N__18805;
    wire N__18802;
    wire N__18797;
    wire N__18796;
    wire N__18793;
    wire N__18790;
    wire N__18787;
    wire N__18782;
    wire N__18779;
    wire N__18778;
    wire N__18775;
    wire N__18772;
    wire N__18769;
    wire N__18764;
    wire N__18761;
    wire N__18760;
    wire N__18757;
    wire N__18754;
    wire N__18751;
    wire N__18746;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18734;
    wire N__18733;
    wire N__18728;
    wire N__18725;
    wire N__18722;
    wire N__18719;
    wire N__18716;
    wire N__18713;
    wire N__18710;
    wire N__18707;
    wire N__18704;
    wire N__18701;
    wire N__18700;
    wire N__18695;
    wire N__18692;
    wire N__18689;
    wire N__18686;
    wire N__18683;
    wire N__18680;
    wire N__18677;
    wire N__18674;
    wire N__18671;
    wire N__18668;
    wire N__18667;
    wire N__18664;
    wire N__18661;
    wire N__18656;
    wire N__18653;
    wire N__18650;
    wire N__18647;
    wire N__18646;
    wire N__18645;
    wire N__18638;
    wire N__18635;
    wire N__18632;
    wire N__18629;
    wire N__18626;
    wire N__18625;
    wire N__18622;
    wire N__18619;
    wire N__18618;
    wire N__18613;
    wire N__18610;
    wire N__18605;
    wire N__18602;
    wire N__18601;
    wire N__18596;
    wire N__18593;
    wire N__18590;
    wire N__18587;
    wire N__18584;
    wire N__18581;
    wire N__18578;
    wire N__18575;
    wire N__18572;
    wire N__18569;
    wire N__18566;
    wire N__18563;
    wire N__18560;
    wire N__18557;
    wire N__18554;
    wire N__18551;
    wire N__18548;
    wire N__18545;
    wire N__18542;
    wire N__18539;
    wire N__18536;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18482;
    wire N__18479;
    wire N__18476;
    wire delay_tr_input_ibuf_gb_io_gb_input;
    wire delay_hc_input_ibuf_gb_io_gb_input;
    wire GNDG0;
    wire VCCG0;
    wire \pll_inst.red_c_i ;
    wire bfn_1_14_0_;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_0 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_1 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_2 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_3 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_4 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_5 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_7 ;
    wire bfn_1_15_0_;
    wire \pwm_generator_inst.un3_threshold_acc_cry_8 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_9 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_10 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_11 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_12 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_13 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_15 ;
    wire bfn_1_16_0_;
    wire \pwm_generator_inst.un3_threshold_acc_cry_16 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_17 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_19 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_ ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_ ;
    wire N_38_i_i;
    wire rgb_drv_RNOZ0;
    wire \pwm_generator_inst.un2_threshold_acc_2_1_15 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1_16 ;
    wire \current_shift_inst.PI_CTRL.N_154 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_3 ;
    wire pwm_duty_input_4;
    wire pwm_duty_input_3;
    wire pwm_duty_input_0;
    wire pwm_duty_input_1;
    wire pwm_duty_input_2;
    wire \pwm_generator_inst.un1_duty_inputlt3 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire \current_shift_inst.PI_CTRL.N_31_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_149 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_27 ;
    wire \current_shift_inst.PI_CTRL.N_27_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_153 ;
    wire \current_shift_inst.PI_CTRL.N_155 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_15 ;
    wire \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ;
    wire bfn_2_13_0_;
    wire \pwm_generator_inst.un2_threshold_acc_2_1 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_16 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_2 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_17 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_18 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_19 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_20 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_21 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_6 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_22 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_23 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ;
    wire bfn_2_14_0_;
    wire \pwm_generator_inst.un2_threshold_acc_2_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_24 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_14 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_25 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ;
    wire bfn_2_15_0_;
    wire \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_ ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_ ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_14_cascade_ ;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_0 ;
    wire bfn_2_16_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_2 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_7 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_8 ;
    wire bfn_2_17_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_9 ;
    wire \pwm_generator_inst.un3_threshold_acc ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_12 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_11 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_12 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_14 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_13 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_15 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_14 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_15 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_16 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ;
    wire bfn_2_18_0_;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_17 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_16 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_17 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_18 ;
    wire \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_5 ;
    wire pwm_duty_input_8;
    wire pwm_duty_input_9;
    wire pwm_duty_input_6;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ;
    wire pwm_duty_input_7;
    wire pwm_duty_input_5;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_53 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ;
    wire \current_shift_inst.PI_CTRL.N_118 ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_3_12_0_;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.thresholdZ0Z_5 ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_3_13_0_;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire \pwm_generator_inst.thresholdZ0Z_0 ;
    wire \pwm_generator_inst.thresholdZ0Z_1 ;
    wire \pwm_generator_inst.thresholdZ0Z_4 ;
    wire \pwm_generator_inst.thresholdZ0Z_6 ;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_0 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_6 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_7 ;
    wire \pwm_generator_inst.thresholdZ0Z_7 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_4 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_1 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_0 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ;
    wire bfn_3_17_0_;
    wire \pwm_generator_inst.un19_threshold_acc_axb_1 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_0 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_2 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_1 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_2 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_4 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_3 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_5 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_4 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_6 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_5 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_7 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_6 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_7 ;
    wire bfn_3_18_0_;
    wire \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_8 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_18 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_8 ;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ;
    wire \pwm_generator_inst.un1_counterlto2_0_cascade_ ;
    wire \pwm_generator_inst.un1_counterlto9_2_cascade_ ;
    wire \pwm_generator_inst.un1_counterlt9 ;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire bfn_4_13_0_;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire bfn_4_14_0_;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire \pwm_generator_inst.thresholdZ0Z_2 ;
    wire \pwm_generator_inst.thresholdZ0Z_9 ;
    wire \pwm_generator_inst.thresholdZ0Z_3 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_2 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_3 ;
    wire \pwm_generator_inst.thresholdZ0Z_8 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_8 ;
    wire \pwm_generator_inst.N_16 ;
    wire \pwm_generator_inst.N_17 ;
    wire N_19_1;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_13 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_3 ;
    wire il_max_comp2_c;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire bfn_5_9_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire bfn_5_10_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire bfn_5_11_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire bfn_5_12_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire il_max_comp2_D1;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_16_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_20_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_75_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31 ;
    wire \current_shift_inst.PI_CTRL.N_62 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_7_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_18 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire bfn_7_13_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire bfn_7_14_0_;
    wire \phase_controller_inst1.stoper_hc.un6_running_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_16 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_17 ;
    wire bfn_7_15_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_19 ;
    wire \phase_controller_inst2.start_timer_hc_0_sqmuxa_cascade_ ;
    wire \phase_controller_inst2.start_timer_hc_RNOZ0Z_0 ;
    wire \phase_controller_inst2.stoper_hc.un2_start_0_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ;
    wire \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.un2_start_0 ;
    wire il_max_comp1_c;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ;
    wire \current_shift_inst.PI_CTRL.N_74_16 ;
    wire \current_shift_inst.PI_CTRL.N_74_21 ;
    wire \current_shift_inst.PI_CTRL.N_103_cascade_ ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire bfn_8_13_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire bfn_8_14_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire bfn_8_15_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.running_1_sqmuxa ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ;
    wire \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNIQVTIZ0Z1 ;
    wire \phase_controller_inst1.stoper_hc.runningZ0 ;
    wire \phase_controller_inst1.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_6 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_2 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_4 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_5 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_8 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_3 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_1 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ;
    wire bfn_8_19_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNINJBZ0Z21 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ;
    wire bfn_8_20_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ;
    wire bfn_8_21_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.N_434_i ;
    wire bfn_9_8_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_0 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_3 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_2 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_5 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire bfn_9_9_0_;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_14 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire bfn_9_10_0_;
    wire \current_shift_inst.PI_CTRL.integrator_i_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire bfn_9_11_0_;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_29 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_30 ;
    wire bfn_9_12_0_;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_15 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_22 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_9 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_13 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_19 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_18 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_17 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_16 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_15 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_7 ;
    wire \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ;
    wire elapsed_time_ns_1_RNI62CED1_0_19_cascade_;
    wire \phase_controller_inst1.stoper_hc.N_315_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18_cascade_ ;
    wire elapsed_time_ns_1_RNIQ4OD11_0_31_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_time_4_f0_i_1Z0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_f0_i_1Z0Z_9_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.N_315 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.N_283_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.N_307 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6_cascade_ ;
    wire elapsed_time_ns_1_RNIIU2KD1_0_6;
    wire elapsed_time_ns_1_RNIIU2KD1_0_6_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0Z0Z_6_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_ ;
    wire elapsed_time_ns_1_RNIDP2KD1_0_1;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.N_327 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_1 ;
    wire bfn_9_19_0_;
    wire \phase_controller_inst2.stoper_hc.un6_running_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_6 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_9 ;
    wire bfn_9_20_0_;
    wire \phase_controller_inst2.stoper_hc.un6_running_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_14 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_16 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_17 ;
    wire bfn_9_21_0_;
    wire \phase_controller_inst2.stoper_hc.un6_running_18 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_17 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_19 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_19 ;
    wire s3_phy_c;
    wire \current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3 ;
    wire \current_shift_inst.PI_CTRL.N_72 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_2 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc5_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0 ;
    wire elapsed_time_ns_1_RNIL13KD1_0_9_cascade_;
    wire elapsed_time_ns_1_RNI1BND11_0_29;
    wire elapsed_time_ns_1_RNI1BND11_0_29_cascade_;
    wire elapsed_time_ns_1_RNIT6ND11_0_25;
    wire elapsed_time_ns_1_RNI0AND11_0_28;
    wire elapsed_time_ns_1_RNIV8ND11_0_27;
    wire elapsed_time_ns_1_RNIT6ND11_0_25_cascade_;
    wire elapsed_time_ns_1_RNIU7ND11_0_26;
    wire elapsed_time_ns_1_RNIP2ND11_0_21;
    wire elapsed_time_ns_1_RNIS5ND11_0_24;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.un6_running_17 ;
    wire elapsed_time_ns_1_RNIQ3ND11_0_22;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17_cascade_ ;
    wire elapsed_time_ns_1_RNIR4ND11_0_23;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa ;
    wire elapsed_time_ns_1_RNI3VBED1_0_16_cascade_;
    wire elapsed_time_ns_1_RNIA3DJ11_0_4;
    wire elapsed_time_ns_1_RNI40CED1_0_17;
    wire elapsed_time_ns_1_RNIA3DJ11_0_4_cascade_;
    wire elapsed_time_ns_1_RNI51CED1_0_18;
    wire elapsed_time_ns_1_RNI62CED1_0_19;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.N_328 ;
    wire \phase_controller_inst1.stoper_hc.N_337 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_4 ;
    wire elapsed_time_ns_1_RNIQURR91_0_3;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_5 ;
    wire elapsed_time_ns_1_RNINVLD11_0_10;
    wire elapsed_time_ns_1_RNIQ2MD11_0_13;
    wire elapsed_time_ns_1_RNINVLD11_0_10_cascade_;
    wire elapsed_time_ns_1_RNIP1MD11_0_12;
    wire \phase_controller_inst1.stoper_hc.N_319_cascade_ ;
    wire elapsed_time_ns_1_RNI1TBED1_0_14;
    wire \phase_controller_inst1.stoper_hc.N_275 ;
    wire \phase_controller_inst1.stoper_hc.N_319 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a5_1_0Z0Z_9 ;
    wire elapsed_time_ns_1_RNIQ4OD11_0_31;
    wire \phase_controller_inst1.stoper_hc.N_278 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_15 ;
    wire \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ;
    wire elapsed_time_ns_1_RNID6DJ11_0_7;
    wire elapsed_time_ns_1_RNIE7DJ11_0_8;
    wire elapsed_time_ns_1_RNIB4DJ11_0_5;
    wire elapsed_time_ns_1_RNIS4MD11_0_15;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_CO ;
    wire \phase_controller_inst2.stoper_hc.running_1_sqmuxa ;
    wire \phase_controller_inst2.start_timer_hcZ0 ;
    wire \phase_controller_inst2.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst2.stoper_hc.running_1_sqmuxa_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.runningZ0 ;
    wire \phase_controller_inst2.stoper_hc.un1_start_latched2_0 ;
    wire s4_phy_c;
    wire il_max_comp1_D1;
    wire il_min_comp2_c;
    wire il_min_comp2_D1;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_19 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.N_103 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ;
    wire bfn_11_10_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_6 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_8 ;
    wire bfn_11_11_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO ;
    wire bfn_11_12_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO ;
    wire bfn_11_13_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_31 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.N_382_i_cascade_ ;
    wire elapsed_time_ns_1_RNIP3OD11_0_30;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91Z0Z_7_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2Z0Z_15_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719Z0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992Z0Z_24 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9Z0Z_24 ;
    wire bfn_11_15_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire bfn_11_16_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire bfn_11_17_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire bfn_11_18_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire bfn_11_19_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire bfn_11_20_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_11_21_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire bfn_11_22_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \delay_measurement_inst.delay_hc_timer.N_432_i ;
    wire il_min_comp1_c;
    wire il_min_comp1_D1;
    wire delay_hc_input_c_g;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_1 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_i_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_24 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_8 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_21 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axb_0 ;
    wire bfn_12_11_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_1 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_2 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_3 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_4 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_5 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_7 ;
    wire bfn_12_12_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_9 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_11 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_8 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ;
    wire elapsed_time_ns_1_RNIO0MD11_0_11;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc5lto15 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKRZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847Z0Z_31 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4Z0Z_31 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_a3_1_3 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_6_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_5 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58FZ0Z_31 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc5lto14 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc5lto6 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2 ;
    wire T01_c;
    wire T12_c;
    wire \phase_controller_inst2.stateZ0Z_2 ;
    wire \phase_controller_inst2.hc_time_passed ;
    wire il_max_comp2_D2;
    wire \phase_controller_inst2.time_passed_RNI9M3O_cascade_ ;
    wire \phase_controller_inst2.time_passed_RNI9M3O ;
    wire T23_c;
    wire \phase_controller_inst2.stateZ0Z_3 ;
    wire \phase_controller_inst2.stateZ0Z_0 ;
    wire T45_c;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.N_433_i ;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire bfn_13_5_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire bfn_13_6_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire bfn_13_7_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire bfn_13_8_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire bfn_13_9_0_;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire bfn_13_10_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire bfn_13_11_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire bfn_13_12_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.N_435_i ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.un2_start_0_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.running_1_sqmuxa_cascade_ ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire delay_tr_input_c_g;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_12 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_i_0_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ;
    wire \phase_controller_inst2.stateZ0Z_1 ;
    wire il_min_comp2_D2;
    wire \phase_controller_inst2.start_timer_tr_0_sqmuxa ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ;
    wire elapsed_time_ns_1_RNI3VBED1_0_16;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16 ;
    wire start_stop_c;
    wire \current_shift_inst.elapsed_time_ns_s1_fast_31 ;
    wire s2_phy_c;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.delay_tr_timer.N_359_1_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_345 ;
    wire \delay_measurement_inst.delay_tr_timer.N_345_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5 ;
    wire \delay_measurement_inst.delay_tr_timer.N_341 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ;
    wire \delay_measurement_inst.delay_tr_timer.N_434_i_g ;
    wire \delay_measurement_inst.delay_tr_timer.N_348 ;
    wire \delay_measurement_inst.delay_tr_timer.N_367 ;
    wire \delay_measurement_inst.delay_tr_timer.N_349_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_363_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_380 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_378 ;
    wire \delay_measurement_inst.delay_tr_timer.N_359_1 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8 ;
    wire \delay_measurement_inst.delay_tr_timer.N_347 ;
    wire \delay_measurement_inst.delay_tr_timer.N_347_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_365 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_7 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire elapsed_time_ns_1_RNITCIF91_0_23;
    wire elapsed_time_ns_1_RNITCIF91_0_23_cascade_;
    wire elapsed_time_ns_1_RNIUDIF91_0_24;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ;
    wire \phase_controller_inst1.N_55_cascade_ ;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire \phase_controller_inst1.start_timer_tr_0_sqmuxa_cascade_ ;
    wire phase_controller_inst1_state_4;
    wire \phase_controller_inst2.stoper_tr.un1_start_latched2_0 ;
    wire \phase_controller_inst2.tr_time_passed ;
    wire \phase_controller_inst2.stoper_tr.running_1_sqmuxa ;
    wire \phase_controller_inst2.stoper_tr.runningZ0 ;
    wire \phase_controller_inst2.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst2.start_timer_trZ0 ;
    wire \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ;
    wire \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.un2_start_0 ;
    wire bfn_14_14_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s0 ;
    wire \current_shift_inst.un38_control_input_cry_1_s0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_2_s0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0 ;
    wire bfn_14_15_0_;
    wire \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_8_s0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0 ;
    wire bfn_14_16_0_;
    wire \current_shift_inst.un38_control_input_cry_16_s0 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ;
    wire \current_shift_inst.un38_control_input_cry_20_s0 ;
    wire \current_shift_inst.un38_control_input_cry_21_s0 ;
    wire \current_shift_inst.un38_control_input_cry_22_s0 ;
    wire \current_shift_inst.un38_control_input_cry_23_s0 ;
    wire bfn_14_17_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ;
    wire \current_shift_inst.un38_control_input_cry_24_s0 ;
    wire \current_shift_inst.un38_control_input_cry_25_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ;
    wire \current_shift_inst.un38_control_input_cry_26_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ;
    wire \current_shift_inst.un38_control_input_cry_27_s0 ;
    wire \current_shift_inst.un38_control_input_cry_28_s0 ;
    wire \current_shift_inst.un38_control_input_cry_29_s0 ;
    wire \current_shift_inst.un38_control_input_axb_31_s0 ;
    wire \current_shift_inst.un38_control_input_cry_30_s0 ;
    wire \current_shift_inst.un38_control_input_5_0 ;
    wire bfn_14_18_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1 ;
    wire bfn_14_19_0_;
    wire \current_shift_inst.un38_control_input_cry_8_s1 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1 ;
    wire bfn_14_20_0_;
    wire \current_shift_inst.un38_control_input_cry_16_s1 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ;
    wire \current_shift_inst.un38_control_input_cry_20_s1 ;
    wire \current_shift_inst.un38_control_input_cry_21_s1 ;
    wire \current_shift_inst.un38_control_input_cry_22_s1 ;
    wire \current_shift_inst.un38_control_input_cry_23_s1 ;
    wire bfn_14_21_0_;
    wire \current_shift_inst.un38_control_input_cry_24_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ;
    wire \current_shift_inst.un38_control_input_cry_25_s1 ;
    wire \current_shift_inst.un38_control_input_cry_26_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ;
    wire \current_shift_inst.un38_control_input_cry_27_s1 ;
    wire \current_shift_inst.un38_control_input_cry_28_s1 ;
    wire \current_shift_inst.un38_control_input_cry_29_s1 ;
    wire \current_shift_inst.un38_control_input_cry_30_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_31 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ;
    wire \delay_measurement_inst.delay_tr_timer.N_381 ;
    wire \delay_measurement_inst.delay_tr_timer.N_358 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ;
    wire elapsed_time_ns_1_RNIIJ4DM1_0_19_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ;
    wire elapsed_time_ns_1_RNISAHF91_0_13_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire elapsed_time_ns_1_RNIVEIF91_0_25;
    wire elapsed_time_ns_1_RNI1HIF91_0_27;
    wire elapsed_time_ns_1_RNIVEIF91_0_25_cascade_;
    wire elapsed_time_ns_1_RNI0GIF91_0_26;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire elapsed_time_ns_1_RNI2IIF91_0_28;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_1 ;
    wire bfn_15_10_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_9 ;
    wire bfn_15_11_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_17 ;
    wire bfn_15_12_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_19 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc5 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc5lto9 ;
    wire elapsed_time_ns_1_RNIL13KD1_0_9;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ;
    wire bfn_15_13_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNI2FGQZ0Z1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ;
    wire bfn_15_14_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ;
    wire bfn_15_15_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_start_latched2_0 ;
    wire \phase_controller_inst1.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire \phase_controller_inst1.hc_time_passed ;
    wire \current_shift_inst.control_inputZ0Z_0 ;
    wire bfn_15_16_0_;
    wire \current_shift_inst.control_inputZ0Z_1 ;
    wire \current_shift_inst.control_input_1_cry_0 ;
    wire \current_shift_inst.control_inputZ0Z_2 ;
    wire \current_shift_inst.control_input_1_cry_1 ;
    wire \current_shift_inst.control_inputZ0Z_3 ;
    wire \current_shift_inst.control_input_1_cry_2 ;
    wire \current_shift_inst.control_inputZ0Z_4 ;
    wire \current_shift_inst.control_input_1_cry_3 ;
    wire \current_shift_inst.control_inputZ0Z_5 ;
    wire \current_shift_inst.control_input_1_cry_4 ;
    wire \current_shift_inst.control_inputZ0Z_6 ;
    wire \current_shift_inst.control_input_1_cry_5 ;
    wire \current_shift_inst.control_inputZ0Z_7 ;
    wire \current_shift_inst.control_input_1_cry_6 ;
    wire \current_shift_inst.control_input_1_cry_7 ;
    wire \current_shift_inst.control_inputZ0Z_8 ;
    wire bfn_15_17_0_;
    wire \current_shift_inst.control_inputZ0Z_9 ;
    wire \current_shift_inst.control_input_1_cry_8 ;
    wire \current_shift_inst.control_inputZ0Z_10 ;
    wire \current_shift_inst.control_input_1_cry_9 ;
    wire \current_shift_inst.control_input_1_axb_11 ;
    wire \current_shift_inst.control_input_1_cry_10 ;
    wire \current_shift_inst.control_inputZ0Z_11 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ;
    wire \current_shift_inst.N_1609_i ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ;
    wire \current_shift_inst.un38_control_input_0_s0_27 ;
    wire \current_shift_inst.un38_control_input_0_s1_27 ;
    wire \current_shift_inst.control_input_1_axb_7 ;
    wire \current_shift_inst.un38_control_input_0_s1_28 ;
    wire \current_shift_inst.un38_control_input_0_s0_28 ;
    wire \current_shift_inst.control_input_1_axb_8 ;
    wire \current_shift_inst.un38_control_input_0_s0_29 ;
    wire \current_shift_inst.un38_control_input_0_s1_29 ;
    wire \current_shift_inst.control_input_1_axb_9 ;
    wire \current_shift_inst.un38_control_input_0_s1_30 ;
    wire \current_shift_inst.un38_control_input_0_s0_30 ;
    wire \current_shift_inst.control_input_1_axb_10 ;
    wire elapsed_time_ns_1_RNI81DJ11_0_2;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ;
    wire \delay_measurement_inst.delay_hc_timer.N_432_i_g ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire \delay_measurement_inst.delay_hc_timer.N_382_i ;
    wire elapsed_time_ns_1_RNIO1ND11_0_20;
    wire \current_shift_inst.un38_control_input_0_s0_20 ;
    wire \current_shift_inst.un38_control_input_0_s1_20 ;
    wire \current_shift_inst.control_input_1_axb_0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ;
    wire \current_shift_inst.un38_control_input_0_s0_21 ;
    wire \current_shift_inst.un38_control_input_0_s1_21 ;
    wire \current_shift_inst.control_input_1_axb_1 ;
    wire \current_shift_inst.un38_control_input_0_s0_22 ;
    wire \current_shift_inst.un38_control_input_0_s1_22 ;
    wire \current_shift_inst.control_input_1_axb_2 ;
    wire \current_shift_inst.un38_control_input_0_s1_23 ;
    wire \current_shift_inst.un38_control_input_0_s0_23 ;
    wire \current_shift_inst.control_input_1_axb_3 ;
    wire \current_shift_inst.un38_control_input_0_s1_24 ;
    wire \current_shift_inst.un38_control_input_0_s0_24 ;
    wire \current_shift_inst.control_input_1_axb_4 ;
    wire \current_shift_inst.un38_control_input_0_s1_25 ;
    wire \current_shift_inst.un38_control_input_0_s0_25 ;
    wire \current_shift_inst.control_input_1_axb_5 ;
    wire \current_shift_inst.un38_control_input_0_s0_26 ;
    wire \current_shift_inst.un38_control_input_0_s1_26 ;
    wire \current_shift_inst.control_input_1_axb_6 ;
    wire \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ;
    wire \current_shift_inst.timer_s1.N_166_i ;
    wire s1_phy_c;
    wire state_ns_i_a3_1;
    wire state_3;
    wire il_max_comp1_D2;
    wire \phase_controller_inst1.start_timer_hc_0_sqmuxa ;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17_cascade_ ;
    wire elapsed_time_ns_1_RNIGH4DM1_0_17_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ;
    wire elapsed_time_ns_1_RNICG2591_0_4_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2_cascade_ ;
    wire elapsed_time_ns_1_RNIDE4DM1_0_14_cascade_;
    wire \phase_controller_inst1.stoper_tr.N_241_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.un6_running_14 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_10 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_11 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_12 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_13 ;
    wire elapsed_time_ns_1_RNISAHF91_0_13;
    wire elapsed_time_ns_1_RNIQ8HF91_0_11;
    wire elapsed_time_ns_1_RNIP7HF91_0_10;
    wire elapsed_time_ns_1_RNIR9HF91_0_12;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire elapsed_time_ns_1_RNIRAIF91_0_21;
    wire elapsed_time_ns_1_RNIRBJF91_0_30;
    wire elapsed_time_ns_1_RNI3JIF91_0_29;
    wire elapsed_time_ns_1_RNIRAIF91_0_21_cascade_;
    wire elapsed_time_ns_1_RNIQ9IF91_0_20;
    wire elapsed_time_ns_1_RNISBIF91_0_22;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18 ;
    wire elapsed_time_ns_1_RNIHI4DM1_0_18;
    wire elapsed_time_ns_1_RNIHI4DM1_0_18_cascade_;
    wire \phase_controller_inst2.stoper_tr.un6_running_18 ;
    wire elapsed_time_ns_1_RNIGH4DM1_0_17;
    wire \phase_controller_inst2.stoper_tr.un6_running_17 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9 ;
    wire elapsed_time_ns_1_RNISCJF91_0_31_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.N_241 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.un6_running_9 ;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire il_min_comp1_D2;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire \phase_controller_inst1.N_56 ;
    wire \phase_controller_inst1.tr_time_passed ;
    wire \current_shift_inst.un38_control_input_cry_0_s0_sf ;
    wire \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ;
    wire bfn_16_16_0_;
    wire \current_shift_inst.un10_control_input_cry_0 ;
    wire \current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_1 ;
    wire \current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_2 ;
    wire \current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_3 ;
    wire \current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_4 ;
    wire \current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_5 ;
    wire \current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_6 ;
    wire \current_shift_inst.un10_control_input_cry_7 ;
    wire \current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ;
    wire bfn_16_17_0_;
    wire \current_shift_inst.un10_control_input_cry_8 ;
    wire \current_shift_inst.un10_control_input_cry_9 ;
    wire \current_shift_inst.un10_control_input_cry_10 ;
    wire \current_shift_inst.un10_control_input_cry_11 ;
    wire \current_shift_inst.un10_control_input_cry_12 ;
    wire \current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_13 ;
    wire \current_shift_inst.un10_control_input_cry_14 ;
    wire \current_shift_inst.un10_control_input_cry_15 ;
    wire bfn_16_18_0_;
    wire \current_shift_inst.un10_control_input_cry_16 ;
    wire \current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_17 ;
    wire \current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_18 ;
    wire \current_shift_inst.un10_control_input_cry_19 ;
    wire \current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_20 ;
    wire \current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_21 ;
    wire \current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_22 ;
    wire \current_shift_inst.un10_control_input_cry_23 ;
    wire bfn_16_19_0_;
    wire \current_shift_inst.un10_control_input_cry_24 ;
    wire \current_shift_inst.un10_control_input_cry_25 ;
    wire \current_shift_inst.un10_control_input_cry_26 ;
    wire \current_shift_inst.un10_control_input_cry_27 ;
    wire \current_shift_inst.un10_control_input_cry_28 ;
    wire CONSTANT_ONE_NET;
    wire \current_shift_inst.un10_control_input_cry_29 ;
    wire \current_shift_inst.un10_control_input_cry_30 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ;
    wire bfn_16_21_0_;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire bfn_16_22_0_;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire bfn_16_23_0_;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire bfn_16_24_0_;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.running_i ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire \current_shift_inst.timer_s1.N_167_i ;
    wire elapsed_time_ns_1_RNIIJ4DM1_0_19;
    wire \phase_controller_inst2.stoper_tr.un6_running_19 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_16 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_15 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_7 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_8 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_2 ;
    wire \phase_controller_inst1.stoper_tr.N_219 ;
    wire elapsed_time_ns_1_RNIAE2591_0_2;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1Z0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6 ;
    wire elapsed_time_ns_1_RNIGK2591_0_8;
    wire elapsed_time_ns_1_RNIUKL2M1_0_6_cascade_;
    wire \phase_controller_inst1.stoper_tr.N_247 ;
    wire \phase_controller_inst1.stoper_tr.N_247_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.un6_running_6 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto15 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ;
    wire elapsed_time_ns_1_RNIUCHF91_0_15_cascade_;
    wire \phase_controller_inst1.stoper_tr.N_251 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9 ;
    wire elapsed_time_ns_1_RNI1OL2M1_0_9;
    wire elapsed_time_ns_1_RNIDE4DM1_0_14;
    wire elapsed_time_ns_1_RNI1OL2M1_0_9_cascade_;
    wire \phase_controller_inst1.stoper_tr.N_244 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2Z0Z_9 ;
    wire elapsed_time_ns_1_RNIUCHF91_0_15;
    wire \phase_controller_inst1.stoper_tr.N_211_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_0_6_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.un6_running_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_17_10_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_17_11_0_;
    wire \phase_controller_inst1.stoper_tr.un6_running_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_17 ;
    wire bfn_17_12_0_;
    wire \phase_controller_inst1.stoper_tr.un6_running_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_19 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_28 ;
    wire \current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_1 ;
    wire \current_shift_inst.un4_control_input1_1_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_30 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_13 ;
    wire \current_shift_inst.elapsed_time_ns_s1_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1 ;
    wire bfn_17_15_0_;
    wire \current_shift_inst.un4_control_input1_3 ;
    wire \current_shift_inst.un4_control_input_1_cry_1 ;
    wire \current_shift_inst.un4_control_input1_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_2 ;
    wire \current_shift_inst.un4_control_input_1_axb_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_3 ;
    wire \current_shift_inst.un4_control_input_1_axb_5 ;
    wire \current_shift_inst.un4_control_input1_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_4 ;
    wire \current_shift_inst.un4_control_input1_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_5 ;
    wire \current_shift_inst.un4_control_input1_8 ;
    wire \current_shift_inst.un4_control_input_1_cry_6 ;
    wire \current_shift_inst.un4_control_input1_9 ;
    wire \current_shift_inst.un4_control_input_1_cry_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_8 ;
    wire bfn_17_16_0_;
    wire \current_shift_inst.un4_control_input_1_cry_9 ;
    wire \current_shift_inst.un4_control_input_1_cry_10 ;
    wire \current_shift_inst.un4_control_input_1_cry_11 ;
    wire \current_shift_inst.un4_control_input_1_cry_12 ;
    wire \current_shift_inst.un4_control_input_1_cry_13 ;
    wire \current_shift_inst.un4_control_input_1_cry_14 ;
    wire \current_shift_inst.un4_control_input_1_cry_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_16 ;
    wire bfn_17_17_0_;
    wire \current_shift_inst.un4_control_input_1_cry_17 ;
    wire \current_shift_inst.un4_control_input1_20 ;
    wire \current_shift_inst.un4_control_input_1_cry_18 ;
    wire \current_shift_inst.un4_control_input_1_cry_19 ;
    wire \current_shift_inst.un4_control_input1_22 ;
    wire \current_shift_inst.un4_control_input_1_cry_20 ;
    wire \current_shift_inst.un4_control_input1_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_21 ;
    wire \current_shift_inst.un4_control_input1_24 ;
    wire \current_shift_inst.un4_control_input_1_cry_22 ;
    wire \current_shift_inst.un4_control_input_1_cry_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_24 ;
    wire bfn_17_18_0_;
    wire \current_shift_inst.un4_control_input_1_cry_25 ;
    wire \current_shift_inst.un4_control_input1_28 ;
    wire \current_shift_inst.un4_control_input_1_cry_26 ;
    wire \current_shift_inst.un4_control_input_1_cry_27 ;
    wire \current_shift_inst.un4_control_input_1_cry_28 ;
    wire \current_shift_inst.un4_control_input1_31 ;
    wire \current_shift_inst.un4_control_input1_21 ;
    wire \current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_29 ;
    wire \current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_12 ;
    wire \current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_12 ;
    wire \current_shift_inst.un4_control_input1_19 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_21 ;
    wire \current_shift_inst.un4_control_input_1_axb_10 ;
    wire \current_shift_inst.un4_control_input_1_axb_14 ;
    wire \current_shift_inst.un4_control_input_1_axb_18 ;
    wire \current_shift_inst.un4_control_input_1_axb_26 ;
    wire \current_shift_inst.un4_control_input_1_axb_15 ;
    wire \current_shift_inst.un4_control_input_1_axb_24 ;
    wire \current_shift_inst.un4_control_input_1_axb_16 ;
    wire \current_shift_inst.un4_control_input_1_axb_25 ;
    wire \current_shift_inst.un4_control_input_1_axb_23 ;
    wire \current_shift_inst.un4_control_input_1_axb_28 ;
    wire \current_shift_inst.un4_control_input_1_axb_29 ;
    wire \current_shift_inst.un4_control_input_1_axb_27 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ;
    wire elapsed_time_ns_1_RNIFG4DM1_0_16;
    wire \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1 ;
    wire elapsed_time_ns_1_RNIPFL2M1_0_1;
    wire \phase_controller_inst1.stoper_tr.N_235 ;
    wire elapsed_time_ns_1_RNIPFL2M1_0_1_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_1 ;
    wire elapsed_time_ns_1_RNIUKL2M1_0_6;
    wire \phase_controller_inst1.stoper_tr.un6_running_6 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_2 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_4 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_5 ;
    wire elapsed_time_ns_1_RNIFJ2591_0_7;
    wire \phase_controller_inst1.stoper_tr.un6_running_7 ;
    wire elapsed_time_ns_1_RNICG2591_0_4;
    wire \phase_controller_inst2.stoper_tr.un6_running_4 ;
    wire elapsed_time_ns_1_RNISCJF91_0_31;
    wire elapsed_time_ns_1_RNIDH2591_0_5;
    wire \phase_controller_inst2.stoper_tr.un6_running_5 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_0_6 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ;
    wire elapsed_time_ns_1_RNIRHL2M1_0_3;
    wire \phase_controller_inst2.stoper_tr.un6_running_3 ;
    wire \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.running_1_sqmuxa ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst1.stoper_tr.running_1_sqmuxa_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.runningZ0 ;
    wire \phase_controller_inst1.stoper_tr.un1_start_latched2_0 ;
    wire \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ;
    wire \phase_controller_inst1.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire bfn_18_11_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNISF8IZ0Z2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire bfn_18_12_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire bfn_18_13_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \current_shift_inst.un4_control_input1_5 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_20 ;
    wire \current_shift_inst.un4_control_input1_17 ;
    wire \current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_18 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_13 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_15 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_16 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_3 ;
    wire \current_shift_inst.un4_control_input_1_axb_7 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_10 ;
    wire \current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_2 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ;
    wire \current_shift_inst.un4_control_input_1_axb_1 ;
    wire \current_shift_inst.un38_control_input_5_1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO ;
    wire \current_shift_inst.un4_control_input_0_31 ;
    wire \current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ;
    wire \current_shift_inst.un4_control_input_1_axb_11 ;
    wire \current_shift_inst.un4_control_input1_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ;
    wire \current_shift_inst.un4_control_input_1_axb_13 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31_rep1 ;
    wire \current_shift_inst.un4_control_input1_11 ;
    wire \current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ;
    wire \current_shift_inst.un4_control_input1_14 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_9 ;
    wire \current_shift_inst.un4_control_input_1_axb_17 ;
    wire \current_shift_inst.un4_control_input1_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ;
    wire \current_shift_inst.un4_control_input_1_axb_22 ;
    wire \current_shift_inst.un4_control_input1_26 ;
    wire \current_shift_inst.un38_control_input_5_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_26 ;
    wire \current_shift_inst.un4_control_input_1_axb_6 ;
    wire \current_shift_inst.un4_control_input_1_axb_8 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_3 ;
    wire bfn_18_19_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.elapsed_time_ns_s1_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire \current_shift_inst.elapsed_time_ns_s1_11 ;
    wire bfn_18_20_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire \current_shift_inst.elapsed_time_ns_s1_19 ;
    wire bfn_18_21_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.elapsed_time_ns_s1_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire \current_shift_inst.elapsed_time_ns_s1_27 ;
    wire bfn_18_22_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire clk_100mhz_0;
    wire \current_shift_inst.timer_s1.N_166_i_g ;
    wire red_c_g;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire _gnd_net_;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__20615),
            .RESETB(N__18575),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clk_100mhz_0));
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__39010),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__39056),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({dangling_wire_16,N__21356,N__21349,N__21354,N__21348,N__21355,N__21347,N__21357,N__21344,N__21350,N__21343,N__21351,N__21345,N__21352,N__21346,N__21353}),
            .C({dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32}),
            .B({dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,N__39009,N__39059,dangling_wire_40,dangling_wire_41,dangling_wire_42,N__39057,N__39008,N__39058,N__39007}),
            .OHOLDTOP(),
            .O({dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,\pwm_generator_inst.un2_threshold_acc_2_1_16 ,\pwm_generator_inst.un2_threshold_acc_2_1_15 ,\pwm_generator_inst.un2_threshold_acc_2_14 ,\pwm_generator_inst.un2_threshold_acc_2_13 ,\pwm_generator_inst.un2_threshold_acc_2_12 ,\pwm_generator_inst.un2_threshold_acc_2_11 ,\pwm_generator_inst.un2_threshold_acc_2_10 ,\pwm_generator_inst.un2_threshold_acc_2_9 ,\pwm_generator_inst.un2_threshold_acc_2_8 ,\pwm_generator_inst.un2_threshold_acc_2_7 ,\pwm_generator_inst.un2_threshold_acc_2_6 ,\pwm_generator_inst.un2_threshold_acc_2_5 ,\pwm_generator_inst.un2_threshold_acc_2_4 ,\pwm_generator_inst.un2_threshold_acc_2_3 ,\pwm_generator_inst.un2_threshold_acc_2_2 ,\pwm_generator_inst.un2_threshold_acc_2_1 ,\pwm_generator_inst.un2_threshold_acc_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__38997),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__38990),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73}),
            .ADDSUBBOT(),
            .A({dangling_wire_74,N__21395,N__21440,N__21396,N__21441,N__21397,N__19998,N__20025,N__19917,N__19956,N__20286,N__18845,N__18825,N__18764,N__18782,N__18797}),
            .C({dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90}),
            .B({dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,N__38996,N__38993,dangling_wire_98,dangling_wire_99,dangling_wire_100,N__38991,N__38995,N__38992,N__38994}),
            .OHOLDTOP(),
            .O({dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,\pwm_generator_inst.un2_threshold_acc_1_25 ,\pwm_generator_inst.un2_threshold_acc_1_24 ,\pwm_generator_inst.un2_threshold_acc_1_23 ,\pwm_generator_inst.un2_threshold_acc_1_22 ,\pwm_generator_inst.un2_threshold_acc_1_21 ,\pwm_generator_inst.un2_threshold_acc_1_20 ,\pwm_generator_inst.un2_threshold_acc_1_19 ,\pwm_generator_inst.un2_threshold_acc_1_18 ,\pwm_generator_inst.un2_threshold_acc_1_17 ,\pwm_generator_inst.un2_threshold_acc_1_16 ,\pwm_generator_inst.un2_threshold_acc_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.un3_threshold_acc ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__48426),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__48428),
            .DIN(N__48427),
            .DOUT(N__48426),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__48428),
            .PADOUT(N__48427),
            .PADIN(N__48426),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T01_obuf_iopad (
            .OE(N__48417),
            .DIN(N__48416),
            .DOUT(N__48415),
            .PACKAGEPIN(T01));
    defparam T01_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T01_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T01_obuf_preio (
            .PADOEN(N__48417),
            .PADOUT(N__48416),
            .PADIN(N__48415),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__31658),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__48408),
            .DIN(N__48407),
            .DOUT(N__48406),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__48408),
            .PADOUT(N__48407),
            .PADIN(N__48406),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__48399),
            .DIN(N__48398),
            .DOUT(N__48397),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__48399),
            .PADOUT(N__48398),
            .PADIN(N__48397),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T23_obuf_iopad (
            .OE(N__48390),
            .DIN(N__48389),
            .DOUT(N__48388),
            .PACKAGEPIN(T23));
    defparam T23_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T23_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T23_obuf_preio (
            .PADOEN(N__48390),
            .PADOUT(N__48389),
            .PADIN(N__48388),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__32039),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__48381),
            .DIN(N__48380),
            .DOUT(N__48379),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__48381),
            .PADOUT(N__48380),
            .PADIN(N__48379),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20333),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__48372),
            .DIN(N__48371),
            .DOUT(N__48370),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__48372),
            .PADOUT(N__48371),
            .PADIN(N__48370),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__48363),
            .DIN(N__48362),
            .DOUT(N__48361),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__48363),
            .PADOUT(N__48362),
            .PADIN(N__48361),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__34076),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T12_obuf_iopad (
            .OE(N__48354),
            .DIN(N__48353),
            .DOUT(N__48352),
            .PACKAGEPIN(T12));
    defparam T12_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T12_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T12_obuf_preio (
            .PADOEN(N__48354),
            .PADOUT(N__48353),
            .PADIN(N__48352),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__32183),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__48345),
            .DIN(N__48344),
            .DOUT(N__48343),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__48345),
            .PADOUT(N__48344),
            .PADIN(N__48343),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__48336),
            .DIN(N__48335),
            .DOUT(N__48334),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__48336),
            .PADOUT(N__48335),
            .PADIN(N__48334),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__37613),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__48327),
            .DIN(N__48326),
            .DOUT(N__48325),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__48327),
            .PADOUT(N__48326),
            .PADIN(N__48325),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__27644),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__48318),
            .DIN(N__48317),
            .DOUT(N__48316),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__48318),
            .PADOUT(N__48317),
            .PADIN(N__48316),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__48309),
            .DIN(N__48308),
            .DOUT(N__48307),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__48309),
            .PADOUT(N__48308),
            .PADIN(N__48307),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__25190),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T45_obuf_iopad (
            .OE(N__48300),
            .DIN(N__48299),
            .DOUT(N__48298),
            .PACKAGEPIN(T45));
    defparam T45_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T45_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T45_obuf_preio (
            .PADOEN(N__48300),
            .PADOUT(N__48299),
            .PADIN(N__48298),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__32348),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_gb_io_iopad (
            .OE(N__48291),
            .DIN(N__48290),
            .DOUT(N__48289),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_gb_io_preio (
            .PADOEN(N__48291),
            .PADOUT(N__48290),
            .PADIN(N__48289),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_gb_io_iopad (
            .OE(N__48282),
            .DIN(N__48281),
            .DOUT(N__48280),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_gb_io_preio (
            .PADOEN(N__48282),
            .PADOUT(N__48281),
            .PADIN(N__48280),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__11474 (
            .O(N__48263),
            .I(N__48257));
    InMux I__11473 (
            .O(N__48262),
            .I(N__48257));
    LocalMux I__11472 (
            .O(N__48257),
            .I(N__48253));
    InMux I__11471 (
            .O(N__48256),
            .I(N__48250));
    Span4Mux_h I__11470 (
            .O(N__48253),
            .I(N__48247));
    LocalMux I__11469 (
            .O(N__48250),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    Odrv4 I__11468 (
            .O(N__48247),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__11467 (
            .O(N__48242),
            .I(N__48239));
    LocalMux I__11466 (
            .O(N__48239),
            .I(N__48234));
    InMux I__11465 (
            .O(N__48238),
            .I(N__48231));
    InMux I__11464 (
            .O(N__48237),
            .I(N__48228));
    Span4Mux_v I__11463 (
            .O(N__48234),
            .I(N__48225));
    LocalMux I__11462 (
            .O(N__48231),
            .I(N__48220));
    LocalMux I__11461 (
            .O(N__48228),
            .I(N__48220));
    Span4Mux_h I__11460 (
            .O(N__48225),
            .I(N__48214));
    Span4Mux_v I__11459 (
            .O(N__48220),
            .I(N__48214));
    InMux I__11458 (
            .O(N__48219),
            .I(N__48211));
    Odrv4 I__11457 (
            .O(N__48214),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    LocalMux I__11456 (
            .O(N__48211),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    InMux I__11455 (
            .O(N__48206),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__11454 (
            .O(N__48203),
            .I(N__48199));
    CascadeMux I__11453 (
            .O(N__48202),
            .I(N__48196));
    InMux I__11452 (
            .O(N__48199),
            .I(N__48193));
    InMux I__11451 (
            .O(N__48196),
            .I(N__48190));
    LocalMux I__11450 (
            .O(N__48193),
            .I(N__48186));
    LocalMux I__11449 (
            .O(N__48190),
            .I(N__48183));
    InMux I__11448 (
            .O(N__48189),
            .I(N__48180));
    Span4Mux_h I__11447 (
            .O(N__48186),
            .I(N__48177));
    Span4Mux_h I__11446 (
            .O(N__48183),
            .I(N__48174));
    LocalMux I__11445 (
            .O(N__48180),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv4 I__11444 (
            .O(N__48177),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv4 I__11443 (
            .O(N__48174),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    InMux I__11442 (
            .O(N__48167),
            .I(N__48163));
    CascadeMux I__11441 (
            .O(N__48166),
            .I(N__48160));
    LocalMux I__11440 (
            .O(N__48163),
            .I(N__48156));
    InMux I__11439 (
            .O(N__48160),
            .I(N__48153));
    CascadeMux I__11438 (
            .O(N__48159),
            .I(N__48150));
    Span4Mux_v I__11437 (
            .O(N__48156),
            .I(N__48147));
    LocalMux I__11436 (
            .O(N__48153),
            .I(N__48144));
    InMux I__11435 (
            .O(N__48150),
            .I(N__48141));
    Span4Mux_h I__11434 (
            .O(N__48147),
            .I(N__48133));
    Span4Mux_v I__11433 (
            .O(N__48144),
            .I(N__48133));
    LocalMux I__11432 (
            .O(N__48141),
            .I(N__48133));
    InMux I__11431 (
            .O(N__48140),
            .I(N__48130));
    Odrv4 I__11430 (
            .O(N__48133),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    LocalMux I__11429 (
            .O(N__48130),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    InMux I__11428 (
            .O(N__48125),
            .I(bfn_18_22_0_));
    CascadeMux I__11427 (
            .O(N__48122),
            .I(N__48118));
    CascadeMux I__11426 (
            .O(N__48121),
            .I(N__48115));
    InMux I__11425 (
            .O(N__48118),
            .I(N__48112));
    InMux I__11424 (
            .O(N__48115),
            .I(N__48109));
    LocalMux I__11423 (
            .O(N__48112),
            .I(N__48105));
    LocalMux I__11422 (
            .O(N__48109),
            .I(N__48102));
    InMux I__11421 (
            .O(N__48108),
            .I(N__48099));
    Span4Mux_h I__11420 (
            .O(N__48105),
            .I(N__48096));
    Span4Mux_h I__11419 (
            .O(N__48102),
            .I(N__48093));
    LocalMux I__11418 (
            .O(N__48099),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__11417 (
            .O(N__48096),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__11416 (
            .O(N__48093),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    InMux I__11415 (
            .O(N__48086),
            .I(N__48079));
    InMux I__11414 (
            .O(N__48085),
            .I(N__48079));
    InMux I__11413 (
            .O(N__48084),
            .I(N__48076));
    LocalMux I__11412 (
            .O(N__48079),
            .I(N__48073));
    LocalMux I__11411 (
            .O(N__48076),
            .I(N__48070));
    Span4Mux_v I__11410 (
            .O(N__48073),
            .I(N__48067));
    Span12Mux_v I__11409 (
            .O(N__48070),
            .I(N__48063));
    Span4Mux_v I__11408 (
            .O(N__48067),
            .I(N__48060));
    InMux I__11407 (
            .O(N__48066),
            .I(N__48057));
    Odrv12 I__11406 (
            .O(N__48063),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    Odrv4 I__11405 (
            .O(N__48060),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    LocalMux I__11404 (
            .O(N__48057),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    InMux I__11403 (
            .O(N__48050),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    InMux I__11402 (
            .O(N__48047),
            .I(N__48044));
    LocalMux I__11401 (
            .O(N__48044),
            .I(N__48040));
    InMux I__11400 (
            .O(N__48043),
            .I(N__48037));
    Span4Mux_h I__11399 (
            .O(N__48040),
            .I(N__48034));
    LocalMux I__11398 (
            .O(N__48037),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    Odrv4 I__11397 (
            .O(N__48034),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    CascadeMux I__11396 (
            .O(N__48029),
            .I(N__48026));
    InMux I__11395 (
            .O(N__48026),
            .I(N__48021));
    InMux I__11394 (
            .O(N__48025),
            .I(N__48018));
    InMux I__11393 (
            .O(N__48024),
            .I(N__48015));
    LocalMux I__11392 (
            .O(N__48021),
            .I(N__48010));
    LocalMux I__11391 (
            .O(N__48018),
            .I(N__48010));
    LocalMux I__11390 (
            .O(N__48015),
            .I(N__48005));
    Span4Mux_v I__11389 (
            .O(N__48010),
            .I(N__48005));
    Odrv4 I__11388 (
            .O(N__48005),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__11387 (
            .O(N__48002),
            .I(N__47998));
    InMux I__11386 (
            .O(N__48001),
            .I(N__47995));
    LocalMux I__11385 (
            .O(N__47998),
            .I(N__47992));
    LocalMux I__11384 (
            .O(N__47995),
            .I(N__47988));
    Span4Mux_v I__11383 (
            .O(N__47992),
            .I(N__47985));
    InMux I__11382 (
            .O(N__47991),
            .I(N__47982));
    Span12Mux_h I__11381 (
            .O(N__47988),
            .I(N__47978));
    Span4Mux_h I__11380 (
            .O(N__47985),
            .I(N__47973));
    LocalMux I__11379 (
            .O(N__47982),
            .I(N__47973));
    InMux I__11378 (
            .O(N__47981),
            .I(N__47970));
    Odrv12 I__11377 (
            .O(N__47978),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    Odrv4 I__11376 (
            .O(N__47973),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    LocalMux I__11375 (
            .O(N__47970),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    InMux I__11374 (
            .O(N__47963),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    InMux I__11373 (
            .O(N__47960),
            .I(N__47957));
    LocalMux I__11372 (
            .O(N__47957),
            .I(N__47953));
    InMux I__11371 (
            .O(N__47956),
            .I(N__47950));
    Span4Mux_h I__11370 (
            .O(N__47953),
            .I(N__47947));
    LocalMux I__11369 (
            .O(N__47950),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    Odrv4 I__11368 (
            .O(N__47947),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    CascadeMux I__11367 (
            .O(N__47942),
            .I(N__47939));
    InMux I__11366 (
            .O(N__47939),
            .I(N__47935));
    InMux I__11365 (
            .O(N__47938),
            .I(N__47932));
    LocalMux I__11364 (
            .O(N__47935),
            .I(N__47926));
    LocalMux I__11363 (
            .O(N__47932),
            .I(N__47926));
    InMux I__11362 (
            .O(N__47931),
            .I(N__47923));
    Span4Mux_v I__11361 (
            .O(N__47926),
            .I(N__47920));
    LocalMux I__11360 (
            .O(N__47923),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    Odrv4 I__11359 (
            .O(N__47920),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    InMux I__11358 (
            .O(N__47915),
            .I(N__47911));
    InMux I__11357 (
            .O(N__47914),
            .I(N__47908));
    LocalMux I__11356 (
            .O(N__47911),
            .I(N__47904));
    LocalMux I__11355 (
            .O(N__47908),
            .I(N__47901));
    InMux I__11354 (
            .O(N__47907),
            .I(N__47898));
    Span4Mux_v I__11353 (
            .O(N__47904),
            .I(N__47894));
    Span4Mux_v I__11352 (
            .O(N__47901),
            .I(N__47889));
    LocalMux I__11351 (
            .O(N__47898),
            .I(N__47889));
    InMux I__11350 (
            .O(N__47897),
            .I(N__47886));
    Odrv4 I__11349 (
            .O(N__47894),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    Odrv4 I__11348 (
            .O(N__47889),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    LocalMux I__11347 (
            .O(N__47886),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    InMux I__11346 (
            .O(N__47879),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    ClkMux I__11345 (
            .O(N__47876),
            .I(N__47519));
    ClkMux I__11344 (
            .O(N__47875),
            .I(N__47519));
    ClkMux I__11343 (
            .O(N__47874),
            .I(N__47519));
    ClkMux I__11342 (
            .O(N__47873),
            .I(N__47519));
    ClkMux I__11341 (
            .O(N__47872),
            .I(N__47519));
    ClkMux I__11340 (
            .O(N__47871),
            .I(N__47519));
    ClkMux I__11339 (
            .O(N__47870),
            .I(N__47519));
    ClkMux I__11338 (
            .O(N__47869),
            .I(N__47519));
    ClkMux I__11337 (
            .O(N__47868),
            .I(N__47519));
    ClkMux I__11336 (
            .O(N__47867),
            .I(N__47519));
    ClkMux I__11335 (
            .O(N__47866),
            .I(N__47519));
    ClkMux I__11334 (
            .O(N__47865),
            .I(N__47519));
    ClkMux I__11333 (
            .O(N__47864),
            .I(N__47519));
    ClkMux I__11332 (
            .O(N__47863),
            .I(N__47519));
    ClkMux I__11331 (
            .O(N__47862),
            .I(N__47519));
    ClkMux I__11330 (
            .O(N__47861),
            .I(N__47519));
    ClkMux I__11329 (
            .O(N__47860),
            .I(N__47519));
    ClkMux I__11328 (
            .O(N__47859),
            .I(N__47519));
    ClkMux I__11327 (
            .O(N__47858),
            .I(N__47519));
    ClkMux I__11326 (
            .O(N__47857),
            .I(N__47519));
    ClkMux I__11325 (
            .O(N__47856),
            .I(N__47519));
    ClkMux I__11324 (
            .O(N__47855),
            .I(N__47519));
    ClkMux I__11323 (
            .O(N__47854),
            .I(N__47519));
    ClkMux I__11322 (
            .O(N__47853),
            .I(N__47519));
    ClkMux I__11321 (
            .O(N__47852),
            .I(N__47519));
    ClkMux I__11320 (
            .O(N__47851),
            .I(N__47519));
    ClkMux I__11319 (
            .O(N__47850),
            .I(N__47519));
    ClkMux I__11318 (
            .O(N__47849),
            .I(N__47519));
    ClkMux I__11317 (
            .O(N__47848),
            .I(N__47519));
    ClkMux I__11316 (
            .O(N__47847),
            .I(N__47519));
    ClkMux I__11315 (
            .O(N__47846),
            .I(N__47519));
    ClkMux I__11314 (
            .O(N__47845),
            .I(N__47519));
    ClkMux I__11313 (
            .O(N__47844),
            .I(N__47519));
    ClkMux I__11312 (
            .O(N__47843),
            .I(N__47519));
    ClkMux I__11311 (
            .O(N__47842),
            .I(N__47519));
    ClkMux I__11310 (
            .O(N__47841),
            .I(N__47519));
    ClkMux I__11309 (
            .O(N__47840),
            .I(N__47519));
    ClkMux I__11308 (
            .O(N__47839),
            .I(N__47519));
    ClkMux I__11307 (
            .O(N__47838),
            .I(N__47519));
    ClkMux I__11306 (
            .O(N__47837),
            .I(N__47519));
    ClkMux I__11305 (
            .O(N__47836),
            .I(N__47519));
    ClkMux I__11304 (
            .O(N__47835),
            .I(N__47519));
    ClkMux I__11303 (
            .O(N__47834),
            .I(N__47519));
    ClkMux I__11302 (
            .O(N__47833),
            .I(N__47519));
    ClkMux I__11301 (
            .O(N__47832),
            .I(N__47519));
    ClkMux I__11300 (
            .O(N__47831),
            .I(N__47519));
    ClkMux I__11299 (
            .O(N__47830),
            .I(N__47519));
    ClkMux I__11298 (
            .O(N__47829),
            .I(N__47519));
    ClkMux I__11297 (
            .O(N__47828),
            .I(N__47519));
    ClkMux I__11296 (
            .O(N__47827),
            .I(N__47519));
    ClkMux I__11295 (
            .O(N__47826),
            .I(N__47519));
    ClkMux I__11294 (
            .O(N__47825),
            .I(N__47519));
    ClkMux I__11293 (
            .O(N__47824),
            .I(N__47519));
    ClkMux I__11292 (
            .O(N__47823),
            .I(N__47519));
    ClkMux I__11291 (
            .O(N__47822),
            .I(N__47519));
    ClkMux I__11290 (
            .O(N__47821),
            .I(N__47519));
    ClkMux I__11289 (
            .O(N__47820),
            .I(N__47519));
    ClkMux I__11288 (
            .O(N__47819),
            .I(N__47519));
    ClkMux I__11287 (
            .O(N__47818),
            .I(N__47519));
    ClkMux I__11286 (
            .O(N__47817),
            .I(N__47519));
    ClkMux I__11285 (
            .O(N__47816),
            .I(N__47519));
    ClkMux I__11284 (
            .O(N__47815),
            .I(N__47519));
    ClkMux I__11283 (
            .O(N__47814),
            .I(N__47519));
    ClkMux I__11282 (
            .O(N__47813),
            .I(N__47519));
    ClkMux I__11281 (
            .O(N__47812),
            .I(N__47519));
    ClkMux I__11280 (
            .O(N__47811),
            .I(N__47519));
    ClkMux I__11279 (
            .O(N__47810),
            .I(N__47519));
    ClkMux I__11278 (
            .O(N__47809),
            .I(N__47519));
    ClkMux I__11277 (
            .O(N__47808),
            .I(N__47519));
    ClkMux I__11276 (
            .O(N__47807),
            .I(N__47519));
    ClkMux I__11275 (
            .O(N__47806),
            .I(N__47519));
    ClkMux I__11274 (
            .O(N__47805),
            .I(N__47519));
    ClkMux I__11273 (
            .O(N__47804),
            .I(N__47519));
    ClkMux I__11272 (
            .O(N__47803),
            .I(N__47519));
    ClkMux I__11271 (
            .O(N__47802),
            .I(N__47519));
    ClkMux I__11270 (
            .O(N__47801),
            .I(N__47519));
    ClkMux I__11269 (
            .O(N__47800),
            .I(N__47519));
    ClkMux I__11268 (
            .O(N__47799),
            .I(N__47519));
    ClkMux I__11267 (
            .O(N__47798),
            .I(N__47519));
    ClkMux I__11266 (
            .O(N__47797),
            .I(N__47519));
    ClkMux I__11265 (
            .O(N__47796),
            .I(N__47519));
    ClkMux I__11264 (
            .O(N__47795),
            .I(N__47519));
    ClkMux I__11263 (
            .O(N__47794),
            .I(N__47519));
    ClkMux I__11262 (
            .O(N__47793),
            .I(N__47519));
    ClkMux I__11261 (
            .O(N__47792),
            .I(N__47519));
    ClkMux I__11260 (
            .O(N__47791),
            .I(N__47519));
    ClkMux I__11259 (
            .O(N__47790),
            .I(N__47519));
    ClkMux I__11258 (
            .O(N__47789),
            .I(N__47519));
    ClkMux I__11257 (
            .O(N__47788),
            .I(N__47519));
    ClkMux I__11256 (
            .O(N__47787),
            .I(N__47519));
    ClkMux I__11255 (
            .O(N__47786),
            .I(N__47519));
    ClkMux I__11254 (
            .O(N__47785),
            .I(N__47519));
    ClkMux I__11253 (
            .O(N__47784),
            .I(N__47519));
    ClkMux I__11252 (
            .O(N__47783),
            .I(N__47519));
    ClkMux I__11251 (
            .O(N__47782),
            .I(N__47519));
    ClkMux I__11250 (
            .O(N__47781),
            .I(N__47519));
    ClkMux I__11249 (
            .O(N__47780),
            .I(N__47519));
    ClkMux I__11248 (
            .O(N__47779),
            .I(N__47519));
    ClkMux I__11247 (
            .O(N__47778),
            .I(N__47519));
    ClkMux I__11246 (
            .O(N__47777),
            .I(N__47519));
    ClkMux I__11245 (
            .O(N__47776),
            .I(N__47519));
    ClkMux I__11244 (
            .O(N__47775),
            .I(N__47519));
    ClkMux I__11243 (
            .O(N__47774),
            .I(N__47519));
    ClkMux I__11242 (
            .O(N__47773),
            .I(N__47519));
    ClkMux I__11241 (
            .O(N__47772),
            .I(N__47519));
    ClkMux I__11240 (
            .O(N__47771),
            .I(N__47519));
    ClkMux I__11239 (
            .O(N__47770),
            .I(N__47519));
    ClkMux I__11238 (
            .O(N__47769),
            .I(N__47519));
    ClkMux I__11237 (
            .O(N__47768),
            .I(N__47519));
    ClkMux I__11236 (
            .O(N__47767),
            .I(N__47519));
    ClkMux I__11235 (
            .O(N__47766),
            .I(N__47519));
    ClkMux I__11234 (
            .O(N__47765),
            .I(N__47519));
    ClkMux I__11233 (
            .O(N__47764),
            .I(N__47519));
    ClkMux I__11232 (
            .O(N__47763),
            .I(N__47519));
    ClkMux I__11231 (
            .O(N__47762),
            .I(N__47519));
    ClkMux I__11230 (
            .O(N__47761),
            .I(N__47519));
    ClkMux I__11229 (
            .O(N__47760),
            .I(N__47519));
    ClkMux I__11228 (
            .O(N__47759),
            .I(N__47519));
    ClkMux I__11227 (
            .O(N__47758),
            .I(N__47519));
    GlobalMux I__11226 (
            .O(N__47519),
            .I(clk_100mhz_0));
    CEMux I__11225 (
            .O(N__47516),
            .I(N__47489));
    CEMux I__11224 (
            .O(N__47515),
            .I(N__47489));
    CEMux I__11223 (
            .O(N__47514),
            .I(N__47489));
    CEMux I__11222 (
            .O(N__47513),
            .I(N__47489));
    CEMux I__11221 (
            .O(N__47512),
            .I(N__47489));
    CEMux I__11220 (
            .O(N__47511),
            .I(N__47489));
    CEMux I__11219 (
            .O(N__47510),
            .I(N__47489));
    CEMux I__11218 (
            .O(N__47509),
            .I(N__47489));
    CEMux I__11217 (
            .O(N__47508),
            .I(N__47489));
    GlobalMux I__11216 (
            .O(N__47489),
            .I(N__47486));
    gio2CtrlBuf I__11215 (
            .O(N__47486),
            .I(\current_shift_inst.timer_s1.N_166_i_g ));
    InMux I__11214 (
            .O(N__47483),
            .I(N__47466));
    InMux I__11213 (
            .O(N__47482),
            .I(N__47463));
    InMux I__11212 (
            .O(N__47481),
            .I(N__47460));
    InMux I__11211 (
            .O(N__47480),
            .I(N__47457));
    InMux I__11210 (
            .O(N__47479),
            .I(N__47454));
    InMux I__11209 (
            .O(N__47478),
            .I(N__47449));
    InMux I__11208 (
            .O(N__47477),
            .I(N__47449));
    InMux I__11207 (
            .O(N__47476),
            .I(N__47444));
    InMux I__11206 (
            .O(N__47475),
            .I(N__47444));
    InMux I__11205 (
            .O(N__47474),
            .I(N__47439));
    InMux I__11204 (
            .O(N__47473),
            .I(N__47439));
    InMux I__11203 (
            .O(N__47472),
            .I(N__47434));
    InMux I__11202 (
            .O(N__47471),
            .I(N__47434));
    InMux I__11201 (
            .O(N__47470),
            .I(N__47431));
    InMux I__11200 (
            .O(N__47469),
            .I(N__47428));
    LocalMux I__11199 (
            .O(N__47466),
            .I(N__47425));
    LocalMux I__11198 (
            .O(N__47463),
            .I(N__47422));
    LocalMux I__11197 (
            .O(N__47460),
            .I(N__47419));
    LocalMux I__11196 (
            .O(N__47457),
            .I(N__47411));
    LocalMux I__11195 (
            .O(N__47454),
            .I(N__47355));
    LocalMux I__11194 (
            .O(N__47449),
            .I(N__47346));
    LocalMux I__11193 (
            .O(N__47444),
            .I(N__47343));
    LocalMux I__11192 (
            .O(N__47439),
            .I(N__47336));
    LocalMux I__11191 (
            .O(N__47434),
            .I(N__47308));
    LocalMux I__11190 (
            .O(N__47431),
            .I(N__47296));
    LocalMux I__11189 (
            .O(N__47428),
            .I(N__47290));
    Glb2LocalMux I__11188 (
            .O(N__47425),
            .I(N__47030));
    Glb2LocalMux I__11187 (
            .O(N__47422),
            .I(N__47030));
    Glb2LocalMux I__11186 (
            .O(N__47419),
            .I(N__47030));
    SRMux I__11185 (
            .O(N__47418),
            .I(N__47030));
    SRMux I__11184 (
            .O(N__47417),
            .I(N__47030));
    SRMux I__11183 (
            .O(N__47416),
            .I(N__47030));
    SRMux I__11182 (
            .O(N__47415),
            .I(N__47030));
    SRMux I__11181 (
            .O(N__47414),
            .I(N__47030));
    Glb2LocalMux I__11180 (
            .O(N__47411),
            .I(N__47030));
    SRMux I__11179 (
            .O(N__47410),
            .I(N__47030));
    SRMux I__11178 (
            .O(N__47409),
            .I(N__47030));
    SRMux I__11177 (
            .O(N__47408),
            .I(N__47030));
    SRMux I__11176 (
            .O(N__47407),
            .I(N__47030));
    SRMux I__11175 (
            .O(N__47406),
            .I(N__47030));
    SRMux I__11174 (
            .O(N__47405),
            .I(N__47030));
    SRMux I__11173 (
            .O(N__47404),
            .I(N__47030));
    SRMux I__11172 (
            .O(N__47403),
            .I(N__47030));
    SRMux I__11171 (
            .O(N__47402),
            .I(N__47030));
    SRMux I__11170 (
            .O(N__47401),
            .I(N__47030));
    SRMux I__11169 (
            .O(N__47400),
            .I(N__47030));
    SRMux I__11168 (
            .O(N__47399),
            .I(N__47030));
    SRMux I__11167 (
            .O(N__47398),
            .I(N__47030));
    SRMux I__11166 (
            .O(N__47397),
            .I(N__47030));
    SRMux I__11165 (
            .O(N__47396),
            .I(N__47030));
    SRMux I__11164 (
            .O(N__47395),
            .I(N__47030));
    SRMux I__11163 (
            .O(N__47394),
            .I(N__47030));
    SRMux I__11162 (
            .O(N__47393),
            .I(N__47030));
    SRMux I__11161 (
            .O(N__47392),
            .I(N__47030));
    SRMux I__11160 (
            .O(N__47391),
            .I(N__47030));
    SRMux I__11159 (
            .O(N__47390),
            .I(N__47030));
    SRMux I__11158 (
            .O(N__47389),
            .I(N__47030));
    SRMux I__11157 (
            .O(N__47388),
            .I(N__47030));
    SRMux I__11156 (
            .O(N__47387),
            .I(N__47030));
    SRMux I__11155 (
            .O(N__47386),
            .I(N__47030));
    SRMux I__11154 (
            .O(N__47385),
            .I(N__47030));
    SRMux I__11153 (
            .O(N__47384),
            .I(N__47030));
    SRMux I__11152 (
            .O(N__47383),
            .I(N__47030));
    SRMux I__11151 (
            .O(N__47382),
            .I(N__47030));
    SRMux I__11150 (
            .O(N__47381),
            .I(N__47030));
    SRMux I__11149 (
            .O(N__47380),
            .I(N__47030));
    SRMux I__11148 (
            .O(N__47379),
            .I(N__47030));
    SRMux I__11147 (
            .O(N__47378),
            .I(N__47030));
    SRMux I__11146 (
            .O(N__47377),
            .I(N__47030));
    SRMux I__11145 (
            .O(N__47376),
            .I(N__47030));
    SRMux I__11144 (
            .O(N__47375),
            .I(N__47030));
    SRMux I__11143 (
            .O(N__47374),
            .I(N__47030));
    SRMux I__11142 (
            .O(N__47373),
            .I(N__47030));
    SRMux I__11141 (
            .O(N__47372),
            .I(N__47030));
    SRMux I__11140 (
            .O(N__47371),
            .I(N__47030));
    SRMux I__11139 (
            .O(N__47370),
            .I(N__47030));
    SRMux I__11138 (
            .O(N__47369),
            .I(N__47030));
    SRMux I__11137 (
            .O(N__47368),
            .I(N__47030));
    SRMux I__11136 (
            .O(N__47367),
            .I(N__47030));
    SRMux I__11135 (
            .O(N__47366),
            .I(N__47030));
    SRMux I__11134 (
            .O(N__47365),
            .I(N__47030));
    SRMux I__11133 (
            .O(N__47364),
            .I(N__47030));
    SRMux I__11132 (
            .O(N__47363),
            .I(N__47030));
    SRMux I__11131 (
            .O(N__47362),
            .I(N__47030));
    SRMux I__11130 (
            .O(N__47361),
            .I(N__47030));
    SRMux I__11129 (
            .O(N__47360),
            .I(N__47030));
    SRMux I__11128 (
            .O(N__47359),
            .I(N__47030));
    SRMux I__11127 (
            .O(N__47358),
            .I(N__47030));
    Glb2LocalMux I__11126 (
            .O(N__47355),
            .I(N__47030));
    SRMux I__11125 (
            .O(N__47354),
            .I(N__47030));
    SRMux I__11124 (
            .O(N__47353),
            .I(N__47030));
    SRMux I__11123 (
            .O(N__47352),
            .I(N__47030));
    SRMux I__11122 (
            .O(N__47351),
            .I(N__47030));
    SRMux I__11121 (
            .O(N__47350),
            .I(N__47030));
    SRMux I__11120 (
            .O(N__47349),
            .I(N__47030));
    Glb2LocalMux I__11119 (
            .O(N__47346),
            .I(N__47030));
    Glb2LocalMux I__11118 (
            .O(N__47343),
            .I(N__47030));
    SRMux I__11117 (
            .O(N__47342),
            .I(N__47030));
    SRMux I__11116 (
            .O(N__47341),
            .I(N__47030));
    SRMux I__11115 (
            .O(N__47340),
            .I(N__47030));
    SRMux I__11114 (
            .O(N__47339),
            .I(N__47030));
    Glb2LocalMux I__11113 (
            .O(N__47336),
            .I(N__47030));
    SRMux I__11112 (
            .O(N__47335),
            .I(N__47030));
    SRMux I__11111 (
            .O(N__47334),
            .I(N__47030));
    SRMux I__11110 (
            .O(N__47333),
            .I(N__47030));
    SRMux I__11109 (
            .O(N__47332),
            .I(N__47030));
    SRMux I__11108 (
            .O(N__47331),
            .I(N__47030));
    SRMux I__11107 (
            .O(N__47330),
            .I(N__47030));
    SRMux I__11106 (
            .O(N__47329),
            .I(N__47030));
    SRMux I__11105 (
            .O(N__47328),
            .I(N__47030));
    SRMux I__11104 (
            .O(N__47327),
            .I(N__47030));
    SRMux I__11103 (
            .O(N__47326),
            .I(N__47030));
    SRMux I__11102 (
            .O(N__47325),
            .I(N__47030));
    SRMux I__11101 (
            .O(N__47324),
            .I(N__47030));
    SRMux I__11100 (
            .O(N__47323),
            .I(N__47030));
    SRMux I__11099 (
            .O(N__47322),
            .I(N__47030));
    SRMux I__11098 (
            .O(N__47321),
            .I(N__47030));
    SRMux I__11097 (
            .O(N__47320),
            .I(N__47030));
    SRMux I__11096 (
            .O(N__47319),
            .I(N__47030));
    SRMux I__11095 (
            .O(N__47318),
            .I(N__47030));
    SRMux I__11094 (
            .O(N__47317),
            .I(N__47030));
    SRMux I__11093 (
            .O(N__47316),
            .I(N__47030));
    SRMux I__11092 (
            .O(N__47315),
            .I(N__47030));
    SRMux I__11091 (
            .O(N__47314),
            .I(N__47030));
    SRMux I__11090 (
            .O(N__47313),
            .I(N__47030));
    SRMux I__11089 (
            .O(N__47312),
            .I(N__47030));
    SRMux I__11088 (
            .O(N__47311),
            .I(N__47030));
    Glb2LocalMux I__11087 (
            .O(N__47308),
            .I(N__47030));
    SRMux I__11086 (
            .O(N__47307),
            .I(N__47030));
    SRMux I__11085 (
            .O(N__47306),
            .I(N__47030));
    SRMux I__11084 (
            .O(N__47305),
            .I(N__47030));
    SRMux I__11083 (
            .O(N__47304),
            .I(N__47030));
    SRMux I__11082 (
            .O(N__47303),
            .I(N__47030));
    SRMux I__11081 (
            .O(N__47302),
            .I(N__47030));
    SRMux I__11080 (
            .O(N__47301),
            .I(N__47030));
    SRMux I__11079 (
            .O(N__47300),
            .I(N__47030));
    SRMux I__11078 (
            .O(N__47299),
            .I(N__47030));
    Glb2LocalMux I__11077 (
            .O(N__47296),
            .I(N__47030));
    SRMux I__11076 (
            .O(N__47295),
            .I(N__47030));
    SRMux I__11075 (
            .O(N__47294),
            .I(N__47030));
    SRMux I__11074 (
            .O(N__47293),
            .I(N__47030));
    Glb2LocalMux I__11073 (
            .O(N__47290),
            .I(N__47030));
    SRMux I__11072 (
            .O(N__47289),
            .I(N__47030));
    SRMux I__11071 (
            .O(N__47288),
            .I(N__47030));
    SRMux I__11070 (
            .O(N__47287),
            .I(N__47030));
    SRMux I__11069 (
            .O(N__47286),
            .I(N__47030));
    SRMux I__11068 (
            .O(N__47285),
            .I(N__47030));
    SRMux I__11067 (
            .O(N__47284),
            .I(N__47030));
    SRMux I__11066 (
            .O(N__47283),
            .I(N__47030));
    SRMux I__11065 (
            .O(N__47282),
            .I(N__47030));
    SRMux I__11064 (
            .O(N__47281),
            .I(N__47030));
    GlobalMux I__11063 (
            .O(N__47030),
            .I(N__47027));
    gio2CtrlBuf I__11062 (
            .O(N__47027),
            .I(red_c_g));
    InMux I__11061 (
            .O(N__47024),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    InMux I__11060 (
            .O(N__47021),
            .I(N__47016));
    InMux I__11059 (
            .O(N__47020),
            .I(N__47013));
    InMux I__11058 (
            .O(N__47019),
            .I(N__47010));
    LocalMux I__11057 (
            .O(N__47016),
            .I(N__47007));
    LocalMux I__11056 (
            .O(N__47013),
            .I(N__47004));
    LocalMux I__11055 (
            .O(N__47010),
            .I(N__47001));
    Span4Mux_v I__11054 (
            .O(N__47007),
            .I(N__46998));
    Span4Mux_h I__11053 (
            .O(N__47004),
            .I(N__46995));
    Sp12to4 I__11052 (
            .O(N__47001),
            .I(N__46992));
    Span4Mux_h I__11051 (
            .O(N__46998),
            .I(N__46987));
    Span4Mux_h I__11050 (
            .O(N__46995),
            .I(N__46987));
    Odrv12 I__11049 (
            .O(N__46992),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    Odrv4 I__11048 (
            .O(N__46987),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    CascadeMux I__11047 (
            .O(N__46982),
            .I(N__46978));
    CascadeMux I__11046 (
            .O(N__46981),
            .I(N__46975));
    InMux I__11045 (
            .O(N__46978),
            .I(N__46972));
    InMux I__11044 (
            .O(N__46975),
            .I(N__46969));
    LocalMux I__11043 (
            .O(N__46972),
            .I(N__46965));
    LocalMux I__11042 (
            .O(N__46969),
            .I(N__46962));
    InMux I__11041 (
            .O(N__46968),
            .I(N__46959));
    Span4Mux_h I__11040 (
            .O(N__46965),
            .I(N__46956));
    Span4Mux_h I__11039 (
            .O(N__46962),
            .I(N__46953));
    LocalMux I__11038 (
            .O(N__46959),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv4 I__11037 (
            .O(N__46956),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv4 I__11036 (
            .O(N__46953),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    InMux I__11035 (
            .O(N__46946),
            .I(N__46942));
    InMux I__11034 (
            .O(N__46945),
            .I(N__46939));
    LocalMux I__11033 (
            .O(N__46942),
            .I(N__46936));
    LocalMux I__11032 (
            .O(N__46939),
            .I(N__46930));
    Span4Mux_h I__11031 (
            .O(N__46936),
            .I(N__46930));
    InMux I__11030 (
            .O(N__46935),
            .I(N__46926));
    Span4Mux_h I__11029 (
            .O(N__46930),
            .I(N__46923));
    InMux I__11028 (
            .O(N__46929),
            .I(N__46920));
    LocalMux I__11027 (
            .O(N__46926),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    Odrv4 I__11026 (
            .O(N__46923),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    LocalMux I__11025 (
            .O(N__46920),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    InMux I__11024 (
            .O(N__46913),
            .I(bfn_18_21_0_));
    CascadeMux I__11023 (
            .O(N__46910),
            .I(N__46906));
    CascadeMux I__11022 (
            .O(N__46909),
            .I(N__46903));
    InMux I__11021 (
            .O(N__46906),
            .I(N__46900));
    InMux I__11020 (
            .O(N__46903),
            .I(N__46897));
    LocalMux I__11019 (
            .O(N__46900),
            .I(N__46893));
    LocalMux I__11018 (
            .O(N__46897),
            .I(N__46890));
    InMux I__11017 (
            .O(N__46896),
            .I(N__46887));
    Span4Mux_h I__11016 (
            .O(N__46893),
            .I(N__46884));
    Span4Mux_h I__11015 (
            .O(N__46890),
            .I(N__46881));
    LocalMux I__11014 (
            .O(N__46887),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__11013 (
            .O(N__46884),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__11012 (
            .O(N__46881),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    InMux I__11011 (
            .O(N__46874),
            .I(N__46869));
    InMux I__11010 (
            .O(N__46873),
            .I(N__46864));
    InMux I__11009 (
            .O(N__46872),
            .I(N__46864));
    LocalMux I__11008 (
            .O(N__46869),
            .I(N__46859));
    LocalMux I__11007 (
            .O(N__46864),
            .I(N__46859));
    Span12Mux_v I__11006 (
            .O(N__46859),
            .I(N__46855));
    InMux I__11005 (
            .O(N__46858),
            .I(N__46852));
    Odrv12 I__11004 (
            .O(N__46855),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    LocalMux I__11003 (
            .O(N__46852),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    InMux I__11002 (
            .O(N__46847),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__11001 (
            .O(N__46844),
            .I(N__46841));
    InMux I__11000 (
            .O(N__46841),
            .I(N__46836));
    InMux I__10999 (
            .O(N__46840),
            .I(N__46833));
    InMux I__10998 (
            .O(N__46839),
            .I(N__46830));
    LocalMux I__10997 (
            .O(N__46836),
            .I(N__46825));
    LocalMux I__10996 (
            .O(N__46833),
            .I(N__46825));
    LocalMux I__10995 (
            .O(N__46830),
            .I(N__46820));
    Span4Mux_v I__10994 (
            .O(N__46825),
            .I(N__46820));
    Odrv4 I__10993 (
            .O(N__46820),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    InMux I__10992 (
            .O(N__46817),
            .I(N__46814));
    LocalMux I__10991 (
            .O(N__46814),
            .I(N__46809));
    InMux I__10990 (
            .O(N__46813),
            .I(N__46806));
    InMux I__10989 (
            .O(N__46812),
            .I(N__46802));
    Span4Mux_v I__10988 (
            .O(N__46809),
            .I(N__46797));
    LocalMux I__10987 (
            .O(N__46806),
            .I(N__46797));
    InMux I__10986 (
            .O(N__46805),
            .I(N__46794));
    LocalMux I__10985 (
            .O(N__46802),
            .I(N__46791));
    Span4Mux_v I__10984 (
            .O(N__46797),
            .I(N__46788));
    LocalMux I__10983 (
            .O(N__46794),
            .I(N__46785));
    Span4Mux_v I__10982 (
            .O(N__46791),
            .I(N__46782));
    Odrv4 I__10981 (
            .O(N__46788),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    Odrv4 I__10980 (
            .O(N__46785),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    Odrv4 I__10979 (
            .O(N__46782),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    InMux I__10978 (
            .O(N__46775),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    InMux I__10977 (
            .O(N__46772),
            .I(N__46766));
    InMux I__10976 (
            .O(N__46771),
            .I(N__46766));
    LocalMux I__10975 (
            .O(N__46766),
            .I(N__46762));
    InMux I__10974 (
            .O(N__46765),
            .I(N__46759));
    Span4Mux_v I__10973 (
            .O(N__46762),
            .I(N__46756));
    LocalMux I__10972 (
            .O(N__46759),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    Odrv4 I__10971 (
            .O(N__46756),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    InMux I__10970 (
            .O(N__46751),
            .I(N__46742));
    InMux I__10969 (
            .O(N__46750),
            .I(N__46742));
    InMux I__10968 (
            .O(N__46749),
            .I(N__46742));
    LocalMux I__10967 (
            .O(N__46742),
            .I(N__46739));
    Span4Mux_v I__10966 (
            .O(N__46739),
            .I(N__46736));
    Span4Mux_h I__10965 (
            .O(N__46736),
            .I(N__46732));
    InMux I__10964 (
            .O(N__46735),
            .I(N__46729));
    Odrv4 I__10963 (
            .O(N__46732),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    LocalMux I__10962 (
            .O(N__46729),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    InMux I__10961 (
            .O(N__46724),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__10960 (
            .O(N__46721),
            .I(N__46718));
    InMux I__10959 (
            .O(N__46718),
            .I(N__46714));
    InMux I__10958 (
            .O(N__46717),
            .I(N__46711));
    LocalMux I__10957 (
            .O(N__46714),
            .I(N__46705));
    LocalMux I__10956 (
            .O(N__46711),
            .I(N__46705));
    InMux I__10955 (
            .O(N__46710),
            .I(N__46702));
    Span4Mux_h I__10954 (
            .O(N__46705),
            .I(N__46699));
    LocalMux I__10953 (
            .O(N__46702),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    Odrv4 I__10952 (
            .O(N__46699),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    InMux I__10951 (
            .O(N__46694),
            .I(N__46689));
    InMux I__10950 (
            .O(N__46693),
            .I(N__46686));
    InMux I__10949 (
            .O(N__46692),
            .I(N__46683));
    LocalMux I__10948 (
            .O(N__46689),
            .I(N__46677));
    LocalMux I__10947 (
            .O(N__46686),
            .I(N__46677));
    LocalMux I__10946 (
            .O(N__46683),
            .I(N__46674));
    InMux I__10945 (
            .O(N__46682),
            .I(N__46671));
    Span4Mux_h I__10944 (
            .O(N__46677),
            .I(N__46668));
    Span4Mux_h I__10943 (
            .O(N__46674),
            .I(N__46663));
    LocalMux I__10942 (
            .O(N__46671),
            .I(N__46663));
    Odrv4 I__10941 (
            .O(N__46668),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    Odrv4 I__10940 (
            .O(N__46663),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    InMux I__10939 (
            .O(N__46658),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__10938 (
            .O(N__46655),
            .I(N__46651));
    CascadeMux I__10937 (
            .O(N__46654),
            .I(N__46648));
    InMux I__10936 (
            .O(N__46651),
            .I(N__46643));
    InMux I__10935 (
            .O(N__46648),
            .I(N__46643));
    LocalMux I__10934 (
            .O(N__46643),
            .I(N__46639));
    InMux I__10933 (
            .O(N__46642),
            .I(N__46636));
    Span4Mux_h I__10932 (
            .O(N__46639),
            .I(N__46633));
    LocalMux I__10931 (
            .O(N__46636),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    Odrv4 I__10930 (
            .O(N__46633),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    CascadeMux I__10929 (
            .O(N__46628),
            .I(N__46624));
    CascadeMux I__10928 (
            .O(N__46627),
            .I(N__46621));
    InMux I__10927 (
            .O(N__46624),
            .I(N__46617));
    InMux I__10926 (
            .O(N__46621),
            .I(N__46612));
    InMux I__10925 (
            .O(N__46620),
            .I(N__46612));
    LocalMux I__10924 (
            .O(N__46617),
            .I(N__46609));
    LocalMux I__10923 (
            .O(N__46612),
            .I(N__46606));
    Span4Mux_h I__10922 (
            .O(N__46609),
            .I(N__46602));
    Span4Mux_h I__10921 (
            .O(N__46606),
            .I(N__46599));
    InMux I__10920 (
            .O(N__46605),
            .I(N__46596));
    Odrv4 I__10919 (
            .O(N__46602),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv4 I__10918 (
            .O(N__46599),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    LocalMux I__10917 (
            .O(N__46596),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    InMux I__10916 (
            .O(N__46589),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    InMux I__10915 (
            .O(N__46586),
            .I(N__46580));
    InMux I__10914 (
            .O(N__46585),
            .I(N__46580));
    LocalMux I__10913 (
            .O(N__46580),
            .I(N__46576));
    InMux I__10912 (
            .O(N__46579),
            .I(N__46573));
    Span4Mux_h I__10911 (
            .O(N__46576),
            .I(N__46570));
    LocalMux I__10910 (
            .O(N__46573),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    Odrv4 I__10909 (
            .O(N__46570),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    CascadeMux I__10908 (
            .O(N__46565),
            .I(N__46562));
    InMux I__10907 (
            .O(N__46562),
            .I(N__46559));
    LocalMux I__10906 (
            .O(N__46559),
            .I(N__46554));
    InMux I__10905 (
            .O(N__46558),
            .I(N__46551));
    InMux I__10904 (
            .O(N__46557),
            .I(N__46548));
    Span4Mux_v I__10903 (
            .O(N__46554),
            .I(N__46543));
    LocalMux I__10902 (
            .O(N__46551),
            .I(N__46543));
    LocalMux I__10901 (
            .O(N__46548),
            .I(N__46539));
    Span4Mux_h I__10900 (
            .O(N__46543),
            .I(N__46536));
    InMux I__10899 (
            .O(N__46542),
            .I(N__46533));
    Odrv12 I__10898 (
            .O(N__46539),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv4 I__10897 (
            .O(N__46536),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    LocalMux I__10896 (
            .O(N__46533),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    InMux I__10895 (
            .O(N__46526),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__10894 (
            .O(N__46523),
            .I(N__46520));
    InMux I__10893 (
            .O(N__46520),
            .I(N__46516));
    InMux I__10892 (
            .O(N__46519),
            .I(N__46513));
    LocalMux I__10891 (
            .O(N__46516),
            .I(N__46509));
    LocalMux I__10890 (
            .O(N__46513),
            .I(N__46506));
    InMux I__10889 (
            .O(N__46512),
            .I(N__46503));
    Span4Mux_h I__10888 (
            .O(N__46509),
            .I(N__46500));
    Span4Mux_h I__10887 (
            .O(N__46506),
            .I(N__46497));
    LocalMux I__10886 (
            .O(N__46503),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv4 I__10885 (
            .O(N__46500),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv4 I__10884 (
            .O(N__46497),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    CascadeMux I__10883 (
            .O(N__46490),
            .I(N__46487));
    InMux I__10882 (
            .O(N__46487),
            .I(N__46484));
    LocalMux I__10881 (
            .O(N__46484),
            .I(N__46479));
    InMux I__10880 (
            .O(N__46483),
            .I(N__46474));
    InMux I__10879 (
            .O(N__46482),
            .I(N__46474));
    Span4Mux_v I__10878 (
            .O(N__46479),
            .I(N__46468));
    LocalMux I__10877 (
            .O(N__46474),
            .I(N__46468));
    InMux I__10876 (
            .O(N__46473),
            .I(N__46465));
    Odrv4 I__10875 (
            .O(N__46468),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    LocalMux I__10874 (
            .O(N__46465),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    InMux I__10873 (
            .O(N__46460),
            .I(bfn_18_20_0_));
    CascadeMux I__10872 (
            .O(N__46457),
            .I(N__46454));
    InMux I__10871 (
            .O(N__46454),
            .I(N__46450));
    InMux I__10870 (
            .O(N__46453),
            .I(N__46447));
    LocalMux I__10869 (
            .O(N__46450),
            .I(N__46443));
    LocalMux I__10868 (
            .O(N__46447),
            .I(N__46440));
    InMux I__10867 (
            .O(N__46446),
            .I(N__46437));
    Span4Mux_h I__10866 (
            .O(N__46443),
            .I(N__46434));
    Span4Mux_h I__10865 (
            .O(N__46440),
            .I(N__46431));
    LocalMux I__10864 (
            .O(N__46437),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__10863 (
            .O(N__46434),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__10862 (
            .O(N__46431),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    InMux I__10861 (
            .O(N__46424),
            .I(N__46420));
    InMux I__10860 (
            .O(N__46423),
            .I(N__46416));
    LocalMux I__10859 (
            .O(N__46420),
            .I(N__46413));
    InMux I__10858 (
            .O(N__46419),
            .I(N__46409));
    LocalMux I__10857 (
            .O(N__46416),
            .I(N__46404));
    Span12Mux_v I__10856 (
            .O(N__46413),
            .I(N__46404));
    InMux I__10855 (
            .O(N__46412),
            .I(N__46401));
    LocalMux I__10854 (
            .O(N__46409),
            .I(N__46398));
    Odrv12 I__10853 (
            .O(N__46404),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    LocalMux I__10852 (
            .O(N__46401),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    Odrv4 I__10851 (
            .O(N__46398),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    InMux I__10850 (
            .O(N__46391),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__10849 (
            .O(N__46388),
            .I(N__46385));
    InMux I__10848 (
            .O(N__46385),
            .I(N__46380));
    InMux I__10847 (
            .O(N__46384),
            .I(N__46377));
    InMux I__10846 (
            .O(N__46383),
            .I(N__46374));
    LocalMux I__10845 (
            .O(N__46380),
            .I(N__46369));
    LocalMux I__10844 (
            .O(N__46377),
            .I(N__46369));
    LocalMux I__10843 (
            .O(N__46374),
            .I(N__46364));
    Span4Mux_v I__10842 (
            .O(N__46369),
            .I(N__46364));
    Odrv4 I__10841 (
            .O(N__46364),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    CascadeMux I__10840 (
            .O(N__46361),
            .I(N__46358));
    InMux I__10839 (
            .O(N__46358),
            .I(N__46355));
    LocalMux I__10838 (
            .O(N__46355),
            .I(N__46352));
    Span4Mux_h I__10837 (
            .O(N__46352),
            .I(N__46348));
    InMux I__10836 (
            .O(N__46351),
            .I(N__46345));
    Span4Mux_h I__10835 (
            .O(N__46348),
            .I(N__46340));
    LocalMux I__10834 (
            .O(N__46345),
            .I(N__46337));
    InMux I__10833 (
            .O(N__46344),
            .I(N__46334));
    InMux I__10832 (
            .O(N__46343),
            .I(N__46331));
    Odrv4 I__10831 (
            .O(N__46340),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    Odrv12 I__10830 (
            .O(N__46337),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    LocalMux I__10829 (
            .O(N__46334),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    LocalMux I__10828 (
            .O(N__46331),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    InMux I__10827 (
            .O(N__46322),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    InMux I__10826 (
            .O(N__46319),
            .I(N__46313));
    InMux I__10825 (
            .O(N__46318),
            .I(N__46313));
    LocalMux I__10824 (
            .O(N__46313),
            .I(N__46309));
    InMux I__10823 (
            .O(N__46312),
            .I(N__46306));
    Span4Mux_v I__10822 (
            .O(N__46309),
            .I(N__46303));
    LocalMux I__10821 (
            .O(N__46306),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    Odrv4 I__10820 (
            .O(N__46303),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__10819 (
            .O(N__46298),
            .I(N__46295));
    LocalMux I__10818 (
            .O(N__46295),
            .I(N__46289));
    InMux I__10817 (
            .O(N__46294),
            .I(N__46284));
    InMux I__10816 (
            .O(N__46293),
            .I(N__46284));
    InMux I__10815 (
            .O(N__46292),
            .I(N__46281));
    Span4Mux_v I__10814 (
            .O(N__46289),
            .I(N__46276));
    LocalMux I__10813 (
            .O(N__46284),
            .I(N__46276));
    LocalMux I__10812 (
            .O(N__46281),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    Odrv4 I__10811 (
            .O(N__46276),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    InMux I__10810 (
            .O(N__46271),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__10809 (
            .O(N__46268),
            .I(N__46265));
    InMux I__10808 (
            .O(N__46265),
            .I(N__46261));
    InMux I__10807 (
            .O(N__46264),
            .I(N__46258));
    LocalMux I__10806 (
            .O(N__46261),
            .I(N__46252));
    LocalMux I__10805 (
            .O(N__46258),
            .I(N__46252));
    InMux I__10804 (
            .O(N__46257),
            .I(N__46249));
    Span4Mux_h I__10803 (
            .O(N__46252),
            .I(N__46246));
    LocalMux I__10802 (
            .O(N__46249),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    Odrv4 I__10801 (
            .O(N__46246),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    CascadeMux I__10800 (
            .O(N__46241),
            .I(N__46238));
    InMux I__10799 (
            .O(N__46238),
            .I(N__46235));
    LocalMux I__10798 (
            .O(N__46235),
            .I(N__46231));
    InMux I__10797 (
            .O(N__46234),
            .I(N__46228));
    Span4Mux_h I__10796 (
            .O(N__46231),
            .I(N__46222));
    LocalMux I__10795 (
            .O(N__46228),
            .I(N__46222));
    InMux I__10794 (
            .O(N__46227),
            .I(N__46219));
    Span4Mux_v I__10793 (
            .O(N__46222),
            .I(N__46216));
    LocalMux I__10792 (
            .O(N__46219),
            .I(N__46212));
    Span4Mux_h I__10791 (
            .O(N__46216),
            .I(N__46209));
    InMux I__10790 (
            .O(N__46215),
            .I(N__46206));
    Odrv12 I__10789 (
            .O(N__46212),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    Odrv4 I__10788 (
            .O(N__46209),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    LocalMux I__10787 (
            .O(N__46206),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    InMux I__10786 (
            .O(N__46199),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__10785 (
            .O(N__46196),
            .I(N__46192));
    CascadeMux I__10784 (
            .O(N__46195),
            .I(N__46189));
    InMux I__10783 (
            .O(N__46192),
            .I(N__46184));
    InMux I__10782 (
            .O(N__46189),
            .I(N__46184));
    LocalMux I__10781 (
            .O(N__46184),
            .I(N__46180));
    InMux I__10780 (
            .O(N__46183),
            .I(N__46177));
    Span4Mux_h I__10779 (
            .O(N__46180),
            .I(N__46174));
    LocalMux I__10778 (
            .O(N__46177),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    Odrv4 I__10777 (
            .O(N__46174),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    CascadeMux I__10776 (
            .O(N__46169),
            .I(N__46166));
    InMux I__10775 (
            .O(N__46166),
            .I(N__46161));
    InMux I__10774 (
            .O(N__46165),
            .I(N__46158));
    InMux I__10773 (
            .O(N__46164),
            .I(N__46155));
    LocalMux I__10772 (
            .O(N__46161),
            .I(N__46151));
    LocalMux I__10771 (
            .O(N__46158),
            .I(N__46146));
    LocalMux I__10770 (
            .O(N__46155),
            .I(N__46146));
    InMux I__10769 (
            .O(N__46154),
            .I(N__46143));
    Odrv4 I__10768 (
            .O(N__46151),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    Odrv12 I__10767 (
            .O(N__46146),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    LocalMux I__10766 (
            .O(N__46143),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    InMux I__10765 (
            .O(N__46136),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    InMux I__10764 (
            .O(N__46133),
            .I(N__46127));
    InMux I__10763 (
            .O(N__46132),
            .I(N__46127));
    LocalMux I__10762 (
            .O(N__46127),
            .I(N__46123));
    InMux I__10761 (
            .O(N__46126),
            .I(N__46120));
    Span4Mux_h I__10760 (
            .O(N__46123),
            .I(N__46117));
    LocalMux I__10759 (
            .O(N__46120),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    Odrv4 I__10758 (
            .O(N__46117),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    CascadeMux I__10757 (
            .O(N__46112),
            .I(N__46107));
    InMux I__10756 (
            .O(N__46111),
            .I(N__46102));
    InMux I__10755 (
            .O(N__46110),
            .I(N__46102));
    InMux I__10754 (
            .O(N__46107),
            .I(N__46099));
    LocalMux I__10753 (
            .O(N__46102),
            .I(N__46096));
    LocalMux I__10752 (
            .O(N__46099),
            .I(N__46092));
    Span4Mux_v I__10751 (
            .O(N__46096),
            .I(N__46089));
    InMux I__10750 (
            .O(N__46095),
            .I(N__46086));
    Odrv4 I__10749 (
            .O(N__46092),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    Odrv4 I__10748 (
            .O(N__46089),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    LocalMux I__10747 (
            .O(N__46086),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    InMux I__10746 (
            .O(N__46079),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    InMux I__10745 (
            .O(N__46076),
            .I(N__46070));
    InMux I__10744 (
            .O(N__46075),
            .I(N__46070));
    LocalMux I__10743 (
            .O(N__46070),
            .I(N__46066));
    InMux I__10742 (
            .O(N__46069),
            .I(N__46063));
    Span4Mux_h I__10741 (
            .O(N__46066),
            .I(N__46060));
    LocalMux I__10740 (
            .O(N__46063),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    Odrv4 I__10739 (
            .O(N__46060),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__10738 (
            .O(N__46055),
            .I(N__46051));
    InMux I__10737 (
            .O(N__46054),
            .I(N__46047));
    LocalMux I__10736 (
            .O(N__46051),
            .I(N__46043));
    InMux I__10735 (
            .O(N__46050),
            .I(N__46040));
    LocalMux I__10734 (
            .O(N__46047),
            .I(N__46037));
    InMux I__10733 (
            .O(N__46046),
            .I(N__46034));
    Span4Mux_v I__10732 (
            .O(N__46043),
            .I(N__46029));
    LocalMux I__10731 (
            .O(N__46040),
            .I(N__46029));
    Odrv4 I__10730 (
            .O(N__46037),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    LocalMux I__10729 (
            .O(N__46034),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    Odrv4 I__10728 (
            .O(N__46029),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    InMux I__10727 (
            .O(N__46022),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    InMux I__10726 (
            .O(N__46019),
            .I(N__46015));
    InMux I__10725 (
            .O(N__46018),
            .I(N__46012));
    LocalMux I__10724 (
            .O(N__46015),
            .I(N__46009));
    LocalMux I__10723 (
            .O(N__46012),
            .I(N__46005));
    Span4Mux_v I__10722 (
            .O(N__46009),
            .I(N__46002));
    InMux I__10721 (
            .O(N__46008),
            .I(N__45999));
    Span4Mux_h I__10720 (
            .O(N__46005),
            .I(N__45996));
    Odrv4 I__10719 (
            .O(N__46002),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    LocalMux I__10718 (
            .O(N__45999),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    Odrv4 I__10717 (
            .O(N__45996),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    CascadeMux I__10716 (
            .O(N__45989),
            .I(N__45986));
    InMux I__10715 (
            .O(N__45986),
            .I(N__45979));
    InMux I__10714 (
            .O(N__45985),
            .I(N__45979));
    InMux I__10713 (
            .O(N__45984),
            .I(N__45976));
    LocalMux I__10712 (
            .O(N__45979),
            .I(N__45972));
    LocalMux I__10711 (
            .O(N__45976),
            .I(N__45969));
    InMux I__10710 (
            .O(N__45975),
            .I(N__45966));
    Span4Mux_v I__10709 (
            .O(N__45972),
            .I(N__45963));
    Span4Mux_h I__10708 (
            .O(N__45969),
            .I(N__45960));
    LocalMux I__10707 (
            .O(N__45966),
            .I(N__45957));
    Odrv4 I__10706 (
            .O(N__45963),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    Odrv4 I__10705 (
            .O(N__45960),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    Odrv12 I__10704 (
            .O(N__45957),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    InMux I__10703 (
            .O(N__45950),
            .I(N__45947));
    LocalMux I__10702 (
            .O(N__45947),
            .I(N__45943));
    InMux I__10701 (
            .O(N__45946),
            .I(N__45940));
    Span4Mux_v I__10700 (
            .O(N__45943),
            .I(N__45937));
    LocalMux I__10699 (
            .O(N__45940),
            .I(N__45933));
    Span4Mux_v I__10698 (
            .O(N__45937),
            .I(N__45930));
    InMux I__10697 (
            .O(N__45936),
            .I(N__45927));
    Span4Mux_h I__10696 (
            .O(N__45933),
            .I(N__45924));
    Odrv4 I__10695 (
            .O(N__45930),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    LocalMux I__10694 (
            .O(N__45927),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    Odrv4 I__10693 (
            .O(N__45924),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    CascadeMux I__10692 (
            .O(N__45917),
            .I(N__45912));
    InMux I__10691 (
            .O(N__45916),
            .I(N__45909));
    InMux I__10690 (
            .O(N__45915),
            .I(N__45906));
    InMux I__10689 (
            .O(N__45912),
            .I(N__45903));
    LocalMux I__10688 (
            .O(N__45909),
            .I(N__45900));
    LocalMux I__10687 (
            .O(N__45906),
            .I(N__45894));
    LocalMux I__10686 (
            .O(N__45903),
            .I(N__45894));
    Span4Mux_h I__10685 (
            .O(N__45900),
            .I(N__45891));
    InMux I__10684 (
            .O(N__45899),
            .I(N__45888));
    Span12Mux_v I__10683 (
            .O(N__45894),
            .I(N__45885));
    Span4Mux_h I__10682 (
            .O(N__45891),
            .I(N__45882));
    LocalMux I__10681 (
            .O(N__45888),
            .I(N__45879));
    Odrv12 I__10680 (
            .O(N__45885),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    Odrv4 I__10679 (
            .O(N__45882),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    Odrv12 I__10678 (
            .O(N__45879),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    InMux I__10677 (
            .O(N__45872),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__10676 (
            .O(N__45869),
            .I(N__45865));
    CascadeMux I__10675 (
            .O(N__45868),
            .I(N__45862));
    InMux I__10674 (
            .O(N__45865),
            .I(N__45856));
    InMux I__10673 (
            .O(N__45862),
            .I(N__45856));
    InMux I__10672 (
            .O(N__45861),
            .I(N__45853));
    LocalMux I__10671 (
            .O(N__45856),
            .I(N__45850));
    LocalMux I__10670 (
            .O(N__45853),
            .I(N__45845));
    Span4Mux_v I__10669 (
            .O(N__45850),
            .I(N__45845));
    Odrv4 I__10668 (
            .O(N__45845),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    InMux I__10667 (
            .O(N__45842),
            .I(N__45839));
    LocalMux I__10666 (
            .O(N__45839),
            .I(N__45833));
    InMux I__10665 (
            .O(N__45838),
            .I(N__45830));
    InMux I__10664 (
            .O(N__45837),
            .I(N__45827));
    InMux I__10663 (
            .O(N__45836),
            .I(N__45824));
    Span4Mux_h I__10662 (
            .O(N__45833),
            .I(N__45821));
    LocalMux I__10661 (
            .O(N__45830),
            .I(N__45818));
    LocalMux I__10660 (
            .O(N__45827),
            .I(N__45813));
    LocalMux I__10659 (
            .O(N__45824),
            .I(N__45813));
    Span4Mux_v I__10658 (
            .O(N__45821),
            .I(N__45810));
    Span4Mux_h I__10657 (
            .O(N__45818),
            .I(N__45807));
    Span4Mux_v I__10656 (
            .O(N__45813),
            .I(N__45804));
    Odrv4 I__10655 (
            .O(N__45810),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    Odrv4 I__10654 (
            .O(N__45807),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    Odrv4 I__10653 (
            .O(N__45804),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    InMux I__10652 (
            .O(N__45797),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__10651 (
            .O(N__45794),
            .I(N__45790));
    CascadeMux I__10650 (
            .O(N__45793),
            .I(N__45787));
    InMux I__10649 (
            .O(N__45790),
            .I(N__45782));
    InMux I__10648 (
            .O(N__45787),
            .I(N__45782));
    LocalMux I__10647 (
            .O(N__45782),
            .I(N__45778));
    InMux I__10646 (
            .O(N__45781),
            .I(N__45775));
    Span4Mux_v I__10645 (
            .O(N__45778),
            .I(N__45772));
    LocalMux I__10644 (
            .O(N__45775),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    Odrv4 I__10643 (
            .O(N__45772),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    CascadeMux I__10642 (
            .O(N__45767),
            .I(N__45764));
    InMux I__10641 (
            .O(N__45764),
            .I(N__45758));
    InMux I__10640 (
            .O(N__45763),
            .I(N__45758));
    LocalMux I__10639 (
            .O(N__45758),
            .I(N__45753));
    InMux I__10638 (
            .O(N__45757),
            .I(N__45750));
    InMux I__10637 (
            .O(N__45756),
            .I(N__45747));
    Span4Mux_h I__10636 (
            .O(N__45753),
            .I(N__45744));
    LocalMux I__10635 (
            .O(N__45750),
            .I(N__45741));
    LocalMux I__10634 (
            .O(N__45747),
            .I(N__45738));
    Span4Mux_v I__10633 (
            .O(N__45744),
            .I(N__45735));
    Span4Mux_h I__10632 (
            .O(N__45741),
            .I(N__45732));
    Span4Mux_v I__10631 (
            .O(N__45738),
            .I(N__45729));
    Odrv4 I__10630 (
            .O(N__45735),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    Odrv4 I__10629 (
            .O(N__45732),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    Odrv4 I__10628 (
            .O(N__45729),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    InMux I__10627 (
            .O(N__45722),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__10626 (
            .O(N__45719),
            .I(N__45716));
    InMux I__10625 (
            .O(N__45716),
            .I(N__45712));
    InMux I__10624 (
            .O(N__45715),
            .I(N__45709));
    LocalMux I__10623 (
            .O(N__45712),
            .I(N__45703));
    LocalMux I__10622 (
            .O(N__45709),
            .I(N__45703));
    InMux I__10621 (
            .O(N__45708),
            .I(N__45700));
    Span4Mux_h I__10620 (
            .O(N__45703),
            .I(N__45697));
    LocalMux I__10619 (
            .O(N__45700),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    Odrv4 I__10618 (
            .O(N__45697),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    CascadeMux I__10617 (
            .O(N__45692),
            .I(N__45688));
    InMux I__10616 (
            .O(N__45691),
            .I(N__45683));
    InMux I__10615 (
            .O(N__45688),
            .I(N__45683));
    LocalMux I__10614 (
            .O(N__45683),
            .I(N__45679));
    InMux I__10613 (
            .O(N__45682),
            .I(N__45676));
    Span4Mux_h I__10612 (
            .O(N__45679),
            .I(N__45673));
    LocalMux I__10611 (
            .O(N__45676),
            .I(N__45670));
    Span4Mux_v I__10610 (
            .O(N__45673),
            .I(N__45666));
    Span4Mux_h I__10609 (
            .O(N__45670),
            .I(N__45663));
    InMux I__10608 (
            .O(N__45669),
            .I(N__45660));
    Odrv4 I__10607 (
            .O(N__45666),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    Odrv4 I__10606 (
            .O(N__45663),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    LocalMux I__10605 (
            .O(N__45660),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    InMux I__10604 (
            .O(N__45653),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__10603 (
            .O(N__45650),
            .I(N__45647));
    InMux I__10602 (
            .O(N__45647),
            .I(N__45643));
    InMux I__10601 (
            .O(N__45646),
            .I(N__45640));
    LocalMux I__10600 (
            .O(N__45643),
            .I(N__45634));
    LocalMux I__10599 (
            .O(N__45640),
            .I(N__45634));
    InMux I__10598 (
            .O(N__45639),
            .I(N__45631));
    Span4Mux_h I__10597 (
            .O(N__45634),
            .I(N__45628));
    LocalMux I__10596 (
            .O(N__45631),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    Odrv4 I__10595 (
            .O(N__45628),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    CascadeMux I__10594 (
            .O(N__45623),
            .I(N__45619));
    CascadeMux I__10593 (
            .O(N__45622),
            .I(N__45616));
    InMux I__10592 (
            .O(N__45619),
            .I(N__45611));
    InMux I__10591 (
            .O(N__45616),
            .I(N__45611));
    LocalMux I__10590 (
            .O(N__45611),
            .I(N__45607));
    InMux I__10589 (
            .O(N__45610),
            .I(N__45604));
    Span4Mux_h I__10588 (
            .O(N__45607),
            .I(N__45600));
    LocalMux I__10587 (
            .O(N__45604),
            .I(N__45597));
    InMux I__10586 (
            .O(N__45603),
            .I(N__45594));
    Span4Mux_v I__10585 (
            .O(N__45600),
            .I(N__45591));
    Span4Mux_h I__10584 (
            .O(N__45597),
            .I(N__45588));
    LocalMux I__10583 (
            .O(N__45594),
            .I(N__45585));
    Odrv4 I__10582 (
            .O(N__45591),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    Odrv4 I__10581 (
            .O(N__45588),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    Odrv12 I__10580 (
            .O(N__45585),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    InMux I__10579 (
            .O(N__45578),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__10578 (
            .O(N__45575),
            .I(N__45572));
    InMux I__10577 (
            .O(N__45572),
            .I(N__45568));
    InMux I__10576 (
            .O(N__45571),
            .I(N__45565));
    LocalMux I__10575 (
            .O(N__45568),
            .I(N__45559));
    LocalMux I__10574 (
            .O(N__45565),
            .I(N__45559));
    InMux I__10573 (
            .O(N__45564),
            .I(N__45556));
    Span4Mux_h I__10572 (
            .O(N__45559),
            .I(N__45553));
    LocalMux I__10571 (
            .O(N__45556),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    Odrv4 I__10570 (
            .O(N__45553),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    CascadeMux I__10569 (
            .O(N__45548),
            .I(N__45545));
    InMux I__10568 (
            .O(N__45545),
            .I(N__45540));
    InMux I__10567 (
            .O(N__45544),
            .I(N__45535));
    InMux I__10566 (
            .O(N__45543),
            .I(N__45535));
    LocalMux I__10565 (
            .O(N__45540),
            .I(N__45530));
    LocalMux I__10564 (
            .O(N__45535),
            .I(N__45530));
    Span12Mux_v I__10563 (
            .O(N__45530),
            .I(N__45526));
    InMux I__10562 (
            .O(N__45529),
            .I(N__45523));
    Odrv12 I__10561 (
            .O(N__45526),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    LocalMux I__10560 (
            .O(N__45523),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    InMux I__10559 (
            .O(N__45518),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__10558 (
            .O(N__45515),
            .I(N__45512));
    InMux I__10557 (
            .O(N__45512),
            .I(N__45508));
    InMux I__10556 (
            .O(N__45511),
            .I(N__45505));
    LocalMux I__10555 (
            .O(N__45508),
            .I(N__45499));
    LocalMux I__10554 (
            .O(N__45505),
            .I(N__45499));
    InMux I__10553 (
            .O(N__45504),
            .I(N__45496));
    Span4Mux_h I__10552 (
            .O(N__45499),
            .I(N__45493));
    LocalMux I__10551 (
            .O(N__45496),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    Odrv4 I__10550 (
            .O(N__45493),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    CascadeMux I__10549 (
            .O(N__45488),
            .I(N__45485));
    InMux I__10548 (
            .O(N__45485),
            .I(N__45482));
    LocalMux I__10547 (
            .O(N__45482),
            .I(N__45479));
    Span4Mux_h I__10546 (
            .O(N__45479),
            .I(N__45474));
    InMux I__10545 (
            .O(N__45478),
            .I(N__45471));
    InMux I__10544 (
            .O(N__45477),
            .I(N__45467));
    Span4Mux_h I__10543 (
            .O(N__45474),
            .I(N__45464));
    LocalMux I__10542 (
            .O(N__45471),
            .I(N__45461));
    InMux I__10541 (
            .O(N__45470),
            .I(N__45458));
    LocalMux I__10540 (
            .O(N__45467),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    Odrv4 I__10539 (
            .O(N__45464),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    Odrv12 I__10538 (
            .O(N__45461),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    LocalMux I__10537 (
            .O(N__45458),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    InMux I__10536 (
            .O(N__45449),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__10535 (
            .O(N__45446),
            .I(N__45443));
    InMux I__10534 (
            .O(N__45443),
            .I(N__45440));
    LocalMux I__10533 (
            .O(N__45440),
            .I(N__45437));
    Span4Mux_h I__10532 (
            .O(N__45437),
            .I(N__45434));
    Span4Mux_v I__10531 (
            .O(N__45434),
            .I(N__45431));
    Odrv4 I__10530 (
            .O(N__45431),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ));
    CascadeMux I__10529 (
            .O(N__45428),
            .I(N__45425));
    InMux I__10528 (
            .O(N__45425),
            .I(N__45421));
    CascadeMux I__10527 (
            .O(N__45424),
            .I(N__45418));
    LocalMux I__10526 (
            .O(N__45421),
            .I(N__45414));
    InMux I__10525 (
            .O(N__45418),
            .I(N__45411));
    InMux I__10524 (
            .O(N__45417),
            .I(N__45408));
    Odrv4 I__10523 (
            .O(N__45414),
            .I(\current_shift_inst.un4_control_input1_14 ));
    LocalMux I__10522 (
            .O(N__45411),
            .I(\current_shift_inst.un4_control_input1_14 ));
    LocalMux I__10521 (
            .O(N__45408),
            .I(\current_shift_inst.un4_control_input1_14 ));
    CascadeMux I__10520 (
            .O(N__45401),
            .I(N__45398));
    InMux I__10519 (
            .O(N__45398),
            .I(N__45395));
    LocalMux I__10518 (
            .O(N__45395),
            .I(N__45392));
    Span4Mux_v I__10517 (
            .O(N__45392),
            .I(N__45389));
    Span4Mux_h I__10516 (
            .O(N__45389),
            .I(N__45386));
    Odrv4 I__10515 (
            .O(N__45386),
            .I(\current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ));
    InMux I__10514 (
            .O(N__45383),
            .I(N__45380));
    LocalMux I__10513 (
            .O(N__45380),
            .I(N__45377));
    Odrv4 I__10512 (
            .O(N__45377),
            .I(\current_shift_inst.un4_control_input_1_axb_9 ));
    InMux I__10511 (
            .O(N__45374),
            .I(N__45371));
    LocalMux I__10510 (
            .O(N__45371),
            .I(\current_shift_inst.un4_control_input_1_axb_17 ));
    InMux I__10509 (
            .O(N__45368),
            .I(N__45363));
    InMux I__10508 (
            .O(N__45367),
            .I(N__45360));
    InMux I__10507 (
            .O(N__45366),
            .I(N__45357));
    LocalMux I__10506 (
            .O(N__45363),
            .I(N__45354));
    LocalMux I__10505 (
            .O(N__45360),
            .I(\current_shift_inst.un4_control_input1_25 ));
    LocalMux I__10504 (
            .O(N__45357),
            .I(\current_shift_inst.un4_control_input1_25 ));
    Odrv4 I__10503 (
            .O(N__45354),
            .I(\current_shift_inst.un4_control_input1_25 ));
    CascadeMux I__10502 (
            .O(N__45347),
            .I(N__45344));
    InMux I__10501 (
            .O(N__45344),
            .I(N__45341));
    LocalMux I__10500 (
            .O(N__45341),
            .I(N__45338));
    Span4Mux_v I__10499 (
            .O(N__45338),
            .I(N__45335));
    Span4Mux_h I__10498 (
            .O(N__45335),
            .I(N__45332));
    Odrv4 I__10497 (
            .O(N__45332),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ));
    InMux I__10496 (
            .O(N__45329),
            .I(N__45326));
    LocalMux I__10495 (
            .O(N__45326),
            .I(\current_shift_inst.un4_control_input_1_axb_22 ));
    InMux I__10494 (
            .O(N__45323),
            .I(N__45320));
    LocalMux I__10493 (
            .O(N__45320),
            .I(N__45317));
    Span4Mux_v I__10492 (
            .O(N__45317),
            .I(N__45312));
    InMux I__10491 (
            .O(N__45316),
            .I(N__45309));
    InMux I__10490 (
            .O(N__45315),
            .I(N__45306));
    Span4Mux_h I__10489 (
            .O(N__45312),
            .I(N__45303));
    LocalMux I__10488 (
            .O(N__45309),
            .I(N__45300));
    LocalMux I__10487 (
            .O(N__45306),
            .I(\current_shift_inst.un4_control_input1_26 ));
    Odrv4 I__10486 (
            .O(N__45303),
            .I(\current_shift_inst.un4_control_input1_26 ));
    Odrv4 I__10485 (
            .O(N__45300),
            .I(\current_shift_inst.un4_control_input1_26 ));
    CascadeMux I__10484 (
            .O(N__45293),
            .I(N__45284));
    CascadeMux I__10483 (
            .O(N__45292),
            .I(N__45281));
    CascadeMux I__10482 (
            .O(N__45291),
            .I(N__45275));
    CascadeMux I__10481 (
            .O(N__45290),
            .I(N__45272));
    CascadeMux I__10480 (
            .O(N__45289),
            .I(N__45268));
    CascadeMux I__10479 (
            .O(N__45288),
            .I(N__45260));
    CascadeMux I__10478 (
            .O(N__45287),
            .I(N__45254));
    InMux I__10477 (
            .O(N__45284),
            .I(N__45248));
    InMux I__10476 (
            .O(N__45281),
            .I(N__45248));
    CascadeMux I__10475 (
            .O(N__45280),
            .I(N__45245));
    CascadeMux I__10474 (
            .O(N__45279),
            .I(N__45242));
    CascadeMux I__10473 (
            .O(N__45278),
            .I(N__45238));
    InMux I__10472 (
            .O(N__45275),
            .I(N__45227));
    InMux I__10471 (
            .O(N__45272),
            .I(N__45227));
    InMux I__10470 (
            .O(N__45271),
            .I(N__45216));
    InMux I__10469 (
            .O(N__45268),
            .I(N__45216));
    InMux I__10468 (
            .O(N__45267),
            .I(N__45216));
    InMux I__10467 (
            .O(N__45266),
            .I(N__45216));
    InMux I__10466 (
            .O(N__45265),
            .I(N__45216));
    CascadeMux I__10465 (
            .O(N__45264),
            .I(N__45212));
    CascadeMux I__10464 (
            .O(N__45263),
            .I(N__45203));
    InMux I__10463 (
            .O(N__45260),
            .I(N__45195));
    InMux I__10462 (
            .O(N__45259),
            .I(N__45190));
    InMux I__10461 (
            .O(N__45258),
            .I(N__45190));
    InMux I__10460 (
            .O(N__45257),
            .I(N__45185));
    InMux I__10459 (
            .O(N__45254),
            .I(N__45185));
    CascadeMux I__10458 (
            .O(N__45253),
            .I(N__45182));
    LocalMux I__10457 (
            .O(N__45248),
            .I(N__45173));
    InMux I__10456 (
            .O(N__45245),
            .I(N__45170));
    InMux I__10455 (
            .O(N__45242),
            .I(N__45163));
    InMux I__10454 (
            .O(N__45241),
            .I(N__45163));
    InMux I__10453 (
            .O(N__45238),
            .I(N__45163));
    InMux I__10452 (
            .O(N__45237),
            .I(N__45152));
    InMux I__10451 (
            .O(N__45236),
            .I(N__45152));
    InMux I__10450 (
            .O(N__45235),
            .I(N__45152));
    InMux I__10449 (
            .O(N__45234),
            .I(N__45152));
    InMux I__10448 (
            .O(N__45233),
            .I(N__45152));
    CascadeMux I__10447 (
            .O(N__45232),
            .I(N__45149));
    LocalMux I__10446 (
            .O(N__45227),
            .I(N__45120));
    LocalMux I__10445 (
            .O(N__45216),
            .I(N__45120));
    InMux I__10444 (
            .O(N__45215),
            .I(N__45113));
    InMux I__10443 (
            .O(N__45212),
            .I(N__45113));
    InMux I__10442 (
            .O(N__45211),
            .I(N__45113));
    InMux I__10441 (
            .O(N__45210),
            .I(N__45102));
    InMux I__10440 (
            .O(N__45209),
            .I(N__45102));
    InMux I__10439 (
            .O(N__45208),
            .I(N__45102));
    InMux I__10438 (
            .O(N__45207),
            .I(N__45102));
    InMux I__10437 (
            .O(N__45206),
            .I(N__45102));
    InMux I__10436 (
            .O(N__45203),
            .I(N__45099));
    CascadeMux I__10435 (
            .O(N__45202),
            .I(N__45095));
    CascadeMux I__10434 (
            .O(N__45201),
            .I(N__45092));
    InMux I__10433 (
            .O(N__45200),
            .I(N__45085));
    InMux I__10432 (
            .O(N__45199),
            .I(N__45085));
    InMux I__10431 (
            .O(N__45198),
            .I(N__45085));
    LocalMux I__10430 (
            .O(N__45195),
            .I(N__45080));
    LocalMux I__10429 (
            .O(N__45190),
            .I(N__45080));
    LocalMux I__10428 (
            .O(N__45185),
            .I(N__45077));
    InMux I__10427 (
            .O(N__45182),
            .I(N__45074));
    InMux I__10426 (
            .O(N__45181),
            .I(N__45071));
    CascadeMux I__10425 (
            .O(N__45180),
            .I(N__45067));
    CascadeMux I__10424 (
            .O(N__45179),
            .I(N__45062));
    CascadeMux I__10423 (
            .O(N__45178),
            .I(N__45055));
    CascadeMux I__10422 (
            .O(N__45177),
            .I(N__45052));
    CascadeMux I__10421 (
            .O(N__45176),
            .I(N__45048));
    Span4Mux_v I__10420 (
            .O(N__45173),
            .I(N__45032));
    LocalMux I__10419 (
            .O(N__45170),
            .I(N__45032));
    LocalMux I__10418 (
            .O(N__45163),
            .I(N__45032));
    LocalMux I__10417 (
            .O(N__45152),
            .I(N__45032));
    InMux I__10416 (
            .O(N__45149),
            .I(N__45023));
    InMux I__10415 (
            .O(N__45148),
            .I(N__45023));
    InMux I__10414 (
            .O(N__45147),
            .I(N__45023));
    InMux I__10413 (
            .O(N__45146),
            .I(N__45023));
    CascadeMux I__10412 (
            .O(N__45145),
            .I(N__45019));
    CascadeMux I__10411 (
            .O(N__45144),
            .I(N__45015));
    CascadeMux I__10410 (
            .O(N__45143),
            .I(N__45011));
    CascadeMux I__10409 (
            .O(N__45142),
            .I(N__45005));
    CascadeMux I__10408 (
            .O(N__45141),
            .I(N__45001));
    CascadeMux I__10407 (
            .O(N__45140),
            .I(N__44997));
    CascadeMux I__10406 (
            .O(N__45139),
            .I(N__44992));
    CascadeMux I__10405 (
            .O(N__45138),
            .I(N__44988));
    CascadeMux I__10404 (
            .O(N__45137),
            .I(N__44984));
    CascadeMux I__10403 (
            .O(N__45136),
            .I(N__44980));
    CascadeMux I__10402 (
            .O(N__45135),
            .I(N__44977));
    CascadeMux I__10401 (
            .O(N__45134),
            .I(N__44973));
    CascadeMux I__10400 (
            .O(N__45133),
            .I(N__44969));
    CascadeMux I__10399 (
            .O(N__45132),
            .I(N__44965));
    CascadeMux I__10398 (
            .O(N__45131),
            .I(N__44961));
    CascadeMux I__10397 (
            .O(N__45130),
            .I(N__44957));
    CascadeMux I__10396 (
            .O(N__45129),
            .I(N__44953));
    CascadeMux I__10395 (
            .O(N__45128),
            .I(N__44949));
    CascadeMux I__10394 (
            .O(N__45127),
            .I(N__44945));
    CascadeMux I__10393 (
            .O(N__45126),
            .I(N__44941));
    CascadeMux I__10392 (
            .O(N__45125),
            .I(N__44937));
    Span4Mux_v I__10391 (
            .O(N__45120),
            .I(N__44931));
    LocalMux I__10390 (
            .O(N__45113),
            .I(N__44931));
    LocalMux I__10389 (
            .O(N__45102),
            .I(N__44928));
    LocalMux I__10388 (
            .O(N__45099),
            .I(N__44925));
    InMux I__10387 (
            .O(N__45098),
            .I(N__44922));
    InMux I__10386 (
            .O(N__45095),
            .I(N__44917));
    InMux I__10385 (
            .O(N__45092),
            .I(N__44917));
    LocalMux I__10384 (
            .O(N__45085),
            .I(N__44914));
    Span4Mux_v I__10383 (
            .O(N__45080),
            .I(N__44905));
    Span4Mux_v I__10382 (
            .O(N__45077),
            .I(N__44905));
    LocalMux I__10381 (
            .O(N__45074),
            .I(N__44905));
    LocalMux I__10380 (
            .O(N__45071),
            .I(N__44905));
    CascadeMux I__10379 (
            .O(N__45070),
            .I(N__44902));
    InMux I__10378 (
            .O(N__45067),
            .I(N__44893));
    InMux I__10377 (
            .O(N__45066),
            .I(N__44893));
    InMux I__10376 (
            .O(N__45065),
            .I(N__44893));
    InMux I__10375 (
            .O(N__45062),
            .I(N__44893));
    InMux I__10374 (
            .O(N__45061),
            .I(N__44876));
    InMux I__10373 (
            .O(N__45060),
            .I(N__44876));
    InMux I__10372 (
            .O(N__45059),
            .I(N__44876));
    InMux I__10371 (
            .O(N__45058),
            .I(N__44876));
    InMux I__10370 (
            .O(N__45055),
            .I(N__44876));
    InMux I__10369 (
            .O(N__45052),
            .I(N__44876));
    InMux I__10368 (
            .O(N__45051),
            .I(N__44876));
    InMux I__10367 (
            .O(N__45048),
            .I(N__44876));
    CascadeMux I__10366 (
            .O(N__45047),
            .I(N__44872));
    CascadeMux I__10365 (
            .O(N__45046),
            .I(N__44868));
    CascadeMux I__10364 (
            .O(N__45045),
            .I(N__44864));
    CascadeMux I__10363 (
            .O(N__45044),
            .I(N__44860));
    CascadeMux I__10362 (
            .O(N__45043),
            .I(N__44857));
    CascadeMux I__10361 (
            .O(N__45042),
            .I(N__44853));
    CascadeMux I__10360 (
            .O(N__45041),
            .I(N__44849));
    Span4Mux_v I__10359 (
            .O(N__45032),
            .I(N__44843));
    LocalMux I__10358 (
            .O(N__45023),
            .I(N__44843));
    InMux I__10357 (
            .O(N__45022),
            .I(N__44828));
    InMux I__10356 (
            .O(N__45019),
            .I(N__44828));
    InMux I__10355 (
            .O(N__45018),
            .I(N__44828));
    InMux I__10354 (
            .O(N__45015),
            .I(N__44828));
    InMux I__10353 (
            .O(N__45014),
            .I(N__44828));
    InMux I__10352 (
            .O(N__45011),
            .I(N__44828));
    InMux I__10351 (
            .O(N__45010),
            .I(N__44828));
    InMux I__10350 (
            .O(N__45009),
            .I(N__44811));
    InMux I__10349 (
            .O(N__45008),
            .I(N__44811));
    InMux I__10348 (
            .O(N__45005),
            .I(N__44811));
    InMux I__10347 (
            .O(N__45004),
            .I(N__44811));
    InMux I__10346 (
            .O(N__45001),
            .I(N__44811));
    InMux I__10345 (
            .O(N__45000),
            .I(N__44811));
    InMux I__10344 (
            .O(N__44997),
            .I(N__44811));
    InMux I__10343 (
            .O(N__44996),
            .I(N__44811));
    InMux I__10342 (
            .O(N__44995),
            .I(N__44794));
    InMux I__10341 (
            .O(N__44992),
            .I(N__44794));
    InMux I__10340 (
            .O(N__44991),
            .I(N__44794));
    InMux I__10339 (
            .O(N__44988),
            .I(N__44794));
    InMux I__10338 (
            .O(N__44987),
            .I(N__44794));
    InMux I__10337 (
            .O(N__44984),
            .I(N__44794));
    InMux I__10336 (
            .O(N__44983),
            .I(N__44794));
    InMux I__10335 (
            .O(N__44980),
            .I(N__44794));
    InMux I__10334 (
            .O(N__44977),
            .I(N__44777));
    InMux I__10333 (
            .O(N__44976),
            .I(N__44777));
    InMux I__10332 (
            .O(N__44973),
            .I(N__44777));
    InMux I__10331 (
            .O(N__44972),
            .I(N__44777));
    InMux I__10330 (
            .O(N__44969),
            .I(N__44777));
    InMux I__10329 (
            .O(N__44968),
            .I(N__44777));
    InMux I__10328 (
            .O(N__44965),
            .I(N__44777));
    InMux I__10327 (
            .O(N__44964),
            .I(N__44777));
    InMux I__10326 (
            .O(N__44961),
            .I(N__44760));
    InMux I__10325 (
            .O(N__44960),
            .I(N__44760));
    InMux I__10324 (
            .O(N__44957),
            .I(N__44760));
    InMux I__10323 (
            .O(N__44956),
            .I(N__44760));
    InMux I__10322 (
            .O(N__44953),
            .I(N__44760));
    InMux I__10321 (
            .O(N__44952),
            .I(N__44760));
    InMux I__10320 (
            .O(N__44949),
            .I(N__44760));
    InMux I__10319 (
            .O(N__44948),
            .I(N__44760));
    InMux I__10318 (
            .O(N__44945),
            .I(N__44747));
    InMux I__10317 (
            .O(N__44944),
            .I(N__44747));
    InMux I__10316 (
            .O(N__44941),
            .I(N__44747));
    InMux I__10315 (
            .O(N__44940),
            .I(N__44747));
    InMux I__10314 (
            .O(N__44937),
            .I(N__44747));
    InMux I__10313 (
            .O(N__44936),
            .I(N__44747));
    Span4Mux_h I__10312 (
            .O(N__44931),
            .I(N__44744));
    Span4Mux_v I__10311 (
            .O(N__44928),
            .I(N__44735));
    Span4Mux_v I__10310 (
            .O(N__44925),
            .I(N__44735));
    LocalMux I__10309 (
            .O(N__44922),
            .I(N__44735));
    LocalMux I__10308 (
            .O(N__44917),
            .I(N__44735));
    Span4Mux_v I__10307 (
            .O(N__44914),
            .I(N__44730));
    Span4Mux_v I__10306 (
            .O(N__44905),
            .I(N__44730));
    InMux I__10305 (
            .O(N__44902),
            .I(N__44727));
    LocalMux I__10304 (
            .O(N__44893),
            .I(N__44722));
    LocalMux I__10303 (
            .O(N__44876),
            .I(N__44722));
    InMux I__10302 (
            .O(N__44875),
            .I(N__44705));
    InMux I__10301 (
            .O(N__44872),
            .I(N__44705));
    InMux I__10300 (
            .O(N__44871),
            .I(N__44705));
    InMux I__10299 (
            .O(N__44868),
            .I(N__44705));
    InMux I__10298 (
            .O(N__44867),
            .I(N__44705));
    InMux I__10297 (
            .O(N__44864),
            .I(N__44705));
    InMux I__10296 (
            .O(N__44863),
            .I(N__44705));
    InMux I__10295 (
            .O(N__44860),
            .I(N__44705));
    InMux I__10294 (
            .O(N__44857),
            .I(N__44692));
    InMux I__10293 (
            .O(N__44856),
            .I(N__44692));
    InMux I__10292 (
            .O(N__44853),
            .I(N__44692));
    InMux I__10291 (
            .O(N__44852),
            .I(N__44692));
    InMux I__10290 (
            .O(N__44849),
            .I(N__44692));
    InMux I__10289 (
            .O(N__44848),
            .I(N__44692));
    Sp12to4 I__10288 (
            .O(N__44843),
            .I(N__44677));
    LocalMux I__10287 (
            .O(N__44828),
            .I(N__44677));
    LocalMux I__10286 (
            .O(N__44811),
            .I(N__44677));
    LocalMux I__10285 (
            .O(N__44794),
            .I(N__44677));
    LocalMux I__10284 (
            .O(N__44777),
            .I(N__44677));
    LocalMux I__10283 (
            .O(N__44760),
            .I(N__44677));
    LocalMux I__10282 (
            .O(N__44747),
            .I(N__44677));
    Odrv4 I__10281 (
            .O(N__44744),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10280 (
            .O(N__44735),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10279 (
            .O(N__44730),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10278 (
            .O(N__44727),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv12 I__10277 (
            .O(N__44722),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10276 (
            .O(N__44705),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10275 (
            .O(N__44692),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv12 I__10274 (
            .O(N__44677),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    InMux I__10273 (
            .O(N__44660),
            .I(N__44639));
    InMux I__10272 (
            .O(N__44659),
            .I(N__44639));
    InMux I__10271 (
            .O(N__44658),
            .I(N__44630));
    InMux I__10270 (
            .O(N__44657),
            .I(N__44630));
    InMux I__10269 (
            .O(N__44656),
            .I(N__44630));
    InMux I__10268 (
            .O(N__44655),
            .I(N__44630));
    InMux I__10267 (
            .O(N__44654),
            .I(N__44615));
    InMux I__10266 (
            .O(N__44653),
            .I(N__44612));
    InMux I__10265 (
            .O(N__44652),
            .I(N__44606));
    InMux I__10264 (
            .O(N__44651),
            .I(N__44595));
    InMux I__10263 (
            .O(N__44650),
            .I(N__44595));
    InMux I__10262 (
            .O(N__44649),
            .I(N__44595));
    InMux I__10261 (
            .O(N__44648),
            .I(N__44595));
    InMux I__10260 (
            .O(N__44647),
            .I(N__44595));
    InMux I__10259 (
            .O(N__44646),
            .I(N__44587));
    InMux I__10258 (
            .O(N__44645),
            .I(N__44583));
    InMux I__10257 (
            .O(N__44644),
            .I(N__44580));
    LocalMux I__10256 (
            .O(N__44639),
            .I(N__44568));
    LocalMux I__10255 (
            .O(N__44630),
            .I(N__44568));
    InMux I__10254 (
            .O(N__44629),
            .I(N__44557));
    InMux I__10253 (
            .O(N__44628),
            .I(N__44557));
    InMux I__10252 (
            .O(N__44627),
            .I(N__44557));
    InMux I__10251 (
            .O(N__44626),
            .I(N__44557));
    InMux I__10250 (
            .O(N__44625),
            .I(N__44557));
    InMux I__10249 (
            .O(N__44624),
            .I(N__44554));
    InMux I__10248 (
            .O(N__44623),
            .I(N__44547));
    InMux I__10247 (
            .O(N__44622),
            .I(N__44547));
    InMux I__10246 (
            .O(N__44621),
            .I(N__44547));
    InMux I__10245 (
            .O(N__44620),
            .I(N__44540));
    InMux I__10244 (
            .O(N__44619),
            .I(N__44540));
    InMux I__10243 (
            .O(N__44618),
            .I(N__44540));
    LocalMux I__10242 (
            .O(N__44615),
            .I(N__44535));
    LocalMux I__10241 (
            .O(N__44612),
            .I(N__44535));
    InMux I__10240 (
            .O(N__44611),
            .I(N__44531));
    InMux I__10239 (
            .O(N__44610),
            .I(N__44528));
    InMux I__10238 (
            .O(N__44609),
            .I(N__44525));
    LocalMux I__10237 (
            .O(N__44606),
            .I(N__44520));
    LocalMux I__10236 (
            .O(N__44595),
            .I(N__44520));
    InMux I__10235 (
            .O(N__44594),
            .I(N__44509));
    InMux I__10234 (
            .O(N__44593),
            .I(N__44509));
    InMux I__10233 (
            .O(N__44592),
            .I(N__44509));
    InMux I__10232 (
            .O(N__44591),
            .I(N__44509));
    InMux I__10231 (
            .O(N__44590),
            .I(N__44509));
    LocalMux I__10230 (
            .O(N__44587),
            .I(N__44506));
    InMux I__10229 (
            .O(N__44586),
            .I(N__44503));
    LocalMux I__10228 (
            .O(N__44583),
            .I(N__44500));
    LocalMux I__10227 (
            .O(N__44580),
            .I(N__44497));
    InMux I__10226 (
            .O(N__44579),
            .I(N__44492));
    InMux I__10225 (
            .O(N__44578),
            .I(N__44492));
    InMux I__10224 (
            .O(N__44577),
            .I(N__44481));
    InMux I__10223 (
            .O(N__44576),
            .I(N__44481));
    InMux I__10222 (
            .O(N__44575),
            .I(N__44481));
    InMux I__10221 (
            .O(N__44574),
            .I(N__44481));
    InMux I__10220 (
            .O(N__44573),
            .I(N__44481));
    Span4Mux_v I__10219 (
            .O(N__44568),
            .I(N__44471));
    LocalMux I__10218 (
            .O(N__44557),
            .I(N__44471));
    LocalMux I__10217 (
            .O(N__44554),
            .I(N__44466));
    LocalMux I__10216 (
            .O(N__44547),
            .I(N__44466));
    LocalMux I__10215 (
            .O(N__44540),
            .I(N__44458));
    Span4Mux_v I__10214 (
            .O(N__44535),
            .I(N__44458));
    InMux I__10213 (
            .O(N__44534),
            .I(N__44453));
    LocalMux I__10212 (
            .O(N__44531),
            .I(N__44442));
    LocalMux I__10211 (
            .O(N__44528),
            .I(N__44442));
    LocalMux I__10210 (
            .O(N__44525),
            .I(N__44442));
    Span4Mux_h I__10209 (
            .O(N__44520),
            .I(N__44442));
    LocalMux I__10208 (
            .O(N__44509),
            .I(N__44442));
    Span4Mux_v I__10207 (
            .O(N__44506),
            .I(N__44437));
    LocalMux I__10206 (
            .O(N__44503),
            .I(N__44437));
    Span4Mux_v I__10205 (
            .O(N__44500),
            .I(N__44428));
    Span4Mux_v I__10204 (
            .O(N__44497),
            .I(N__44428));
    LocalMux I__10203 (
            .O(N__44492),
            .I(N__44428));
    LocalMux I__10202 (
            .O(N__44481),
            .I(N__44428));
    CascadeMux I__10201 (
            .O(N__44480),
            .I(N__44414));
    CascadeMux I__10200 (
            .O(N__44479),
            .I(N__44409));
    InMux I__10199 (
            .O(N__44478),
            .I(N__44401));
    InMux I__10198 (
            .O(N__44477),
            .I(N__44401));
    InMux I__10197 (
            .O(N__44476),
            .I(N__44401));
    Span4Mux_h I__10196 (
            .O(N__44471),
            .I(N__44396));
    Span4Mux_v I__10195 (
            .O(N__44466),
            .I(N__44396));
    InMux I__10194 (
            .O(N__44465),
            .I(N__44389));
    InMux I__10193 (
            .O(N__44464),
            .I(N__44389));
    InMux I__10192 (
            .O(N__44463),
            .I(N__44389));
    Span4Mux_v I__10191 (
            .O(N__44458),
            .I(N__44386));
    InMux I__10190 (
            .O(N__44457),
            .I(N__44381));
    InMux I__10189 (
            .O(N__44456),
            .I(N__44381));
    LocalMux I__10188 (
            .O(N__44453),
            .I(N__44376));
    Span4Mux_v I__10187 (
            .O(N__44442),
            .I(N__44376));
    Span4Mux_v I__10186 (
            .O(N__44437),
            .I(N__44371));
    Span4Mux_v I__10185 (
            .O(N__44428),
            .I(N__44371));
    InMux I__10184 (
            .O(N__44427),
            .I(N__44364));
    InMux I__10183 (
            .O(N__44426),
            .I(N__44364));
    InMux I__10182 (
            .O(N__44425),
            .I(N__44364));
    InMux I__10181 (
            .O(N__44424),
            .I(N__44353));
    InMux I__10180 (
            .O(N__44423),
            .I(N__44353));
    InMux I__10179 (
            .O(N__44422),
            .I(N__44353));
    InMux I__10178 (
            .O(N__44421),
            .I(N__44353));
    InMux I__10177 (
            .O(N__44420),
            .I(N__44353));
    InMux I__10176 (
            .O(N__44419),
            .I(N__44348));
    InMux I__10175 (
            .O(N__44418),
            .I(N__44348));
    InMux I__10174 (
            .O(N__44417),
            .I(N__44345));
    InMux I__10173 (
            .O(N__44414),
            .I(N__44334));
    InMux I__10172 (
            .O(N__44413),
            .I(N__44334));
    InMux I__10171 (
            .O(N__44412),
            .I(N__44334));
    InMux I__10170 (
            .O(N__44409),
            .I(N__44334));
    InMux I__10169 (
            .O(N__44408),
            .I(N__44334));
    LocalMux I__10168 (
            .O(N__44401),
            .I(N__44327));
    Span4Mux_h I__10167 (
            .O(N__44396),
            .I(N__44327));
    LocalMux I__10166 (
            .O(N__44389),
            .I(N__44327));
    Odrv4 I__10165 (
            .O(N__44386),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10164 (
            .O(N__44381),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10163 (
            .O(N__44376),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10162 (
            .O(N__44371),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10161 (
            .O(N__44364),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10160 (
            .O(N__44353),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10159 (
            .O(N__44348),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10158 (
            .O(N__44345),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10157 (
            .O(N__44334),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10156 (
            .O(N__44327),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    InMux I__10155 (
            .O(N__44306),
            .I(N__44303));
    LocalMux I__10154 (
            .O(N__44303),
            .I(N__44300));
    Span4Mux_h I__10153 (
            .O(N__44300),
            .I(N__44297));
    Odrv4 I__10152 (
            .O(N__44297),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ));
    InMux I__10151 (
            .O(N__44294),
            .I(N__44291));
    LocalMux I__10150 (
            .O(N__44291),
            .I(N__44288));
    Span4Mux_h I__10149 (
            .O(N__44288),
            .I(N__44285));
    Odrv4 I__10148 (
            .O(N__44285),
            .I(\current_shift_inst.un4_control_input_1_axb_6 ));
    InMux I__10147 (
            .O(N__44282),
            .I(N__44279));
    LocalMux I__10146 (
            .O(N__44279),
            .I(N__44276));
    Span4Mux_h I__10145 (
            .O(N__44276),
            .I(N__44273));
    Odrv4 I__10144 (
            .O(N__44273),
            .I(\current_shift_inst.un4_control_input_1_axb_8 ));
    CascadeMux I__10143 (
            .O(N__44270),
            .I(N__44267));
    InMux I__10142 (
            .O(N__44267),
            .I(N__44264));
    LocalMux I__10141 (
            .O(N__44264),
            .I(N__44261));
    Span4Mux_h I__10140 (
            .O(N__44261),
            .I(N__44258));
    Odrv4 I__10139 (
            .O(N__44258),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ));
    InMux I__10138 (
            .O(N__44255),
            .I(N__44249));
    InMux I__10137 (
            .O(N__44254),
            .I(N__44249));
    LocalMux I__10136 (
            .O(N__44249),
            .I(N__44246));
    Odrv4 I__10135 (
            .O(N__44246),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    CascadeMux I__10134 (
            .O(N__44243),
            .I(N__44239));
    CascadeMux I__10133 (
            .O(N__44242),
            .I(N__44236));
    InMux I__10132 (
            .O(N__44239),
            .I(N__44233));
    InMux I__10131 (
            .O(N__44236),
            .I(N__44230));
    LocalMux I__10130 (
            .O(N__44233),
            .I(N__44227));
    LocalMux I__10129 (
            .O(N__44230),
            .I(N__44224));
    Span4Mux_v I__10128 (
            .O(N__44227),
            .I(N__44219));
    Span4Mux_v I__10127 (
            .O(N__44224),
            .I(N__44219));
    Span4Mux_h I__10126 (
            .O(N__44219),
            .I(N__44216));
    Odrv4 I__10125 (
            .O(N__44216),
            .I(\current_shift_inst.un4_control_input_0_31 ));
    InMux I__10124 (
            .O(N__44213),
            .I(N__44210));
    LocalMux I__10123 (
            .O(N__44210),
            .I(N__44207));
    Span4Mux_h I__10122 (
            .O(N__44207),
            .I(N__44204));
    Odrv4 I__10121 (
            .O(N__44204),
            .I(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ));
    InMux I__10120 (
            .O(N__44201),
            .I(N__44198));
    LocalMux I__10119 (
            .O(N__44198),
            .I(N__44194));
    InMux I__10118 (
            .O(N__44197),
            .I(N__44190));
    Span4Mux_h I__10117 (
            .O(N__44194),
            .I(N__44187));
    InMux I__10116 (
            .O(N__44193),
            .I(N__44184));
    LocalMux I__10115 (
            .O(N__44190),
            .I(\current_shift_inst.un4_control_input1_27 ));
    Odrv4 I__10114 (
            .O(N__44187),
            .I(\current_shift_inst.un4_control_input1_27 ));
    LocalMux I__10113 (
            .O(N__44184),
            .I(\current_shift_inst.un4_control_input1_27 ));
    CascadeMux I__10112 (
            .O(N__44177),
            .I(N__44174));
    InMux I__10111 (
            .O(N__44174),
            .I(N__44171));
    LocalMux I__10110 (
            .O(N__44171),
            .I(N__44168));
    Odrv12 I__10109 (
            .O(N__44168),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ));
    InMux I__10108 (
            .O(N__44165),
            .I(N__44162));
    LocalMux I__10107 (
            .O(N__44162),
            .I(\current_shift_inst.un4_control_input_1_axb_11 ));
    CascadeMux I__10106 (
            .O(N__44159),
            .I(N__44156));
    InMux I__10105 (
            .O(N__44156),
            .I(N__44152));
    CascadeMux I__10104 (
            .O(N__44155),
            .I(N__44149));
    LocalMux I__10103 (
            .O(N__44152),
            .I(N__44146));
    InMux I__10102 (
            .O(N__44149),
            .I(N__44142));
    Span4Mux_h I__10101 (
            .O(N__44146),
            .I(N__44139));
    InMux I__10100 (
            .O(N__44145),
            .I(N__44136));
    LocalMux I__10099 (
            .O(N__44142),
            .I(\current_shift_inst.un4_control_input1_30 ));
    Odrv4 I__10098 (
            .O(N__44139),
            .I(\current_shift_inst.un4_control_input1_30 ));
    LocalMux I__10097 (
            .O(N__44136),
            .I(\current_shift_inst.un4_control_input1_30 ));
    InMux I__10096 (
            .O(N__44129),
            .I(N__44126));
    LocalMux I__10095 (
            .O(N__44126),
            .I(N__44123));
    Odrv12 I__10094 (
            .O(N__44123),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ));
    InMux I__10093 (
            .O(N__44120),
            .I(N__44117));
    LocalMux I__10092 (
            .O(N__44117),
            .I(\current_shift_inst.un4_control_input_1_axb_13 ));
    CascadeMux I__10091 (
            .O(N__44114),
            .I(N__44111));
    InMux I__10090 (
            .O(N__44111),
            .I(N__44108));
    LocalMux I__10089 (
            .O(N__44108),
            .I(N__44105));
    Span4Mux_v I__10088 (
            .O(N__44105),
            .I(N__44102));
    Odrv4 I__10087 (
            .O(N__44102),
            .I(\current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ));
    InMux I__10086 (
            .O(N__44099),
            .I(N__44095));
    CascadeMux I__10085 (
            .O(N__44098),
            .I(N__44089));
    LocalMux I__10084 (
            .O(N__44095),
            .I(N__44072));
    InMux I__10083 (
            .O(N__44094),
            .I(N__44067));
    InMux I__10082 (
            .O(N__44093),
            .I(N__44067));
    InMux I__10081 (
            .O(N__44092),
            .I(N__44062));
    InMux I__10080 (
            .O(N__44089),
            .I(N__44055));
    InMux I__10079 (
            .O(N__44088),
            .I(N__44055));
    InMux I__10078 (
            .O(N__44087),
            .I(N__44055));
    InMux I__10077 (
            .O(N__44086),
            .I(N__44052));
    InMux I__10076 (
            .O(N__44085),
            .I(N__44037));
    InMux I__10075 (
            .O(N__44084),
            .I(N__44037));
    InMux I__10074 (
            .O(N__44083),
            .I(N__44037));
    InMux I__10073 (
            .O(N__44082),
            .I(N__44037));
    InMux I__10072 (
            .O(N__44081),
            .I(N__44037));
    InMux I__10071 (
            .O(N__44080),
            .I(N__44037));
    InMux I__10070 (
            .O(N__44079),
            .I(N__44037));
    InMux I__10069 (
            .O(N__44078),
            .I(N__44034));
    InMux I__10068 (
            .O(N__44077),
            .I(N__44031));
    InMux I__10067 (
            .O(N__44076),
            .I(N__44026));
    InMux I__10066 (
            .O(N__44075),
            .I(N__44026));
    Span4Mux_v I__10065 (
            .O(N__44072),
            .I(N__44020));
    LocalMux I__10064 (
            .O(N__44067),
            .I(N__44020));
    InMux I__10063 (
            .O(N__44066),
            .I(N__44015));
    InMux I__10062 (
            .O(N__44065),
            .I(N__44015));
    LocalMux I__10061 (
            .O(N__44062),
            .I(N__44007));
    LocalMux I__10060 (
            .O(N__44055),
            .I(N__44007));
    LocalMux I__10059 (
            .O(N__44052),
            .I(N__44007));
    LocalMux I__10058 (
            .O(N__44037),
            .I(N__44004));
    LocalMux I__10057 (
            .O(N__44034),
            .I(N__44001));
    LocalMux I__10056 (
            .O(N__44031),
            .I(N__43998));
    LocalMux I__10055 (
            .O(N__44026),
            .I(N__43993));
    InMux I__10054 (
            .O(N__44025),
            .I(N__43990));
    Span4Mux_v I__10053 (
            .O(N__44020),
            .I(N__43987));
    LocalMux I__10052 (
            .O(N__44015),
            .I(N__43984));
    InMux I__10051 (
            .O(N__44014),
            .I(N__43981));
    Span4Mux_v I__10050 (
            .O(N__44007),
            .I(N__43976));
    Span4Mux_v I__10049 (
            .O(N__44004),
            .I(N__43976));
    Span4Mux_h I__10048 (
            .O(N__44001),
            .I(N__43973));
    Span4Mux_h I__10047 (
            .O(N__43998),
            .I(N__43970));
    InMux I__10046 (
            .O(N__43997),
            .I(N__43967));
    InMux I__10045 (
            .O(N__43996),
            .I(N__43964));
    Span12Mux_h I__10044 (
            .O(N__43993),
            .I(N__43961));
    LocalMux I__10043 (
            .O(N__43990),
            .I(N__43956));
    Span4Mux_h I__10042 (
            .O(N__43987),
            .I(N__43956));
    Span4Mux_h I__10041 (
            .O(N__43984),
            .I(N__43947));
    LocalMux I__10040 (
            .O(N__43981),
            .I(N__43947));
    Span4Mux_h I__10039 (
            .O(N__43976),
            .I(N__43947));
    Span4Mux_h I__10038 (
            .O(N__43973),
            .I(N__43947));
    Span4Mux_h I__10037 (
            .O(N__43970),
            .I(N__43944));
    LocalMux I__10036 (
            .O(N__43967),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__10035 (
            .O(N__43964),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv12 I__10034 (
            .O(N__43961),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__10033 (
            .O(N__43956),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__10032 (
            .O(N__43947),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__10031 (
            .O(N__43944),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    InMux I__10030 (
            .O(N__43931),
            .I(N__43928));
    LocalMux I__10029 (
            .O(N__43928),
            .I(N__43924));
    InMux I__10028 (
            .O(N__43927),
            .I(N__43920));
    Span12Mux_s8_h I__10027 (
            .O(N__43924),
            .I(N__43917));
    InMux I__10026 (
            .O(N__43923),
            .I(N__43914));
    LocalMux I__10025 (
            .O(N__43920),
            .I(\current_shift_inst.un4_control_input1_11 ));
    Odrv12 I__10024 (
            .O(N__43917),
            .I(\current_shift_inst.un4_control_input1_11 ));
    LocalMux I__10023 (
            .O(N__43914),
            .I(\current_shift_inst.un4_control_input1_11 ));
    CascadeMux I__10022 (
            .O(N__43907),
            .I(N__43904));
    InMux I__10021 (
            .O(N__43904),
            .I(N__43901));
    LocalMux I__10020 (
            .O(N__43901),
            .I(N__43898));
    Odrv12 I__10019 (
            .O(N__43898),
            .I(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ));
    InMux I__10018 (
            .O(N__43895),
            .I(N__43892));
    LocalMux I__10017 (
            .O(N__43892),
            .I(N__43889));
    Odrv12 I__10016 (
            .O(N__43889),
            .I(\current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ));
    CascadeMux I__10015 (
            .O(N__43886),
            .I(N__43883));
    InMux I__10014 (
            .O(N__43883),
            .I(N__43879));
    InMux I__10013 (
            .O(N__43882),
            .I(N__43876));
    LocalMux I__10012 (
            .O(N__43879),
            .I(N__43873));
    LocalMux I__10011 (
            .O(N__43876),
            .I(N__43869));
    Span4Mux_v I__10010 (
            .O(N__43873),
            .I(N__43866));
    InMux I__10009 (
            .O(N__43872),
            .I(N__43863));
    Odrv12 I__10008 (
            .O(N__43869),
            .I(\current_shift_inst.un4_control_input1_10 ));
    Odrv4 I__10007 (
            .O(N__43866),
            .I(\current_shift_inst.un4_control_input1_10 ));
    LocalMux I__10006 (
            .O(N__43863),
            .I(\current_shift_inst.un4_control_input1_10 ));
    CascadeMux I__10005 (
            .O(N__43856),
            .I(N__43853));
    InMux I__10004 (
            .O(N__43853),
            .I(N__43850));
    LocalMux I__10003 (
            .O(N__43850),
            .I(N__43847));
    Span4Mux_h I__10002 (
            .O(N__43847),
            .I(N__43844));
    Odrv4 I__10001 (
            .O(N__43844),
            .I(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ));
    InMux I__10000 (
            .O(N__43841),
            .I(N__43838));
    LocalMux I__9999 (
            .O(N__43838),
            .I(\current_shift_inst.un4_control_input_1_axb_2 ));
    CascadeMux I__9998 (
            .O(N__43835),
            .I(N__43832));
    InMux I__9997 (
            .O(N__43832),
            .I(N__43829));
    LocalMux I__9996 (
            .O(N__43829),
            .I(N__43826));
    Span4Mux_v I__9995 (
            .O(N__43826),
            .I(N__43823));
    Span4Mux_h I__9994 (
            .O(N__43823),
            .I(N__43820));
    Odrv4 I__9993 (
            .O(N__43820),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ));
    InMux I__9992 (
            .O(N__43817),
            .I(N__43814));
    LocalMux I__9991 (
            .O(N__43814),
            .I(\current_shift_inst.un4_control_input_1_axb_1 ));
    CascadeMux I__9990 (
            .O(N__43811),
            .I(N__43807));
    InMux I__9989 (
            .O(N__43810),
            .I(N__43802));
    InMux I__9988 (
            .O(N__43807),
            .I(N__43802));
    LocalMux I__9987 (
            .O(N__43802),
            .I(N__43798));
    InMux I__9986 (
            .O(N__43801),
            .I(N__43794));
    Span4Mux_h I__9985 (
            .O(N__43798),
            .I(N__43791));
    InMux I__9984 (
            .O(N__43797),
            .I(N__43788));
    LocalMux I__9983 (
            .O(N__43794),
            .I(N__43785));
    Odrv4 I__9982 (
            .O(N__43791),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    LocalMux I__9981 (
            .O(N__43788),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    Odrv12 I__9980 (
            .O(N__43785),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    CascadeMux I__9979 (
            .O(N__43778),
            .I(N__43775));
    InMux I__9978 (
            .O(N__43775),
            .I(N__43772));
    LocalMux I__9977 (
            .O(N__43772),
            .I(N__43769));
    Span4Mux_v I__9976 (
            .O(N__43769),
            .I(N__43766));
    Odrv4 I__9975 (
            .O(N__43766),
            .I(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ));
    CascadeMux I__9974 (
            .O(N__43763),
            .I(N__43760));
    InMux I__9973 (
            .O(N__43760),
            .I(N__43751));
    InMux I__9972 (
            .O(N__43759),
            .I(N__43751));
    InMux I__9971 (
            .O(N__43758),
            .I(N__43751));
    LocalMux I__9970 (
            .O(N__43751),
            .I(\current_shift_inst.un4_control_input1_2 ));
    InMux I__9969 (
            .O(N__43748),
            .I(N__43736));
    InMux I__9968 (
            .O(N__43747),
            .I(N__43736));
    InMux I__9967 (
            .O(N__43746),
            .I(N__43736));
    InMux I__9966 (
            .O(N__43745),
            .I(N__43736));
    LocalMux I__9965 (
            .O(N__43736),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    CascadeMux I__9964 (
            .O(N__43733),
            .I(N__43730));
    InMux I__9963 (
            .O(N__43730),
            .I(N__43727));
    LocalMux I__9962 (
            .O(N__43727),
            .I(N__43724));
    Span4Mux_h I__9961 (
            .O(N__43724),
            .I(N__43721));
    Odrv4 I__9960 (
            .O(N__43721),
            .I(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ));
    InMux I__9959 (
            .O(N__43718),
            .I(N__43715));
    LocalMux I__9958 (
            .O(N__43715),
            .I(N__43712));
    Odrv4 I__9957 (
            .O(N__43712),
            .I(\current_shift_inst.un4_control_input_1_axb_20 ));
    InMux I__9956 (
            .O(N__43709),
            .I(N__43705));
    CascadeMux I__9955 (
            .O(N__43708),
            .I(N__43702));
    LocalMux I__9954 (
            .O(N__43705),
            .I(N__43698));
    InMux I__9953 (
            .O(N__43702),
            .I(N__43693));
    InMux I__9952 (
            .O(N__43701),
            .I(N__43693));
    Span4Mux_v I__9951 (
            .O(N__43698),
            .I(N__43690));
    LocalMux I__9950 (
            .O(N__43693),
            .I(N__43687));
    Odrv4 I__9949 (
            .O(N__43690),
            .I(\current_shift_inst.un4_control_input1_17 ));
    Odrv4 I__9948 (
            .O(N__43687),
            .I(\current_shift_inst.un4_control_input1_17 ));
    CascadeMux I__9947 (
            .O(N__43682),
            .I(N__43679));
    InMux I__9946 (
            .O(N__43679),
            .I(N__43676));
    LocalMux I__9945 (
            .O(N__43676),
            .I(N__43673));
    Span4Mux_v I__9944 (
            .O(N__43673),
            .I(N__43670));
    Odrv4 I__9943 (
            .O(N__43670),
            .I(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ));
    CascadeMux I__9942 (
            .O(N__43667),
            .I(N__43664));
    InMux I__9941 (
            .O(N__43664),
            .I(N__43660));
    CascadeMux I__9940 (
            .O(N__43663),
            .I(N__43657));
    LocalMux I__9939 (
            .O(N__43660),
            .I(N__43654));
    InMux I__9938 (
            .O(N__43657),
            .I(N__43651));
    Span4Mux_v I__9937 (
            .O(N__43654),
            .I(N__43647));
    LocalMux I__9936 (
            .O(N__43651),
            .I(N__43644));
    InMux I__9935 (
            .O(N__43650),
            .I(N__43641));
    Span4Mux_h I__9934 (
            .O(N__43647),
            .I(N__43638));
    Span4Mux_h I__9933 (
            .O(N__43644),
            .I(N__43635));
    LocalMux I__9932 (
            .O(N__43641),
            .I(N__43632));
    Odrv4 I__9931 (
            .O(N__43638),
            .I(\current_shift_inst.un4_control_input1_18 ));
    Odrv4 I__9930 (
            .O(N__43635),
            .I(\current_shift_inst.un4_control_input1_18 ));
    Odrv4 I__9929 (
            .O(N__43632),
            .I(\current_shift_inst.un4_control_input1_18 ));
    InMux I__9928 (
            .O(N__43625),
            .I(N__43622));
    LocalMux I__9927 (
            .O(N__43622),
            .I(N__43619));
    Span4Mux_v I__9926 (
            .O(N__43619),
            .I(N__43616));
    Odrv4 I__9925 (
            .O(N__43616),
            .I(\current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ));
    InMux I__9924 (
            .O(N__43613),
            .I(N__43608));
    InMux I__9923 (
            .O(N__43612),
            .I(N__43605));
    InMux I__9922 (
            .O(N__43611),
            .I(N__43602));
    LocalMux I__9921 (
            .O(N__43608),
            .I(N__43599));
    LocalMux I__9920 (
            .O(N__43605),
            .I(N__43596));
    LocalMux I__9919 (
            .O(N__43602),
            .I(N__43593));
    Odrv12 I__9918 (
            .O(N__43599),
            .I(\current_shift_inst.un4_control_input1_13 ));
    Odrv4 I__9917 (
            .O(N__43596),
            .I(\current_shift_inst.un4_control_input1_13 ));
    Odrv4 I__9916 (
            .O(N__43593),
            .I(\current_shift_inst.un4_control_input1_13 ));
    CascadeMux I__9915 (
            .O(N__43586),
            .I(N__43583));
    InMux I__9914 (
            .O(N__43583),
            .I(N__43580));
    LocalMux I__9913 (
            .O(N__43580),
            .I(N__43577));
    Span4Mux_v I__9912 (
            .O(N__43577),
            .I(N__43574));
    Span4Mux_h I__9911 (
            .O(N__43574),
            .I(N__43571));
    Odrv4 I__9910 (
            .O(N__43571),
            .I(\current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ));
    CascadeMux I__9909 (
            .O(N__43568),
            .I(N__43565));
    InMux I__9908 (
            .O(N__43565),
            .I(N__43562));
    LocalMux I__9907 (
            .O(N__43562),
            .I(N__43559));
    Span4Mux_v I__9906 (
            .O(N__43559),
            .I(N__43556));
    Odrv4 I__9905 (
            .O(N__43556),
            .I(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ));
    InMux I__9904 (
            .O(N__43553),
            .I(N__43549));
    InMux I__9903 (
            .O(N__43552),
            .I(N__43546));
    LocalMux I__9902 (
            .O(N__43549),
            .I(N__43542));
    LocalMux I__9901 (
            .O(N__43546),
            .I(N__43539));
    InMux I__9900 (
            .O(N__43545),
            .I(N__43536));
    Span4Mux_v I__9899 (
            .O(N__43542),
            .I(N__43533));
    Odrv12 I__9898 (
            .O(N__43539),
            .I(\current_shift_inst.un4_control_input1_15 ));
    LocalMux I__9897 (
            .O(N__43536),
            .I(\current_shift_inst.un4_control_input1_15 ));
    Odrv4 I__9896 (
            .O(N__43533),
            .I(\current_shift_inst.un4_control_input1_15 ));
    CascadeMux I__9895 (
            .O(N__43526),
            .I(N__43523));
    InMux I__9894 (
            .O(N__43523),
            .I(N__43520));
    LocalMux I__9893 (
            .O(N__43520),
            .I(N__43517));
    Span4Mux_h I__9892 (
            .O(N__43517),
            .I(N__43514));
    Span4Mux_v I__9891 (
            .O(N__43514),
            .I(N__43511));
    Odrv4 I__9890 (
            .O(N__43511),
            .I(\current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ));
    CascadeMux I__9889 (
            .O(N__43508),
            .I(N__43505));
    InMux I__9888 (
            .O(N__43505),
            .I(N__43501));
    InMux I__9887 (
            .O(N__43504),
            .I(N__43498));
    LocalMux I__9886 (
            .O(N__43501),
            .I(N__43494));
    LocalMux I__9885 (
            .O(N__43498),
            .I(N__43491));
    InMux I__9884 (
            .O(N__43497),
            .I(N__43488));
    Span4Mux_v I__9883 (
            .O(N__43494),
            .I(N__43483));
    Span4Mux_v I__9882 (
            .O(N__43491),
            .I(N__43483));
    LocalMux I__9881 (
            .O(N__43488),
            .I(N__43480));
    Odrv4 I__9880 (
            .O(N__43483),
            .I(\current_shift_inst.un4_control_input1_16 ));
    Odrv4 I__9879 (
            .O(N__43480),
            .I(\current_shift_inst.un4_control_input1_16 ));
    CascadeMux I__9878 (
            .O(N__43475),
            .I(N__43472));
    InMux I__9877 (
            .O(N__43472),
            .I(N__43469));
    LocalMux I__9876 (
            .O(N__43469),
            .I(N__43466));
    Span4Mux_h I__9875 (
            .O(N__43466),
            .I(N__43463));
    Odrv4 I__9874 (
            .O(N__43463),
            .I(\current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ));
    InMux I__9873 (
            .O(N__43460),
            .I(N__43457));
    LocalMux I__9872 (
            .O(N__43457),
            .I(\current_shift_inst.un4_control_input_1_axb_3 ));
    InMux I__9871 (
            .O(N__43454),
            .I(N__43451));
    LocalMux I__9870 (
            .O(N__43451),
            .I(\current_shift_inst.un4_control_input_1_axb_7 ));
    InMux I__9869 (
            .O(N__43448),
            .I(N__43444));
    InMux I__9868 (
            .O(N__43447),
            .I(N__43441));
    LocalMux I__9867 (
            .O(N__43444),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    LocalMux I__9866 (
            .O(N__43441),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__9865 (
            .O(N__43436),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__9864 (
            .O(N__43433),
            .I(N__43429));
    InMux I__9863 (
            .O(N__43432),
            .I(N__43426));
    LocalMux I__9862 (
            .O(N__43429),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    LocalMux I__9861 (
            .O(N__43426),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__9860 (
            .O(N__43421),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ));
    InMux I__9859 (
            .O(N__43418),
            .I(N__43414));
    InMux I__9858 (
            .O(N__43417),
            .I(N__43411));
    LocalMux I__9857 (
            .O(N__43414),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    LocalMux I__9856 (
            .O(N__43411),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__9855 (
            .O(N__43406),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__9854 (
            .O(N__43403),
            .I(N__43399));
    InMux I__9853 (
            .O(N__43402),
            .I(N__43396));
    LocalMux I__9852 (
            .O(N__43399),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__9851 (
            .O(N__43396),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__9850 (
            .O(N__43391),
            .I(bfn_18_13_0_));
    InMux I__9849 (
            .O(N__43388),
            .I(N__43384));
    InMux I__9848 (
            .O(N__43387),
            .I(N__43381));
    LocalMux I__9847 (
            .O(N__43384),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    LocalMux I__9846 (
            .O(N__43381),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__9845 (
            .O(N__43376),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ));
    CEMux I__9844 (
            .O(N__43373),
            .I(N__43364));
    InMux I__9843 (
            .O(N__43372),
            .I(N__43355));
    InMux I__9842 (
            .O(N__43371),
            .I(N__43355));
    InMux I__9841 (
            .O(N__43370),
            .I(N__43355));
    InMux I__9840 (
            .O(N__43369),
            .I(N__43355));
    CEMux I__9839 (
            .O(N__43368),
            .I(N__43352));
    CEMux I__9838 (
            .O(N__43367),
            .I(N__43348));
    LocalMux I__9837 (
            .O(N__43364),
            .I(N__43345));
    LocalMux I__9836 (
            .O(N__43355),
            .I(N__43340));
    LocalMux I__9835 (
            .O(N__43352),
            .I(N__43340));
    InMux I__9834 (
            .O(N__43351),
            .I(N__43323));
    LocalMux I__9833 (
            .O(N__43348),
            .I(N__43318));
    Span4Mux_h I__9832 (
            .O(N__43345),
            .I(N__43318));
    Span4Mux_v I__9831 (
            .O(N__43340),
            .I(N__43315));
    InMux I__9830 (
            .O(N__43339),
            .I(N__43308));
    InMux I__9829 (
            .O(N__43338),
            .I(N__43308));
    InMux I__9828 (
            .O(N__43337),
            .I(N__43308));
    InMux I__9827 (
            .O(N__43336),
            .I(N__43299));
    InMux I__9826 (
            .O(N__43335),
            .I(N__43299));
    InMux I__9825 (
            .O(N__43334),
            .I(N__43299));
    InMux I__9824 (
            .O(N__43333),
            .I(N__43299));
    InMux I__9823 (
            .O(N__43332),
            .I(N__43296));
    InMux I__9822 (
            .O(N__43331),
            .I(N__43291));
    InMux I__9821 (
            .O(N__43330),
            .I(N__43291));
    InMux I__9820 (
            .O(N__43329),
            .I(N__43282));
    InMux I__9819 (
            .O(N__43328),
            .I(N__43282));
    InMux I__9818 (
            .O(N__43327),
            .I(N__43282));
    InMux I__9817 (
            .O(N__43326),
            .I(N__43282));
    LocalMux I__9816 (
            .O(N__43323),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__9815 (
            .O(N__43318),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__9814 (
            .O(N__43315),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    LocalMux I__9813 (
            .O(N__43308),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    LocalMux I__9812 (
            .O(N__43299),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    LocalMux I__9811 (
            .O(N__43296),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    LocalMux I__9810 (
            .O(N__43291),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    LocalMux I__9809 (
            .O(N__43282),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    InMux I__9808 (
            .O(N__43265),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ));
    InMux I__9807 (
            .O(N__43262),
            .I(N__43258));
    InMux I__9806 (
            .O(N__43261),
            .I(N__43255));
    LocalMux I__9805 (
            .O(N__43258),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    LocalMux I__9804 (
            .O(N__43255),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__9803 (
            .O(N__43250),
            .I(N__43245));
    InMux I__9802 (
            .O(N__43249),
            .I(N__43242));
    InMux I__9801 (
            .O(N__43248),
            .I(N__43239));
    LocalMux I__9800 (
            .O(N__43245),
            .I(\current_shift_inst.un4_control_input1_5 ));
    LocalMux I__9799 (
            .O(N__43242),
            .I(\current_shift_inst.un4_control_input1_5 ));
    LocalMux I__9798 (
            .O(N__43239),
            .I(\current_shift_inst.un4_control_input1_5 ));
    CascadeMux I__9797 (
            .O(N__43232),
            .I(N__43229));
    InMux I__9796 (
            .O(N__43229),
            .I(N__43226));
    LocalMux I__9795 (
            .O(N__43226),
            .I(N__43223));
    Span4Mux_h I__9794 (
            .O(N__43223),
            .I(N__43220));
    Span4Mux_v I__9793 (
            .O(N__43220),
            .I(N__43217));
    Odrv4 I__9792 (
            .O(N__43217),
            .I(\current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ));
    CascadeMux I__9791 (
            .O(N__43214),
            .I(N__43211));
    InMux I__9790 (
            .O(N__43211),
            .I(N__43208));
    LocalMux I__9789 (
            .O(N__43208),
            .I(N__43205));
    Span4Mux_h I__9788 (
            .O(N__43205),
            .I(N__43202));
    Odrv4 I__9787 (
            .O(N__43202),
            .I(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ));
    CascadeMux I__9786 (
            .O(N__43199),
            .I(N__43196));
    InMux I__9785 (
            .O(N__43196),
            .I(N__43193));
    LocalMux I__9784 (
            .O(N__43193),
            .I(N__43190));
    Span4Mux_v I__9783 (
            .O(N__43190),
            .I(N__43187));
    Span4Mux_h I__9782 (
            .O(N__43187),
            .I(N__43184));
    Odrv4 I__9781 (
            .O(N__43184),
            .I(\current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ));
    InMux I__9780 (
            .O(N__43181),
            .I(N__43177));
    InMux I__9779 (
            .O(N__43180),
            .I(N__43174));
    LocalMux I__9778 (
            .O(N__43177),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__9777 (
            .O(N__43174),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__9776 (
            .O(N__43169),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__9775 (
            .O(N__43166),
            .I(N__43162));
    InMux I__9774 (
            .O(N__43165),
            .I(N__43159));
    LocalMux I__9773 (
            .O(N__43162),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__9772 (
            .O(N__43159),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__9771 (
            .O(N__43154),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__9770 (
            .O(N__43151),
            .I(N__43147));
    InMux I__9769 (
            .O(N__43150),
            .I(N__43144));
    LocalMux I__9768 (
            .O(N__43147),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    LocalMux I__9767 (
            .O(N__43144),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__9766 (
            .O(N__43139),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__9765 (
            .O(N__43136),
            .I(N__43132));
    InMux I__9764 (
            .O(N__43135),
            .I(N__43129));
    LocalMux I__9763 (
            .O(N__43132),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    LocalMux I__9762 (
            .O(N__43129),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__9761 (
            .O(N__43124),
            .I(bfn_18_12_0_));
    InMux I__9760 (
            .O(N__43121),
            .I(N__43117));
    InMux I__9759 (
            .O(N__43120),
            .I(N__43114));
    LocalMux I__9758 (
            .O(N__43117),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    LocalMux I__9757 (
            .O(N__43114),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__9756 (
            .O(N__43109),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__9755 (
            .O(N__43106),
            .I(N__43102));
    InMux I__9754 (
            .O(N__43105),
            .I(N__43099));
    LocalMux I__9753 (
            .O(N__43102),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    LocalMux I__9752 (
            .O(N__43099),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__9751 (
            .O(N__43094),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__9750 (
            .O(N__43091),
            .I(N__43087));
    InMux I__9749 (
            .O(N__43090),
            .I(N__43084));
    LocalMux I__9748 (
            .O(N__43087),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    LocalMux I__9747 (
            .O(N__43084),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__9746 (
            .O(N__43079),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__9745 (
            .O(N__43076),
            .I(N__43072));
    InMux I__9744 (
            .O(N__43075),
            .I(N__43069));
    LocalMux I__9743 (
            .O(N__43072),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    LocalMux I__9742 (
            .O(N__43069),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__9741 (
            .O(N__43064),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__9740 (
            .O(N__43061),
            .I(N__43058));
    LocalMux I__9739 (
            .O(N__43058),
            .I(N__43055));
    Span4Mux_v I__9738 (
            .O(N__43055),
            .I(N__43051));
    InMux I__9737 (
            .O(N__43054),
            .I(N__43048));
    Odrv4 I__9736 (
            .O(N__43051),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_CO ));
    LocalMux I__9735 (
            .O(N__43048),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_CO ));
    InMux I__9734 (
            .O(N__43043),
            .I(N__43040));
    LocalMux I__9733 (
            .O(N__43040),
            .I(N__43037));
    Span12Mux_h I__9732 (
            .O(N__43037),
            .I(N__43034));
    Odrv12 I__9731 (
            .O(N__43034),
            .I(\phase_controller_inst1.stoper_tr.running_1_sqmuxa ));
    InMux I__9730 (
            .O(N__43031),
            .I(N__43025));
    InMux I__9729 (
            .O(N__43030),
            .I(N__43025));
    LocalMux I__9728 (
            .O(N__43025),
            .I(N__43017));
    InMux I__9727 (
            .O(N__43024),
            .I(N__43013));
    InMux I__9726 (
            .O(N__43023),
            .I(N__43010));
    InMux I__9725 (
            .O(N__43022),
            .I(N__43005));
    InMux I__9724 (
            .O(N__43021),
            .I(N__43005));
    InMux I__9723 (
            .O(N__43020),
            .I(N__43002));
    Span4Mux_h I__9722 (
            .O(N__43017),
            .I(N__42999));
    InMux I__9721 (
            .O(N__43016),
            .I(N__42996));
    LocalMux I__9720 (
            .O(N__43013),
            .I(N__42989));
    LocalMux I__9719 (
            .O(N__43010),
            .I(N__42989));
    LocalMux I__9718 (
            .O(N__43005),
            .I(N__42989));
    LocalMux I__9717 (
            .O(N__43002),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__9716 (
            .O(N__42999),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__9715 (
            .O(N__42996),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv12 I__9714 (
            .O(N__42989),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    CascadeMux I__9713 (
            .O(N__42980),
            .I(N__42976));
    InMux I__9712 (
            .O(N__42979),
            .I(N__42972));
    InMux I__9711 (
            .O(N__42976),
            .I(N__42968));
    CascadeMux I__9710 (
            .O(N__42975),
            .I(N__42965));
    LocalMux I__9709 (
            .O(N__42972),
            .I(N__42962));
    InMux I__9708 (
            .O(N__42971),
            .I(N__42959));
    LocalMux I__9707 (
            .O(N__42968),
            .I(N__42955));
    InMux I__9706 (
            .O(N__42965),
            .I(N__42952));
    Span4Mux_v I__9705 (
            .O(N__42962),
            .I(N__42949));
    LocalMux I__9704 (
            .O(N__42959),
            .I(N__42946));
    InMux I__9703 (
            .O(N__42958),
            .I(N__42941));
    Span4Mux_h I__9702 (
            .O(N__42955),
            .I(N__42938));
    LocalMux I__9701 (
            .O(N__42952),
            .I(N__42931));
    Span4Mux_h I__9700 (
            .O(N__42949),
            .I(N__42931));
    Span4Mux_v I__9699 (
            .O(N__42946),
            .I(N__42931));
    InMux I__9698 (
            .O(N__42945),
            .I(N__42926));
    InMux I__9697 (
            .O(N__42944),
            .I(N__42926));
    LocalMux I__9696 (
            .O(N__42941),
            .I(N__42923));
    Odrv4 I__9695 (
            .O(N__42938),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    Odrv4 I__9694 (
            .O(N__42931),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    LocalMux I__9693 (
            .O(N__42926),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    Odrv12 I__9692 (
            .O(N__42923),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    CascadeMux I__9691 (
            .O(N__42914),
            .I(\phase_controller_inst1.stoper_tr.running_1_sqmuxa_cascade_ ));
    InMux I__9690 (
            .O(N__42911),
            .I(N__42908));
    LocalMux I__9689 (
            .O(N__42908),
            .I(N__42904));
    InMux I__9688 (
            .O(N__42907),
            .I(N__42901));
    Span4Mux_h I__9687 (
            .O(N__42904),
            .I(N__42897));
    LocalMux I__9686 (
            .O(N__42901),
            .I(N__42894));
    InMux I__9685 (
            .O(N__42900),
            .I(N__42891));
    Span4Mux_h I__9684 (
            .O(N__42897),
            .I(N__42888));
    Span4Mux_h I__9683 (
            .O(N__42894),
            .I(N__42885));
    LocalMux I__9682 (
            .O(N__42891),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    Odrv4 I__9681 (
            .O(N__42888),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    Odrv4 I__9680 (
            .O(N__42885),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    InMux I__9679 (
            .O(N__42878),
            .I(N__42875));
    LocalMux I__9678 (
            .O(N__42875),
            .I(N__42872));
    Span4Mux_h I__9677 (
            .O(N__42872),
            .I(N__42869));
    Odrv4 I__9676 (
            .O(N__42869),
            .I(\phase_controller_inst1.stoper_tr.un1_start_latched2_0 ));
    InMux I__9675 (
            .O(N__42866),
            .I(N__42861));
    InMux I__9674 (
            .O(N__42865),
            .I(N__42858));
    InMux I__9673 (
            .O(N__42864),
            .I(N__42855));
    LocalMux I__9672 (
            .O(N__42861),
            .I(N__42852));
    LocalMux I__9671 (
            .O(N__42858),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    LocalMux I__9670 (
            .O(N__42855),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    Odrv4 I__9669 (
            .O(N__42852),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    InMux I__9668 (
            .O(N__42845),
            .I(N__42841));
    InMux I__9667 (
            .O(N__42844),
            .I(N__42836));
    LocalMux I__9666 (
            .O(N__42841),
            .I(N__42833));
    InMux I__9665 (
            .O(N__42840),
            .I(N__42830));
    InMux I__9664 (
            .O(N__42839),
            .I(N__42827));
    LocalMux I__9663 (
            .O(N__42836),
            .I(N__42824));
    Span4Mux_v I__9662 (
            .O(N__42833),
            .I(N__42821));
    LocalMux I__9661 (
            .O(N__42830),
            .I(N__42816));
    LocalMux I__9660 (
            .O(N__42827),
            .I(N__42816));
    Span4Mux_h I__9659 (
            .O(N__42824),
            .I(N__42813));
    Odrv4 I__9658 (
            .O(N__42821),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    Odrv12 I__9657 (
            .O(N__42816),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    Odrv4 I__9656 (
            .O(N__42813),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    InMux I__9655 (
            .O(N__42806),
            .I(N__42803));
    LocalMux I__9654 (
            .O(N__42803),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ));
    CascadeMux I__9653 (
            .O(N__42800),
            .I(N__42797));
    InMux I__9652 (
            .O(N__42797),
            .I(N__42792));
    InMux I__9651 (
            .O(N__42796),
            .I(N__42789));
    CascadeMux I__9650 (
            .O(N__42795),
            .I(N__42786));
    LocalMux I__9649 (
            .O(N__42792),
            .I(N__42783));
    LocalMux I__9648 (
            .O(N__42789),
            .I(N__42780));
    InMux I__9647 (
            .O(N__42786),
            .I(N__42777));
    Span4Mux_h I__9646 (
            .O(N__42783),
            .I(N__42774));
    Span4Mux_v I__9645 (
            .O(N__42780),
            .I(N__42771));
    LocalMux I__9644 (
            .O(N__42777),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__9643 (
            .O(N__42774),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__9642 (
            .O(N__42771),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__9641 (
            .O(N__42764),
            .I(N__42760));
    InMux I__9640 (
            .O(N__42763),
            .I(N__42757));
    LocalMux I__9639 (
            .O(N__42760),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__9638 (
            .O(N__42757),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__9637 (
            .O(N__42752),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ));
    InMux I__9636 (
            .O(N__42749),
            .I(N__42746));
    LocalMux I__9635 (
            .O(N__42746),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNISF8IZ0Z2 ));
    CascadeMux I__9634 (
            .O(N__42743),
            .I(N__42740));
    InMux I__9633 (
            .O(N__42740),
            .I(N__42736));
    InMux I__9632 (
            .O(N__42739),
            .I(N__42733));
    LocalMux I__9631 (
            .O(N__42736),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__9630 (
            .O(N__42733),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__9629 (
            .O(N__42728),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__9628 (
            .O(N__42725),
            .I(N__42721));
    InMux I__9627 (
            .O(N__42724),
            .I(N__42718));
    LocalMux I__9626 (
            .O(N__42721),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__9625 (
            .O(N__42718),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__9624 (
            .O(N__42713),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__9623 (
            .O(N__42710),
            .I(N__42706));
    InMux I__9622 (
            .O(N__42709),
            .I(N__42703));
    LocalMux I__9621 (
            .O(N__42706),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__9620 (
            .O(N__42703),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__9619 (
            .O(N__42698),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ));
    InMux I__9618 (
            .O(N__42695),
            .I(N__42692));
    LocalMux I__9617 (
            .O(N__42692),
            .I(N__42687));
    InMux I__9616 (
            .O(N__42691),
            .I(N__42684));
    InMux I__9615 (
            .O(N__42690),
            .I(N__42681));
    Span4Mux_h I__9614 (
            .O(N__42687),
            .I(N__42678));
    LocalMux I__9613 (
            .O(N__42684),
            .I(elapsed_time_ns_1_RNIUKL2M1_0_6));
    LocalMux I__9612 (
            .O(N__42681),
            .I(elapsed_time_ns_1_RNIUKL2M1_0_6));
    Odrv4 I__9611 (
            .O(N__42678),
            .I(elapsed_time_ns_1_RNIUKL2M1_0_6));
    CascadeMux I__9610 (
            .O(N__42671),
            .I(N__42668));
    InMux I__9609 (
            .O(N__42668),
            .I(N__42665));
    LocalMux I__9608 (
            .O(N__42665),
            .I(\phase_controller_inst1.stoper_tr.un6_running_6 ));
    InMux I__9607 (
            .O(N__42662),
            .I(N__42658));
    InMux I__9606 (
            .O(N__42661),
            .I(N__42655));
    LocalMux I__9605 (
            .O(N__42658),
            .I(N__42652));
    LocalMux I__9604 (
            .O(N__42655),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2 ));
    Odrv12 I__9603 (
            .O(N__42652),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2 ));
    InMux I__9602 (
            .O(N__42647),
            .I(N__42644));
    LocalMux I__9601 (
            .O(N__42644),
            .I(\phase_controller_inst1.stoper_tr.un6_running_2 ));
    InMux I__9600 (
            .O(N__42641),
            .I(N__42638));
    LocalMux I__9599 (
            .O(N__42638),
            .I(\phase_controller_inst1.stoper_tr.un6_running_4 ));
    CascadeMux I__9598 (
            .O(N__42635),
            .I(N__42632));
    InMux I__9597 (
            .O(N__42632),
            .I(N__42629));
    LocalMux I__9596 (
            .O(N__42629),
            .I(\phase_controller_inst1.stoper_tr.un6_running_5 ));
    CascadeMux I__9595 (
            .O(N__42626),
            .I(N__42622));
    InMux I__9594 (
            .O(N__42625),
            .I(N__42618));
    InMux I__9593 (
            .O(N__42622),
            .I(N__42615));
    InMux I__9592 (
            .O(N__42621),
            .I(N__42611));
    LocalMux I__9591 (
            .O(N__42618),
            .I(N__42608));
    LocalMux I__9590 (
            .O(N__42615),
            .I(N__42605));
    InMux I__9589 (
            .O(N__42614),
            .I(N__42602));
    LocalMux I__9588 (
            .O(N__42611),
            .I(elapsed_time_ns_1_RNIFJ2591_0_7));
    Odrv12 I__9587 (
            .O(N__42608),
            .I(elapsed_time_ns_1_RNIFJ2591_0_7));
    Odrv4 I__9586 (
            .O(N__42605),
            .I(elapsed_time_ns_1_RNIFJ2591_0_7));
    LocalMux I__9585 (
            .O(N__42602),
            .I(elapsed_time_ns_1_RNIFJ2591_0_7));
    InMux I__9584 (
            .O(N__42593),
            .I(N__42590));
    LocalMux I__9583 (
            .O(N__42590),
            .I(\phase_controller_inst1.stoper_tr.un6_running_7 ));
    CascadeMux I__9582 (
            .O(N__42587),
            .I(N__42583));
    CascadeMux I__9581 (
            .O(N__42586),
            .I(N__42580));
    InMux I__9580 (
            .O(N__42583),
            .I(N__42577));
    InMux I__9579 (
            .O(N__42580),
            .I(N__42574));
    LocalMux I__9578 (
            .O(N__42577),
            .I(N__42571));
    LocalMux I__9577 (
            .O(N__42574),
            .I(N__42568));
    Span4Mux_h I__9576 (
            .O(N__42571),
            .I(N__42564));
    Span4Mux_h I__9575 (
            .O(N__42568),
            .I(N__42561));
    InMux I__9574 (
            .O(N__42567),
            .I(N__42558));
    Odrv4 I__9573 (
            .O(N__42564),
            .I(elapsed_time_ns_1_RNICG2591_0_4));
    Odrv4 I__9572 (
            .O(N__42561),
            .I(elapsed_time_ns_1_RNICG2591_0_4));
    LocalMux I__9571 (
            .O(N__42558),
            .I(elapsed_time_ns_1_RNICG2591_0_4));
    CascadeMux I__9570 (
            .O(N__42551),
            .I(N__42548));
    InMux I__9569 (
            .O(N__42548),
            .I(N__42545));
    LocalMux I__9568 (
            .O(N__42545),
            .I(N__42542));
    Span4Mux_h I__9567 (
            .O(N__42542),
            .I(N__42539));
    Odrv4 I__9566 (
            .O(N__42539),
            .I(\phase_controller_inst2.stoper_tr.un6_running_4 ));
    InMux I__9565 (
            .O(N__42536),
            .I(N__42499));
    InMux I__9564 (
            .O(N__42535),
            .I(N__42499));
    InMux I__9563 (
            .O(N__42534),
            .I(N__42499));
    InMux I__9562 (
            .O(N__42533),
            .I(N__42499));
    InMux I__9561 (
            .O(N__42532),
            .I(N__42499));
    InMux I__9560 (
            .O(N__42531),
            .I(N__42494));
    InMux I__9559 (
            .O(N__42530),
            .I(N__42494));
    InMux I__9558 (
            .O(N__42529),
            .I(N__42479));
    InMux I__9557 (
            .O(N__42528),
            .I(N__42479));
    InMux I__9556 (
            .O(N__42527),
            .I(N__42479));
    InMux I__9555 (
            .O(N__42526),
            .I(N__42479));
    InMux I__9554 (
            .O(N__42525),
            .I(N__42479));
    InMux I__9553 (
            .O(N__42524),
            .I(N__42479));
    InMux I__9552 (
            .O(N__42523),
            .I(N__42479));
    InMux I__9551 (
            .O(N__42522),
            .I(N__42468));
    InMux I__9550 (
            .O(N__42521),
            .I(N__42468));
    InMux I__9549 (
            .O(N__42520),
            .I(N__42468));
    InMux I__9548 (
            .O(N__42519),
            .I(N__42468));
    InMux I__9547 (
            .O(N__42518),
            .I(N__42468));
    InMux I__9546 (
            .O(N__42517),
            .I(N__42454));
    InMux I__9545 (
            .O(N__42516),
            .I(N__42454));
    InMux I__9544 (
            .O(N__42515),
            .I(N__42454));
    InMux I__9543 (
            .O(N__42514),
            .I(N__42454));
    InMux I__9542 (
            .O(N__42513),
            .I(N__42454));
    InMux I__9541 (
            .O(N__42512),
            .I(N__42454));
    InMux I__9540 (
            .O(N__42511),
            .I(N__42445));
    InMux I__9539 (
            .O(N__42510),
            .I(N__42445));
    LocalMux I__9538 (
            .O(N__42499),
            .I(N__42442));
    LocalMux I__9537 (
            .O(N__42494),
            .I(N__42439));
    LocalMux I__9536 (
            .O(N__42479),
            .I(N__42434));
    LocalMux I__9535 (
            .O(N__42468),
            .I(N__42434));
    InMux I__9534 (
            .O(N__42467),
            .I(N__42428));
    LocalMux I__9533 (
            .O(N__42454),
            .I(N__42425));
    InMux I__9532 (
            .O(N__42453),
            .I(N__42422));
    InMux I__9531 (
            .O(N__42452),
            .I(N__42419));
    InMux I__9530 (
            .O(N__42451),
            .I(N__42414));
    InMux I__9529 (
            .O(N__42450),
            .I(N__42414));
    LocalMux I__9528 (
            .O(N__42445),
            .I(N__42409));
    Span4Mux_h I__9527 (
            .O(N__42442),
            .I(N__42409));
    Span4Mux_h I__9526 (
            .O(N__42439),
            .I(N__42404));
    Span4Mux_v I__9525 (
            .O(N__42434),
            .I(N__42404));
    InMux I__9524 (
            .O(N__42433),
            .I(N__42397));
    InMux I__9523 (
            .O(N__42432),
            .I(N__42397));
    InMux I__9522 (
            .O(N__42431),
            .I(N__42397));
    LocalMux I__9521 (
            .O(N__42428),
            .I(N__42388));
    Span4Mux_v I__9520 (
            .O(N__42425),
            .I(N__42388));
    LocalMux I__9519 (
            .O(N__42422),
            .I(N__42388));
    LocalMux I__9518 (
            .O(N__42419),
            .I(N__42388));
    LocalMux I__9517 (
            .O(N__42414),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    Odrv4 I__9516 (
            .O(N__42409),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    Odrv4 I__9515 (
            .O(N__42404),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    LocalMux I__9514 (
            .O(N__42397),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    Odrv4 I__9513 (
            .O(N__42388),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    InMux I__9512 (
            .O(N__42377),
            .I(N__42374));
    LocalMux I__9511 (
            .O(N__42374),
            .I(N__42370));
    InMux I__9510 (
            .O(N__42373),
            .I(N__42367));
    Span4Mux_v I__9509 (
            .O(N__42370),
            .I(N__42361));
    LocalMux I__9508 (
            .O(N__42367),
            .I(N__42361));
    InMux I__9507 (
            .O(N__42366),
            .I(N__42357));
    Span4Mux_h I__9506 (
            .O(N__42361),
            .I(N__42354));
    InMux I__9505 (
            .O(N__42360),
            .I(N__42351));
    LocalMux I__9504 (
            .O(N__42357),
            .I(elapsed_time_ns_1_RNIDH2591_0_5));
    Odrv4 I__9503 (
            .O(N__42354),
            .I(elapsed_time_ns_1_RNIDH2591_0_5));
    LocalMux I__9502 (
            .O(N__42351),
            .I(elapsed_time_ns_1_RNIDH2591_0_5));
    InMux I__9501 (
            .O(N__42344),
            .I(N__42341));
    LocalMux I__9500 (
            .O(N__42341),
            .I(N__42338));
    Span4Mux_h I__9499 (
            .O(N__42338),
            .I(N__42335));
    Odrv4 I__9498 (
            .O(N__42335),
            .I(\phase_controller_inst2.stoper_tr.un6_running_5 ));
    CascadeMux I__9497 (
            .O(N__42332),
            .I(N__42328));
    InMux I__9496 (
            .O(N__42331),
            .I(N__42325));
    InMux I__9495 (
            .O(N__42328),
            .I(N__42322));
    LocalMux I__9494 (
            .O(N__42325),
            .I(N__42319));
    LocalMux I__9493 (
            .O(N__42322),
            .I(N__42316));
    Span4Mux_h I__9492 (
            .O(N__42319),
            .I(N__42313));
    Odrv12 I__9491 (
            .O(N__42316),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3 ));
    Odrv4 I__9490 (
            .O(N__42313),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3 ));
    CascadeMux I__9489 (
            .O(N__42308),
            .I(N__42300));
    CascadeMux I__9488 (
            .O(N__42307),
            .I(N__42297));
    InMux I__9487 (
            .O(N__42306),
            .I(N__42282));
    InMux I__9486 (
            .O(N__42305),
            .I(N__42282));
    InMux I__9485 (
            .O(N__42304),
            .I(N__42282));
    InMux I__9484 (
            .O(N__42303),
            .I(N__42279));
    InMux I__9483 (
            .O(N__42300),
            .I(N__42268));
    InMux I__9482 (
            .O(N__42297),
            .I(N__42268));
    InMux I__9481 (
            .O(N__42296),
            .I(N__42268));
    InMux I__9480 (
            .O(N__42295),
            .I(N__42268));
    InMux I__9479 (
            .O(N__42294),
            .I(N__42268));
    InMux I__9478 (
            .O(N__42293),
            .I(N__42261));
    InMux I__9477 (
            .O(N__42292),
            .I(N__42261));
    InMux I__9476 (
            .O(N__42291),
            .I(N__42261));
    InMux I__9475 (
            .O(N__42290),
            .I(N__42256));
    InMux I__9474 (
            .O(N__42289),
            .I(N__42256));
    LocalMux I__9473 (
            .O(N__42282),
            .I(N__42253));
    LocalMux I__9472 (
            .O(N__42279),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_0_6 ));
    LocalMux I__9471 (
            .O(N__42268),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_0_6 ));
    LocalMux I__9470 (
            .O(N__42261),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_0_6 ));
    LocalMux I__9469 (
            .O(N__42256),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_0_6 ));
    Odrv4 I__9468 (
            .O(N__42253),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_0_6 ));
    CascadeMux I__9467 (
            .O(N__42242),
            .I(N__42236));
    CascadeMux I__9466 (
            .O(N__42241),
            .I(N__42233));
    CascadeMux I__9465 (
            .O(N__42240),
            .I(N__42228));
    CascadeMux I__9464 (
            .O(N__42239),
            .I(N__42225));
    InMux I__9463 (
            .O(N__42236),
            .I(N__42217));
    InMux I__9462 (
            .O(N__42233),
            .I(N__42212));
    InMux I__9461 (
            .O(N__42232),
            .I(N__42212));
    InMux I__9460 (
            .O(N__42231),
            .I(N__42209));
    InMux I__9459 (
            .O(N__42228),
            .I(N__42206));
    InMux I__9458 (
            .O(N__42225),
            .I(N__42203));
    InMux I__9457 (
            .O(N__42224),
            .I(N__42200));
    InMux I__9456 (
            .O(N__42223),
            .I(N__42191));
    InMux I__9455 (
            .O(N__42222),
            .I(N__42191));
    InMux I__9454 (
            .O(N__42221),
            .I(N__42191));
    InMux I__9453 (
            .O(N__42220),
            .I(N__42191));
    LocalMux I__9452 (
            .O(N__42217),
            .I(N__42186));
    LocalMux I__9451 (
            .O(N__42212),
            .I(N__42186));
    LocalMux I__9450 (
            .O(N__42209),
            .I(N__42183));
    LocalMux I__9449 (
            .O(N__42206),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ));
    LocalMux I__9448 (
            .O(N__42203),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ));
    LocalMux I__9447 (
            .O(N__42200),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ));
    LocalMux I__9446 (
            .O(N__42191),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ));
    Odrv4 I__9445 (
            .O(N__42186),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ));
    Odrv4 I__9444 (
            .O(N__42183),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ));
    InMux I__9443 (
            .O(N__42170),
            .I(N__42166));
    InMux I__9442 (
            .O(N__42169),
            .I(N__42161));
    LocalMux I__9441 (
            .O(N__42166),
            .I(N__42158));
    CascadeMux I__9440 (
            .O(N__42165),
            .I(N__42155));
    InMux I__9439 (
            .O(N__42164),
            .I(N__42151));
    LocalMux I__9438 (
            .O(N__42161),
            .I(N__42148));
    Span4Mux_v I__9437 (
            .O(N__42158),
            .I(N__42145));
    InMux I__9436 (
            .O(N__42155),
            .I(N__42142));
    InMux I__9435 (
            .O(N__42154),
            .I(N__42139));
    LocalMux I__9434 (
            .O(N__42151),
            .I(elapsed_time_ns_1_RNIRHL2M1_0_3));
    Odrv12 I__9433 (
            .O(N__42148),
            .I(elapsed_time_ns_1_RNIRHL2M1_0_3));
    Odrv4 I__9432 (
            .O(N__42145),
            .I(elapsed_time_ns_1_RNIRHL2M1_0_3));
    LocalMux I__9431 (
            .O(N__42142),
            .I(elapsed_time_ns_1_RNIRHL2M1_0_3));
    LocalMux I__9430 (
            .O(N__42139),
            .I(elapsed_time_ns_1_RNIRHL2M1_0_3));
    InMux I__9429 (
            .O(N__42128),
            .I(N__42125));
    LocalMux I__9428 (
            .O(N__42125),
            .I(N__42122));
    Odrv4 I__9427 (
            .O(N__42122),
            .I(\phase_controller_inst2.stoper_tr.un6_running_3 ));
    CEMux I__9426 (
            .O(N__42119),
            .I(N__42112));
    CEMux I__9425 (
            .O(N__42118),
            .I(N__42109));
    CEMux I__9424 (
            .O(N__42117),
            .I(N__42106));
    CEMux I__9423 (
            .O(N__42116),
            .I(N__42103));
    CEMux I__9422 (
            .O(N__42115),
            .I(N__42099));
    LocalMux I__9421 (
            .O(N__42112),
            .I(N__42084));
    LocalMux I__9420 (
            .O(N__42109),
            .I(N__42076));
    LocalMux I__9419 (
            .O(N__42106),
            .I(N__42076));
    LocalMux I__9418 (
            .O(N__42103),
            .I(N__42073));
    InMux I__9417 (
            .O(N__42102),
            .I(N__42066));
    LocalMux I__9416 (
            .O(N__42099),
            .I(N__42063));
    CEMux I__9415 (
            .O(N__42098),
            .I(N__42060));
    InMux I__9414 (
            .O(N__42097),
            .I(N__42051));
    InMux I__9413 (
            .O(N__42096),
            .I(N__42051));
    InMux I__9412 (
            .O(N__42095),
            .I(N__42051));
    InMux I__9411 (
            .O(N__42094),
            .I(N__42051));
    InMux I__9410 (
            .O(N__42093),
            .I(N__42048));
    InMux I__9409 (
            .O(N__42092),
            .I(N__42039));
    InMux I__9408 (
            .O(N__42091),
            .I(N__42039));
    InMux I__9407 (
            .O(N__42090),
            .I(N__42039));
    InMux I__9406 (
            .O(N__42089),
            .I(N__42039));
    InMux I__9405 (
            .O(N__42088),
            .I(N__42034));
    InMux I__9404 (
            .O(N__42087),
            .I(N__42034));
    Span4Mux_v I__9403 (
            .O(N__42084),
            .I(N__42031));
    InMux I__9402 (
            .O(N__42083),
            .I(N__42024));
    InMux I__9401 (
            .O(N__42082),
            .I(N__42024));
    InMux I__9400 (
            .O(N__42081),
            .I(N__42024));
    Span4Mux_v I__9399 (
            .O(N__42076),
            .I(N__42019));
    Span4Mux_v I__9398 (
            .O(N__42073),
            .I(N__42019));
    InMux I__9397 (
            .O(N__42072),
            .I(N__42010));
    InMux I__9396 (
            .O(N__42071),
            .I(N__42010));
    InMux I__9395 (
            .O(N__42070),
            .I(N__42010));
    InMux I__9394 (
            .O(N__42069),
            .I(N__42010));
    LocalMux I__9393 (
            .O(N__42066),
            .I(N__42007));
    Span4Mux_v I__9392 (
            .O(N__42063),
            .I(N__42004));
    LocalMux I__9391 (
            .O(N__42060),
            .I(N__42001));
    LocalMux I__9390 (
            .O(N__42051),
            .I(N__41994));
    LocalMux I__9389 (
            .O(N__42048),
            .I(N__41994));
    LocalMux I__9388 (
            .O(N__42039),
            .I(N__41994));
    LocalMux I__9387 (
            .O(N__42034),
            .I(N__41991));
    Span4Mux_h I__9386 (
            .O(N__42031),
            .I(N__41982));
    LocalMux I__9385 (
            .O(N__42024),
            .I(N__41982));
    Span4Mux_v I__9384 (
            .O(N__42019),
            .I(N__41982));
    LocalMux I__9383 (
            .O(N__42010),
            .I(N__41982));
    Span4Mux_v I__9382 (
            .O(N__42007),
            .I(N__41979));
    Span4Mux_v I__9381 (
            .O(N__42004),
            .I(N__41976));
    Span12Mux_h I__9380 (
            .O(N__42001),
            .I(N__41973));
    Span4Mux_v I__9379 (
            .O(N__41994),
            .I(N__41968));
    Span4Mux_v I__9378 (
            .O(N__41991),
            .I(N__41968));
    Span4Mux_h I__9377 (
            .O(N__41982),
            .I(N__41965));
    Sp12to4 I__9376 (
            .O(N__41979),
            .I(N__41960));
    Sp12to4 I__9375 (
            .O(N__41976),
            .I(N__41960));
    Odrv12 I__9374 (
            .O(N__41973),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv4 I__9373 (
            .O(N__41968),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv4 I__9372 (
            .O(N__41965),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv12 I__9371 (
            .O(N__41960),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    InMux I__9370 (
            .O(N__41951),
            .I(N__41948));
    LocalMux I__9369 (
            .O(N__41948),
            .I(N__41945));
    Odrv4 I__9368 (
            .O(N__41945),
            .I(\current_shift_inst.un4_control_input_1_axb_25 ));
    InMux I__9367 (
            .O(N__41942),
            .I(N__41939));
    LocalMux I__9366 (
            .O(N__41939),
            .I(N__41936));
    Odrv12 I__9365 (
            .O(N__41936),
            .I(\current_shift_inst.un4_control_input_1_axb_23 ));
    InMux I__9364 (
            .O(N__41933),
            .I(N__41930));
    LocalMux I__9363 (
            .O(N__41930),
            .I(N__41927));
    Odrv12 I__9362 (
            .O(N__41927),
            .I(\current_shift_inst.un4_control_input_1_axb_28 ));
    InMux I__9361 (
            .O(N__41924),
            .I(N__41921));
    LocalMux I__9360 (
            .O(N__41921),
            .I(N__41918));
    Odrv12 I__9359 (
            .O(N__41918),
            .I(\current_shift_inst.un4_control_input_1_axb_29 ));
    InMux I__9358 (
            .O(N__41915),
            .I(N__41912));
    LocalMux I__9357 (
            .O(N__41912),
            .I(N__41909));
    Odrv12 I__9356 (
            .O(N__41909),
            .I(\current_shift_inst.un4_control_input_1_axb_27 ));
    CascadeMux I__9355 (
            .O(N__41906),
            .I(N__41903));
    InMux I__9354 (
            .O(N__41903),
            .I(N__41900));
    LocalMux I__9353 (
            .O(N__41900),
            .I(N__41897));
    Span4Mux_v I__9352 (
            .O(N__41897),
            .I(N__41893));
    InMux I__9351 (
            .O(N__41896),
            .I(N__41890));
    Odrv4 I__9350 (
            .O(N__41893),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    LocalMux I__9349 (
            .O(N__41890),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    InMux I__9348 (
            .O(N__41885),
            .I(N__41882));
    LocalMux I__9347 (
            .O(N__41882),
            .I(N__41879));
    Span4Mux_v I__9346 (
            .O(N__41879),
            .I(N__41874));
    InMux I__9345 (
            .O(N__41878),
            .I(N__41869));
    InMux I__9344 (
            .O(N__41877),
            .I(N__41869));
    Span4Mux_h I__9343 (
            .O(N__41874),
            .I(N__41864));
    LocalMux I__9342 (
            .O(N__41869),
            .I(N__41864));
    Odrv4 I__9341 (
            .O(N__41864),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    InMux I__9340 (
            .O(N__41861),
            .I(N__41857));
    InMux I__9339 (
            .O(N__41860),
            .I(N__41853));
    LocalMux I__9338 (
            .O(N__41857),
            .I(N__41850));
    InMux I__9337 (
            .O(N__41856),
            .I(N__41847));
    LocalMux I__9336 (
            .O(N__41853),
            .I(N__41842));
    Span4Mux_v I__9335 (
            .O(N__41850),
            .I(N__41837));
    LocalMux I__9334 (
            .O(N__41847),
            .I(N__41837));
    InMux I__9333 (
            .O(N__41846),
            .I(N__41832));
    InMux I__9332 (
            .O(N__41845),
            .I(N__41832));
    Odrv4 I__9331 (
            .O(N__41842),
            .I(elapsed_time_ns_1_RNIFG4DM1_0_16));
    Odrv4 I__9330 (
            .O(N__41837),
            .I(elapsed_time_ns_1_RNIFG4DM1_0_16));
    LocalMux I__9329 (
            .O(N__41832),
            .I(elapsed_time_ns_1_RNIFG4DM1_0_16));
    CascadeMux I__9328 (
            .O(N__41825),
            .I(N__41817));
    CascadeMux I__9327 (
            .O(N__41824),
            .I(N__41812));
    CascadeMux I__9326 (
            .O(N__41823),
            .I(N__41806));
    CascadeMux I__9325 (
            .O(N__41822),
            .I(N__41800));
    CascadeMux I__9324 (
            .O(N__41821),
            .I(N__41797));
    InMux I__9323 (
            .O(N__41820),
            .I(N__41793));
    InMux I__9322 (
            .O(N__41817),
            .I(N__41790));
    CascadeMux I__9321 (
            .O(N__41816),
            .I(N__41787));
    CascadeMux I__9320 (
            .O(N__41815),
            .I(N__41783));
    InMux I__9319 (
            .O(N__41812),
            .I(N__41780));
    CascadeMux I__9318 (
            .O(N__41811),
            .I(N__41777));
    CascadeMux I__9317 (
            .O(N__41810),
            .I(N__41774));
    InMux I__9316 (
            .O(N__41809),
            .I(N__41771));
    InMux I__9315 (
            .O(N__41806),
            .I(N__41765));
    InMux I__9314 (
            .O(N__41805),
            .I(N__41762));
    InMux I__9313 (
            .O(N__41804),
            .I(N__41755));
    InMux I__9312 (
            .O(N__41803),
            .I(N__41755));
    InMux I__9311 (
            .O(N__41800),
            .I(N__41755));
    InMux I__9310 (
            .O(N__41797),
            .I(N__41747));
    CascadeMux I__9309 (
            .O(N__41796),
            .I(N__41744));
    LocalMux I__9308 (
            .O(N__41793),
            .I(N__41738));
    LocalMux I__9307 (
            .O(N__41790),
            .I(N__41738));
    InMux I__9306 (
            .O(N__41787),
            .I(N__41731));
    InMux I__9305 (
            .O(N__41786),
            .I(N__41731));
    InMux I__9304 (
            .O(N__41783),
            .I(N__41731));
    LocalMux I__9303 (
            .O(N__41780),
            .I(N__41728));
    InMux I__9302 (
            .O(N__41777),
            .I(N__41725));
    InMux I__9301 (
            .O(N__41774),
            .I(N__41722));
    LocalMux I__9300 (
            .O(N__41771),
            .I(N__41718));
    CascadeMux I__9299 (
            .O(N__41770),
            .I(N__41715));
    CascadeMux I__9298 (
            .O(N__41769),
            .I(N__41712));
    CascadeMux I__9297 (
            .O(N__41768),
            .I(N__41709));
    LocalMux I__9296 (
            .O(N__41765),
            .I(N__41706));
    LocalMux I__9295 (
            .O(N__41762),
            .I(N__41701));
    LocalMux I__9294 (
            .O(N__41755),
            .I(N__41701));
    CascadeMux I__9293 (
            .O(N__41754),
            .I(N__41697));
    CascadeMux I__9292 (
            .O(N__41753),
            .I(N__41694));
    CascadeMux I__9291 (
            .O(N__41752),
            .I(N__41691));
    CascadeMux I__9290 (
            .O(N__41751),
            .I(N__41686));
    CascadeMux I__9289 (
            .O(N__41750),
            .I(N__41682));
    LocalMux I__9288 (
            .O(N__41747),
            .I(N__41679));
    InMux I__9287 (
            .O(N__41744),
            .I(N__41674));
    InMux I__9286 (
            .O(N__41743),
            .I(N__41674));
    Span4Mux_v I__9285 (
            .O(N__41738),
            .I(N__41669));
    LocalMux I__9284 (
            .O(N__41731),
            .I(N__41669));
    Span4Mux_v I__9283 (
            .O(N__41728),
            .I(N__41662));
    LocalMux I__9282 (
            .O(N__41725),
            .I(N__41662));
    LocalMux I__9281 (
            .O(N__41722),
            .I(N__41662));
    InMux I__9280 (
            .O(N__41721),
            .I(N__41659));
    Span4Mux_v I__9279 (
            .O(N__41718),
            .I(N__41656));
    InMux I__9278 (
            .O(N__41715),
            .I(N__41653));
    InMux I__9277 (
            .O(N__41712),
            .I(N__41650));
    InMux I__9276 (
            .O(N__41709),
            .I(N__41647));
    Span4Mux_h I__9275 (
            .O(N__41706),
            .I(N__41642));
    Span4Mux_h I__9274 (
            .O(N__41701),
            .I(N__41642));
    InMux I__9273 (
            .O(N__41700),
            .I(N__41635));
    InMux I__9272 (
            .O(N__41697),
            .I(N__41635));
    InMux I__9271 (
            .O(N__41694),
            .I(N__41635));
    InMux I__9270 (
            .O(N__41691),
            .I(N__41622));
    InMux I__9269 (
            .O(N__41690),
            .I(N__41622));
    InMux I__9268 (
            .O(N__41689),
            .I(N__41622));
    InMux I__9267 (
            .O(N__41686),
            .I(N__41622));
    InMux I__9266 (
            .O(N__41685),
            .I(N__41622));
    InMux I__9265 (
            .O(N__41682),
            .I(N__41622));
    Span4Mux_v I__9264 (
            .O(N__41679),
            .I(N__41617));
    LocalMux I__9263 (
            .O(N__41674),
            .I(N__41617));
    Span4Mux_h I__9262 (
            .O(N__41669),
            .I(N__41612));
    Span4Mux_h I__9261 (
            .O(N__41662),
            .I(N__41612));
    LocalMux I__9260 (
            .O(N__41659),
            .I(N__41609));
    Odrv4 I__9259 (
            .O(N__41656),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__9258 (
            .O(N__41653),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__9257 (
            .O(N__41650),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__9256 (
            .O(N__41647),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    Odrv4 I__9255 (
            .O(N__41642),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__9254 (
            .O(N__41635),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__9253 (
            .O(N__41622),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    Odrv4 I__9252 (
            .O(N__41617),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    Odrv4 I__9251 (
            .O(N__41612),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    Odrv12 I__9250 (
            .O(N__41609),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    InMux I__9249 (
            .O(N__41588),
            .I(N__41579));
    InMux I__9248 (
            .O(N__41587),
            .I(N__41576));
    InMux I__9247 (
            .O(N__41586),
            .I(N__41573));
    InMux I__9246 (
            .O(N__41585),
            .I(N__41570));
    InMux I__9245 (
            .O(N__41584),
            .I(N__41565));
    InMux I__9244 (
            .O(N__41583),
            .I(N__41565));
    InMux I__9243 (
            .O(N__41582),
            .I(N__41562));
    LocalMux I__9242 (
            .O(N__41579),
            .I(N__41556));
    LocalMux I__9241 (
            .O(N__41576),
            .I(N__41556));
    LocalMux I__9240 (
            .O(N__41573),
            .I(N__41552));
    LocalMux I__9239 (
            .O(N__41570),
            .I(N__41547));
    LocalMux I__9238 (
            .O(N__41565),
            .I(N__41547));
    LocalMux I__9237 (
            .O(N__41562),
            .I(N__41544));
    InMux I__9236 (
            .O(N__41561),
            .I(N__41541));
    Span4Mux_v I__9235 (
            .O(N__41556),
            .I(N__41538));
    InMux I__9234 (
            .O(N__41555),
            .I(N__41535));
    Span4Mux_v I__9233 (
            .O(N__41552),
            .I(N__41530));
    Span4Mux_v I__9232 (
            .O(N__41547),
            .I(N__41530));
    Span4Mux_v I__9231 (
            .O(N__41544),
            .I(N__41525));
    LocalMux I__9230 (
            .O(N__41541),
            .I(N__41525));
    Odrv4 I__9229 (
            .O(N__41538),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9 ));
    LocalMux I__9228 (
            .O(N__41535),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9 ));
    Odrv4 I__9227 (
            .O(N__41530),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9 ));
    Odrv4 I__9226 (
            .O(N__41525),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9 ));
    InMux I__9225 (
            .O(N__41516),
            .I(N__41513));
    LocalMux I__9224 (
            .O(N__41513),
            .I(N__41510));
    Span4Mux_v I__9223 (
            .O(N__41510),
            .I(N__41507));
    Odrv4 I__9222 (
            .O(N__41507),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16 ));
    InMux I__9221 (
            .O(N__41504),
            .I(N__41500));
    InMux I__9220 (
            .O(N__41503),
            .I(N__41493));
    LocalMux I__9219 (
            .O(N__41500),
            .I(N__41490));
    InMux I__9218 (
            .O(N__41499),
            .I(N__41487));
    InMux I__9217 (
            .O(N__41498),
            .I(N__41484));
    CascadeMux I__9216 (
            .O(N__41497),
            .I(N__41481));
    InMux I__9215 (
            .O(N__41496),
            .I(N__41476));
    LocalMux I__9214 (
            .O(N__41493),
            .I(N__41469));
    Span4Mux_h I__9213 (
            .O(N__41490),
            .I(N__41469));
    LocalMux I__9212 (
            .O(N__41487),
            .I(N__41469));
    LocalMux I__9211 (
            .O(N__41484),
            .I(N__41466));
    InMux I__9210 (
            .O(N__41481),
            .I(N__41461));
    InMux I__9209 (
            .O(N__41480),
            .I(N__41461));
    InMux I__9208 (
            .O(N__41479),
            .I(N__41458));
    LocalMux I__9207 (
            .O(N__41476),
            .I(N__41453));
    Span4Mux_v I__9206 (
            .O(N__41469),
            .I(N__41453));
    Span4Mux_h I__9205 (
            .O(N__41466),
            .I(N__41450));
    LocalMux I__9204 (
            .O(N__41461),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ));
    LocalMux I__9203 (
            .O(N__41458),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ));
    Odrv4 I__9202 (
            .O(N__41453),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ));
    Odrv4 I__9201 (
            .O(N__41450),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ));
    InMux I__9200 (
            .O(N__41441),
            .I(N__41438));
    LocalMux I__9199 (
            .O(N__41438),
            .I(N__41435));
    Odrv4 I__9198 (
            .O(N__41435),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1 ));
    InMux I__9197 (
            .O(N__41432),
            .I(N__41427));
    InMux I__9196 (
            .O(N__41431),
            .I(N__41422));
    InMux I__9195 (
            .O(N__41430),
            .I(N__41422));
    LocalMux I__9194 (
            .O(N__41427),
            .I(N__41419));
    LocalMux I__9193 (
            .O(N__41422),
            .I(elapsed_time_ns_1_RNIPFL2M1_0_1));
    Odrv4 I__9192 (
            .O(N__41419),
            .I(elapsed_time_ns_1_RNIPFL2M1_0_1));
    InMux I__9191 (
            .O(N__41414),
            .I(N__41410));
    InMux I__9190 (
            .O(N__41413),
            .I(N__41407));
    LocalMux I__9189 (
            .O(N__41410),
            .I(\phase_controller_inst1.stoper_tr.N_235 ));
    LocalMux I__9188 (
            .O(N__41407),
            .I(\phase_controller_inst1.stoper_tr.N_235 ));
    CascadeMux I__9187 (
            .O(N__41402),
            .I(elapsed_time_ns_1_RNIPFL2M1_0_1_cascade_));
    InMux I__9186 (
            .O(N__41399),
            .I(N__41396));
    LocalMux I__9185 (
            .O(N__41396),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1 ));
    CascadeMux I__9184 (
            .O(N__41393),
            .I(N__41390));
    InMux I__9183 (
            .O(N__41390),
            .I(N__41387));
    LocalMux I__9182 (
            .O(N__41387),
            .I(\phase_controller_inst1.stoper_tr.un6_running_1 ));
    InMux I__9181 (
            .O(N__41384),
            .I(N__41381));
    LocalMux I__9180 (
            .O(N__41381),
            .I(N__41378));
    Odrv4 I__9179 (
            .O(N__41378),
            .I(\current_shift_inst.un4_control_input_1_axb_19 ));
    InMux I__9178 (
            .O(N__41375),
            .I(N__41372));
    LocalMux I__9177 (
            .O(N__41372),
            .I(N__41369));
    Odrv12 I__9176 (
            .O(N__41369),
            .I(\current_shift_inst.un4_control_input_1_axb_21 ));
    InMux I__9175 (
            .O(N__41366),
            .I(N__41363));
    LocalMux I__9174 (
            .O(N__41363),
            .I(N__41360));
    Odrv12 I__9173 (
            .O(N__41360),
            .I(\current_shift_inst.un4_control_input_1_axb_10 ));
    InMux I__9172 (
            .O(N__41357),
            .I(N__41354));
    LocalMux I__9171 (
            .O(N__41354),
            .I(N__41351));
    Span4Mux_v I__9170 (
            .O(N__41351),
            .I(N__41348));
    Odrv4 I__9169 (
            .O(N__41348),
            .I(\current_shift_inst.un4_control_input_1_axb_14 ));
    InMux I__9168 (
            .O(N__41345),
            .I(N__41342));
    LocalMux I__9167 (
            .O(N__41342),
            .I(N__41339));
    Span4Mux_h I__9166 (
            .O(N__41339),
            .I(N__41336));
    Odrv4 I__9165 (
            .O(N__41336),
            .I(\current_shift_inst.un4_control_input_1_axb_18 ));
    InMux I__9164 (
            .O(N__41333),
            .I(N__41330));
    LocalMux I__9163 (
            .O(N__41330),
            .I(N__41327));
    Odrv4 I__9162 (
            .O(N__41327),
            .I(\current_shift_inst.un4_control_input_1_axb_26 ));
    InMux I__9161 (
            .O(N__41324),
            .I(N__41321));
    LocalMux I__9160 (
            .O(N__41321),
            .I(N__41318));
    Odrv12 I__9159 (
            .O(N__41318),
            .I(\current_shift_inst.un4_control_input_1_axb_15 ));
    InMux I__9158 (
            .O(N__41315),
            .I(N__41312));
    LocalMux I__9157 (
            .O(N__41312),
            .I(N__41309));
    Odrv12 I__9156 (
            .O(N__41309),
            .I(\current_shift_inst.un4_control_input_1_axb_24 ));
    InMux I__9155 (
            .O(N__41306),
            .I(N__41303));
    LocalMux I__9154 (
            .O(N__41303),
            .I(N__41300));
    Odrv12 I__9153 (
            .O(N__41300),
            .I(\current_shift_inst.un4_control_input_1_axb_16 ));
    InMux I__9152 (
            .O(N__41297),
            .I(N__41294));
    LocalMux I__9151 (
            .O(N__41294),
            .I(N__41291));
    Odrv4 I__9150 (
            .O(N__41291),
            .I(\current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ));
    CascadeMux I__9149 (
            .O(N__41288),
            .I(N__41285));
    InMux I__9148 (
            .O(N__41285),
            .I(N__41281));
    InMux I__9147 (
            .O(N__41284),
            .I(N__41278));
    LocalMux I__9146 (
            .O(N__41281),
            .I(N__41273));
    LocalMux I__9145 (
            .O(N__41278),
            .I(N__41273));
    Span4Mux_v I__9144 (
            .O(N__41273),
            .I(N__41269));
    InMux I__9143 (
            .O(N__41272),
            .I(N__41266));
    Odrv4 I__9142 (
            .O(N__41269),
            .I(\current_shift_inst.un4_control_input1_29 ));
    LocalMux I__9141 (
            .O(N__41266),
            .I(\current_shift_inst.un4_control_input1_29 ));
    CascadeMux I__9140 (
            .O(N__41261),
            .I(N__41258));
    InMux I__9139 (
            .O(N__41258),
            .I(N__41255));
    LocalMux I__9138 (
            .O(N__41255),
            .I(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ));
    InMux I__9137 (
            .O(N__41252),
            .I(N__41249));
    LocalMux I__9136 (
            .O(N__41249),
            .I(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ));
    CascadeMux I__9135 (
            .O(N__41246),
            .I(N__41243));
    InMux I__9134 (
            .O(N__41243),
            .I(N__41240));
    LocalMux I__9133 (
            .O(N__41240),
            .I(N__41237));
    Odrv4 I__9132 (
            .O(N__41237),
            .I(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ));
    CascadeMux I__9131 (
            .O(N__41234),
            .I(N__41231));
    InMux I__9130 (
            .O(N__41231),
            .I(N__41228));
    LocalMux I__9129 (
            .O(N__41228),
            .I(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ));
    InMux I__9128 (
            .O(N__41225),
            .I(N__41222));
    LocalMux I__9127 (
            .O(N__41222),
            .I(N__41219));
    Odrv4 I__9126 (
            .O(N__41219),
            .I(\current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ));
    CascadeMux I__9125 (
            .O(N__41216),
            .I(N__41212));
    CascadeMux I__9124 (
            .O(N__41215),
            .I(N__41209));
    InMux I__9123 (
            .O(N__41212),
            .I(N__41205));
    InMux I__9122 (
            .O(N__41209),
            .I(N__41202));
    InMux I__9121 (
            .O(N__41208),
            .I(N__41199));
    LocalMux I__9120 (
            .O(N__41205),
            .I(N__41196));
    LocalMux I__9119 (
            .O(N__41202),
            .I(N__41193));
    LocalMux I__9118 (
            .O(N__41199),
            .I(N__41190));
    Span4Mux_h I__9117 (
            .O(N__41196),
            .I(N__41185));
    Span4Mux_v I__9116 (
            .O(N__41193),
            .I(N__41185));
    Span4Mux_v I__9115 (
            .O(N__41190),
            .I(N__41182));
    Odrv4 I__9114 (
            .O(N__41185),
            .I(\current_shift_inst.un4_control_input1_12 ));
    Odrv4 I__9113 (
            .O(N__41182),
            .I(\current_shift_inst.un4_control_input1_12 ));
    CascadeMux I__9112 (
            .O(N__41177),
            .I(N__41174));
    InMux I__9111 (
            .O(N__41174),
            .I(N__41171));
    LocalMux I__9110 (
            .O(N__41171),
            .I(N__41168));
    Odrv4 I__9109 (
            .O(N__41168),
            .I(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ));
    InMux I__9108 (
            .O(N__41165),
            .I(N__41162));
    LocalMux I__9107 (
            .O(N__41162),
            .I(N__41159));
    Odrv12 I__9106 (
            .O(N__41159),
            .I(\current_shift_inst.un4_control_input_1_axb_12 ));
    InMux I__9105 (
            .O(N__41156),
            .I(N__41152));
    InMux I__9104 (
            .O(N__41155),
            .I(N__41149));
    LocalMux I__9103 (
            .O(N__41152),
            .I(N__41145));
    LocalMux I__9102 (
            .O(N__41149),
            .I(N__41142));
    InMux I__9101 (
            .O(N__41148),
            .I(N__41139));
    Span4Mux_h I__9100 (
            .O(N__41145),
            .I(N__41136));
    Odrv12 I__9099 (
            .O(N__41142),
            .I(\current_shift_inst.un4_control_input1_19 ));
    LocalMux I__9098 (
            .O(N__41139),
            .I(\current_shift_inst.un4_control_input1_19 ));
    Odrv4 I__9097 (
            .O(N__41136),
            .I(\current_shift_inst.un4_control_input1_19 ));
    CascadeMux I__9096 (
            .O(N__41129),
            .I(N__41126));
    InMux I__9095 (
            .O(N__41126),
            .I(N__41123));
    LocalMux I__9094 (
            .O(N__41123),
            .I(N__41120));
    Span4Mux_h I__9093 (
            .O(N__41120),
            .I(N__41117));
    Odrv4 I__9092 (
            .O(N__41117),
            .I(\current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ));
    InMux I__9091 (
            .O(N__41114),
            .I(\current_shift_inst.un4_control_input_1_cry_25 ));
    InMux I__9090 (
            .O(N__41111),
            .I(N__41108));
    LocalMux I__9089 (
            .O(N__41108),
            .I(N__41103));
    InMux I__9088 (
            .O(N__41107),
            .I(N__41098));
    InMux I__9087 (
            .O(N__41106),
            .I(N__41098));
    Span4Mux_h I__9086 (
            .O(N__41103),
            .I(N__41095));
    LocalMux I__9085 (
            .O(N__41098),
            .I(N__41092));
    Odrv4 I__9084 (
            .O(N__41095),
            .I(\current_shift_inst.un4_control_input1_28 ));
    Odrv12 I__9083 (
            .O(N__41092),
            .I(\current_shift_inst.un4_control_input1_28 ));
    InMux I__9082 (
            .O(N__41087),
            .I(\current_shift_inst.un4_control_input_1_cry_26 ));
    InMux I__9081 (
            .O(N__41084),
            .I(\current_shift_inst.un4_control_input_1_cry_27 ));
    InMux I__9080 (
            .O(N__41081),
            .I(\current_shift_inst.un4_control_input_1_cry_28 ));
    InMux I__9079 (
            .O(N__41078),
            .I(\current_shift_inst.un4_control_input1_31 ));
    InMux I__9078 (
            .O(N__41075),
            .I(N__41072));
    LocalMux I__9077 (
            .O(N__41072),
            .I(N__41068));
    InMux I__9076 (
            .O(N__41071),
            .I(N__41065));
    Span4Mux_v I__9075 (
            .O(N__41068),
            .I(N__41061));
    LocalMux I__9074 (
            .O(N__41065),
            .I(N__41058));
    InMux I__9073 (
            .O(N__41064),
            .I(N__41055));
    Odrv4 I__9072 (
            .O(N__41061),
            .I(\current_shift_inst.un4_control_input1_21 ));
    Odrv4 I__9071 (
            .O(N__41058),
            .I(\current_shift_inst.un4_control_input1_21 ));
    LocalMux I__9070 (
            .O(N__41055),
            .I(\current_shift_inst.un4_control_input1_21 ));
    CascadeMux I__9069 (
            .O(N__41048),
            .I(N__41045));
    InMux I__9068 (
            .O(N__41045),
            .I(N__41042));
    LocalMux I__9067 (
            .O(N__41042),
            .I(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ));
    InMux I__9066 (
            .O(N__41039),
            .I(N__41036));
    LocalMux I__9065 (
            .O(N__41036),
            .I(N__41033));
    Span4Mux_h I__9064 (
            .O(N__41033),
            .I(N__41030));
    Odrv4 I__9063 (
            .O(N__41030),
            .I(\current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ));
    InMux I__9062 (
            .O(N__41027),
            .I(N__41024));
    LocalMux I__9061 (
            .O(N__41024),
            .I(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ));
    CascadeMux I__9060 (
            .O(N__41021),
            .I(N__41018));
    InMux I__9059 (
            .O(N__41018),
            .I(N__41015));
    LocalMux I__9058 (
            .O(N__41015),
            .I(N__41012));
    Odrv4 I__9057 (
            .O(N__41012),
            .I(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ));
    InMux I__9056 (
            .O(N__41009),
            .I(bfn_17_17_0_));
    InMux I__9055 (
            .O(N__41006),
            .I(\current_shift_inst.un4_control_input_1_cry_17 ));
    InMux I__9054 (
            .O(N__41003),
            .I(N__40999));
    CascadeMux I__9053 (
            .O(N__41002),
            .I(N__40996));
    LocalMux I__9052 (
            .O(N__40999),
            .I(N__40992));
    InMux I__9051 (
            .O(N__40996),
            .I(N__40987));
    InMux I__9050 (
            .O(N__40995),
            .I(N__40987));
    Span4Mux_h I__9049 (
            .O(N__40992),
            .I(N__40984));
    LocalMux I__9048 (
            .O(N__40987),
            .I(N__40981));
    Odrv4 I__9047 (
            .O(N__40984),
            .I(\current_shift_inst.un4_control_input1_20 ));
    Odrv12 I__9046 (
            .O(N__40981),
            .I(\current_shift_inst.un4_control_input1_20 ));
    InMux I__9045 (
            .O(N__40976),
            .I(\current_shift_inst.un4_control_input_1_cry_18 ));
    InMux I__9044 (
            .O(N__40973),
            .I(\current_shift_inst.un4_control_input_1_cry_19 ));
    CascadeMux I__9043 (
            .O(N__40970),
            .I(N__40966));
    InMux I__9042 (
            .O(N__40969),
            .I(N__40960));
    InMux I__9041 (
            .O(N__40966),
            .I(N__40960));
    InMux I__9040 (
            .O(N__40965),
            .I(N__40957));
    LocalMux I__9039 (
            .O(N__40960),
            .I(N__40952));
    LocalMux I__9038 (
            .O(N__40957),
            .I(N__40952));
    Span4Mux_h I__9037 (
            .O(N__40952),
            .I(N__40949));
    Odrv4 I__9036 (
            .O(N__40949),
            .I(\current_shift_inst.un4_control_input1_22 ));
    InMux I__9035 (
            .O(N__40946),
            .I(\current_shift_inst.un4_control_input_1_cry_20 ));
    InMux I__9034 (
            .O(N__40943),
            .I(N__40938));
    InMux I__9033 (
            .O(N__40942),
            .I(N__40935));
    InMux I__9032 (
            .O(N__40941),
            .I(N__40932));
    LocalMux I__9031 (
            .O(N__40938),
            .I(N__40929));
    LocalMux I__9030 (
            .O(N__40935),
            .I(N__40926));
    LocalMux I__9029 (
            .O(N__40932),
            .I(N__40921));
    Span4Mux_h I__9028 (
            .O(N__40929),
            .I(N__40921));
    Odrv4 I__9027 (
            .O(N__40926),
            .I(\current_shift_inst.un4_control_input1_23 ));
    Odrv4 I__9026 (
            .O(N__40921),
            .I(\current_shift_inst.un4_control_input1_23 ));
    InMux I__9025 (
            .O(N__40916),
            .I(\current_shift_inst.un4_control_input_1_cry_21 ));
    InMux I__9024 (
            .O(N__40913),
            .I(N__40906));
    InMux I__9023 (
            .O(N__40912),
            .I(N__40906));
    InMux I__9022 (
            .O(N__40911),
            .I(N__40903));
    LocalMux I__9021 (
            .O(N__40906),
            .I(N__40900));
    LocalMux I__9020 (
            .O(N__40903),
            .I(N__40897));
    Span4Mux_h I__9019 (
            .O(N__40900),
            .I(N__40894));
    Odrv4 I__9018 (
            .O(N__40897),
            .I(\current_shift_inst.un4_control_input1_24 ));
    Odrv4 I__9017 (
            .O(N__40894),
            .I(\current_shift_inst.un4_control_input1_24 ));
    InMux I__9016 (
            .O(N__40889),
            .I(\current_shift_inst.un4_control_input_1_cry_22 ));
    InMux I__9015 (
            .O(N__40886),
            .I(\current_shift_inst.un4_control_input_1_cry_23 ));
    InMux I__9014 (
            .O(N__40883),
            .I(bfn_17_18_0_));
    CascadeMux I__9013 (
            .O(N__40880),
            .I(N__40876));
    InMux I__9012 (
            .O(N__40879),
            .I(N__40872));
    InMux I__9011 (
            .O(N__40876),
            .I(N__40867));
    InMux I__9010 (
            .O(N__40875),
            .I(N__40867));
    LocalMux I__9009 (
            .O(N__40872),
            .I(\current_shift_inst.un4_control_input1_9 ));
    LocalMux I__9008 (
            .O(N__40867),
            .I(\current_shift_inst.un4_control_input1_9 ));
    InMux I__9007 (
            .O(N__40862),
            .I(\current_shift_inst.un4_control_input_1_cry_7 ));
    InMux I__9006 (
            .O(N__40859),
            .I(bfn_17_16_0_));
    InMux I__9005 (
            .O(N__40856),
            .I(\current_shift_inst.un4_control_input_1_cry_9 ));
    InMux I__9004 (
            .O(N__40853),
            .I(\current_shift_inst.un4_control_input_1_cry_10 ));
    InMux I__9003 (
            .O(N__40850),
            .I(\current_shift_inst.un4_control_input_1_cry_11 ));
    InMux I__9002 (
            .O(N__40847),
            .I(\current_shift_inst.un4_control_input_1_cry_12 ));
    InMux I__9001 (
            .O(N__40844),
            .I(\current_shift_inst.un4_control_input_1_cry_13 ));
    InMux I__9000 (
            .O(N__40841),
            .I(\current_shift_inst.un4_control_input_1_cry_14 ));
    InMux I__8999 (
            .O(N__40838),
            .I(\current_shift_inst.un4_control_input_1_cry_15 ));
    InMux I__8998 (
            .O(N__40835),
            .I(N__40832));
    LocalMux I__8997 (
            .O(N__40832),
            .I(N__40829));
    Sp12to4 I__8996 (
            .O(N__40829),
            .I(N__40823));
    CascadeMux I__8995 (
            .O(N__40828),
            .I(N__40820));
    InMux I__8994 (
            .O(N__40827),
            .I(N__40817));
    InMux I__8993 (
            .O(N__40826),
            .I(N__40814));
    Span12Mux_v I__8992 (
            .O(N__40823),
            .I(N__40811));
    InMux I__8991 (
            .O(N__40820),
            .I(N__40808));
    LocalMux I__8990 (
            .O(N__40817),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__8989 (
            .O(N__40814),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    Odrv12 I__8988 (
            .O(N__40811),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__8987 (
            .O(N__40808),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    InMux I__8986 (
            .O(N__40799),
            .I(N__40793));
    InMux I__8985 (
            .O(N__40798),
            .I(N__40793));
    LocalMux I__8984 (
            .O(N__40793),
            .I(N__40789));
    InMux I__8983 (
            .O(N__40792),
            .I(N__40786));
    Odrv4 I__8982 (
            .O(N__40789),
            .I(\current_shift_inst.un4_control_input1_3 ));
    LocalMux I__8981 (
            .O(N__40786),
            .I(\current_shift_inst.un4_control_input1_3 ));
    InMux I__8980 (
            .O(N__40781),
            .I(\current_shift_inst.un4_control_input_1_cry_1 ));
    InMux I__8979 (
            .O(N__40778),
            .I(N__40775));
    LocalMux I__8978 (
            .O(N__40775),
            .I(N__40771));
    InMux I__8977 (
            .O(N__40774),
            .I(N__40768));
    Span4Mux_v I__8976 (
            .O(N__40771),
            .I(N__40763));
    LocalMux I__8975 (
            .O(N__40768),
            .I(N__40763));
    Span4Mux_h I__8974 (
            .O(N__40763),
            .I(N__40759));
    InMux I__8973 (
            .O(N__40762),
            .I(N__40756));
    Odrv4 I__8972 (
            .O(N__40759),
            .I(\current_shift_inst.un4_control_input1_4 ));
    LocalMux I__8971 (
            .O(N__40756),
            .I(\current_shift_inst.un4_control_input1_4 ));
    InMux I__8970 (
            .O(N__40751),
            .I(\current_shift_inst.un4_control_input_1_cry_2 ));
    InMux I__8969 (
            .O(N__40748),
            .I(N__40745));
    LocalMux I__8968 (
            .O(N__40745),
            .I(\current_shift_inst.un4_control_input_1_axb_4 ));
    InMux I__8967 (
            .O(N__40742),
            .I(\current_shift_inst.un4_control_input_1_cry_3 ));
    InMux I__8966 (
            .O(N__40739),
            .I(N__40736));
    LocalMux I__8965 (
            .O(N__40736),
            .I(\current_shift_inst.un4_control_input_1_axb_5 ));
    InMux I__8964 (
            .O(N__40733),
            .I(N__40726));
    InMux I__8963 (
            .O(N__40732),
            .I(N__40726));
    InMux I__8962 (
            .O(N__40731),
            .I(N__40723));
    LocalMux I__8961 (
            .O(N__40726),
            .I(\current_shift_inst.un4_control_input1_6 ));
    LocalMux I__8960 (
            .O(N__40723),
            .I(\current_shift_inst.un4_control_input1_6 ));
    InMux I__8959 (
            .O(N__40718),
            .I(\current_shift_inst.un4_control_input_1_cry_4 ));
    InMux I__8958 (
            .O(N__40715),
            .I(N__40708));
    InMux I__8957 (
            .O(N__40714),
            .I(N__40708));
    InMux I__8956 (
            .O(N__40713),
            .I(N__40705));
    LocalMux I__8955 (
            .O(N__40708),
            .I(\current_shift_inst.un4_control_input1_7 ));
    LocalMux I__8954 (
            .O(N__40705),
            .I(\current_shift_inst.un4_control_input1_7 ));
    InMux I__8953 (
            .O(N__40700),
            .I(\current_shift_inst.un4_control_input_1_cry_5 ));
    InMux I__8952 (
            .O(N__40697),
            .I(N__40690));
    InMux I__8951 (
            .O(N__40696),
            .I(N__40690));
    InMux I__8950 (
            .O(N__40695),
            .I(N__40687));
    LocalMux I__8949 (
            .O(N__40690),
            .I(\current_shift_inst.un4_control_input1_8 ));
    LocalMux I__8948 (
            .O(N__40687),
            .I(\current_shift_inst.un4_control_input1_8 ));
    InMux I__8947 (
            .O(N__40682),
            .I(\current_shift_inst.un4_control_input_1_cry_6 ));
    CascadeMux I__8946 (
            .O(N__40679),
            .I(N__40676));
    InMux I__8945 (
            .O(N__40676),
            .I(N__40673));
    LocalMux I__8944 (
            .O(N__40673),
            .I(N__40670));
    Span4Mux_h I__8943 (
            .O(N__40670),
            .I(N__40667));
    Odrv4 I__8942 (
            .O(N__40667),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ));
    CascadeMux I__8941 (
            .O(N__40664),
            .I(N__40661));
    InMux I__8940 (
            .O(N__40661),
            .I(N__40658));
    LocalMux I__8939 (
            .O(N__40658),
            .I(N__40655));
    Span4Mux_v I__8938 (
            .O(N__40655),
            .I(N__40652));
    Span4Mux_v I__8937 (
            .O(N__40652),
            .I(N__40649));
    Odrv4 I__8936 (
            .O(N__40649),
            .I(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ));
    InMux I__8935 (
            .O(N__40646),
            .I(N__40643));
    LocalMux I__8934 (
            .O(N__40643),
            .I(\current_shift_inst.un4_control_input1_1 ));
    CascadeMux I__8933 (
            .O(N__40640),
            .I(\current_shift_inst.un4_control_input1_1_cascade_ ));
    InMux I__8932 (
            .O(N__40637),
            .I(N__40633));
    CascadeMux I__8931 (
            .O(N__40636),
            .I(N__40630));
    LocalMux I__8930 (
            .O(N__40633),
            .I(N__40627));
    InMux I__8929 (
            .O(N__40630),
            .I(N__40624));
    Sp12to4 I__8928 (
            .O(N__40627),
            .I(N__40619));
    LocalMux I__8927 (
            .O(N__40624),
            .I(N__40619));
    Span12Mux_v I__8926 (
            .O(N__40619),
            .I(N__40616));
    Odrv12 I__8925 (
            .O(N__40616),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    CascadeMux I__8924 (
            .O(N__40613),
            .I(N__40609));
    InMux I__8923 (
            .O(N__40612),
            .I(N__40606));
    InMux I__8922 (
            .O(N__40609),
            .I(N__40602));
    LocalMux I__8921 (
            .O(N__40606),
            .I(N__40598));
    InMux I__8920 (
            .O(N__40605),
            .I(N__40595));
    LocalMux I__8919 (
            .O(N__40602),
            .I(N__40592));
    InMux I__8918 (
            .O(N__40601),
            .I(N__40589));
    Span4Mux_v I__8917 (
            .O(N__40598),
            .I(N__40586));
    LocalMux I__8916 (
            .O(N__40595),
            .I(N__40583));
    Span4Mux_h I__8915 (
            .O(N__40592),
            .I(N__40578));
    LocalMux I__8914 (
            .O(N__40589),
            .I(N__40578));
    Sp12to4 I__8913 (
            .O(N__40586),
            .I(N__40575));
    Span4Mux_v I__8912 (
            .O(N__40583),
            .I(N__40572));
    Odrv4 I__8911 (
            .O(N__40578),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv12 I__8910 (
            .O(N__40575),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__8909 (
            .O(N__40572),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    CascadeMux I__8908 (
            .O(N__40565),
            .I(N__40562));
    InMux I__8907 (
            .O(N__40562),
            .I(N__40559));
    LocalMux I__8906 (
            .O(N__40559),
            .I(N__40556));
    Span4Mux_h I__8905 (
            .O(N__40556),
            .I(N__40553));
    Span4Mux_h I__8904 (
            .O(N__40553),
            .I(N__40550));
    Odrv4 I__8903 (
            .O(N__40550),
            .I(\current_shift_inst.PI_CTRL.integrator_i_30 ));
    InMux I__8902 (
            .O(N__40547),
            .I(N__40543));
    InMux I__8901 (
            .O(N__40546),
            .I(N__40540));
    LocalMux I__8900 (
            .O(N__40543),
            .I(N__40537));
    LocalMux I__8899 (
            .O(N__40540),
            .I(N__40533));
    Span4Mux_v I__8898 (
            .O(N__40537),
            .I(N__40530));
    InMux I__8897 (
            .O(N__40536),
            .I(N__40527));
    Span4Mux_v I__8896 (
            .O(N__40533),
            .I(N__40524));
    Span4Mux_h I__8895 (
            .O(N__40530),
            .I(N__40521));
    LocalMux I__8894 (
            .O(N__40527),
            .I(N__40512));
    Span4Mux_h I__8893 (
            .O(N__40524),
            .I(N__40512));
    Span4Mux_h I__8892 (
            .O(N__40521),
            .I(N__40512));
    InMux I__8891 (
            .O(N__40520),
            .I(N__40507));
    InMux I__8890 (
            .O(N__40519),
            .I(N__40507));
    Odrv4 I__8889 (
            .O(N__40512),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    LocalMux I__8888 (
            .O(N__40507),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    InMux I__8887 (
            .O(N__40502),
            .I(N__40499));
    LocalMux I__8886 (
            .O(N__40499),
            .I(N__40496));
    Span4Mux_v I__8885 (
            .O(N__40496),
            .I(N__40493));
    Span4Mux_h I__8884 (
            .O(N__40493),
            .I(N__40490));
    Span4Mux_h I__8883 (
            .O(N__40490),
            .I(N__40487));
    Odrv4 I__8882 (
            .O(N__40487),
            .I(\current_shift_inst.PI_CTRL.integrator_i_13 ));
    InMux I__8881 (
            .O(N__40484),
            .I(N__40481));
    LocalMux I__8880 (
            .O(N__40481),
            .I(N__40476));
    InMux I__8879 (
            .O(N__40480),
            .I(N__40472));
    InMux I__8878 (
            .O(N__40479),
            .I(N__40469));
    Span12Mux_v I__8877 (
            .O(N__40476),
            .I(N__40466));
    InMux I__8876 (
            .O(N__40475),
            .I(N__40463));
    LocalMux I__8875 (
            .O(N__40472),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__8874 (
            .O(N__40469),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    Odrv12 I__8873 (
            .O(N__40466),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__8872 (
            .O(N__40463),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    InMux I__8871 (
            .O(N__40454),
            .I(N__40451));
    LocalMux I__8870 (
            .O(N__40451),
            .I(N__40448));
    Span4Mux_v I__8869 (
            .O(N__40448),
            .I(N__40445));
    Odrv4 I__8868 (
            .O(N__40445),
            .I(\phase_controller_inst1.stoper_tr.un6_running_18 ));
    CascadeMux I__8867 (
            .O(N__40442),
            .I(N__40439));
    InMux I__8866 (
            .O(N__40439),
            .I(N__40436));
    LocalMux I__8865 (
            .O(N__40436),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ));
    InMux I__8864 (
            .O(N__40433),
            .I(N__40430));
    LocalMux I__8863 (
            .O(N__40430),
            .I(N__40427));
    Span4Mux_v I__8862 (
            .O(N__40427),
            .I(N__40424));
    Odrv4 I__8861 (
            .O(N__40424),
            .I(\phase_controller_inst1.stoper_tr.un6_running_19 ));
    CascadeMux I__8860 (
            .O(N__40421),
            .I(N__40418));
    InMux I__8859 (
            .O(N__40418),
            .I(N__40415));
    LocalMux I__8858 (
            .O(N__40415),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ));
    InMux I__8857 (
            .O(N__40412),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_19 ));
    InMux I__8856 (
            .O(N__40409),
            .I(N__40406));
    LocalMux I__8855 (
            .O(N__40406),
            .I(N__40403));
    Span12Mux_h I__8854 (
            .O(N__40403),
            .I(N__40400));
    Odrv12 I__8853 (
            .O(N__40400),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ));
    InMux I__8852 (
            .O(N__40397),
            .I(N__40394));
    LocalMux I__8851 (
            .O(N__40394),
            .I(N__40391));
    Span4Mux_v I__8850 (
            .O(N__40391),
            .I(N__40388));
    Odrv4 I__8849 (
            .O(N__40388),
            .I(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ));
    CascadeMux I__8848 (
            .O(N__40385),
            .I(N__40382));
    InMux I__8847 (
            .O(N__40382),
            .I(N__40379));
    LocalMux I__8846 (
            .O(N__40379),
            .I(N__40376));
    Span4Mux_v I__8845 (
            .O(N__40376),
            .I(N__40373));
    Odrv4 I__8844 (
            .O(N__40373),
            .I(\phase_controller_inst1.stoper_tr.un6_running_10 ));
    InMux I__8843 (
            .O(N__40370),
            .I(N__40367));
    LocalMux I__8842 (
            .O(N__40367),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    InMux I__8841 (
            .O(N__40364),
            .I(N__40361));
    LocalMux I__8840 (
            .O(N__40361),
            .I(N__40358));
    Span4Mux_h I__8839 (
            .O(N__40358),
            .I(N__40355));
    Odrv4 I__8838 (
            .O(N__40355),
            .I(\phase_controller_inst1.stoper_tr.un6_running_11 ));
    CascadeMux I__8837 (
            .O(N__40352),
            .I(N__40349));
    InMux I__8836 (
            .O(N__40349),
            .I(N__40346));
    LocalMux I__8835 (
            .O(N__40346),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    InMux I__8834 (
            .O(N__40343),
            .I(N__40340));
    LocalMux I__8833 (
            .O(N__40340),
            .I(N__40337));
    Span4Mux_h I__8832 (
            .O(N__40337),
            .I(N__40334));
    Odrv4 I__8831 (
            .O(N__40334),
            .I(\phase_controller_inst1.stoper_tr.un6_running_12 ));
    CascadeMux I__8830 (
            .O(N__40331),
            .I(N__40328));
    InMux I__8829 (
            .O(N__40328),
            .I(N__40325));
    LocalMux I__8828 (
            .O(N__40325),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    InMux I__8827 (
            .O(N__40322),
            .I(N__40319));
    LocalMux I__8826 (
            .O(N__40319),
            .I(N__40316));
    Span4Mux_h I__8825 (
            .O(N__40316),
            .I(N__40313));
    Odrv4 I__8824 (
            .O(N__40313),
            .I(\phase_controller_inst1.stoper_tr.un6_running_13 ));
    CascadeMux I__8823 (
            .O(N__40310),
            .I(N__40307));
    InMux I__8822 (
            .O(N__40307),
            .I(N__40304));
    LocalMux I__8821 (
            .O(N__40304),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    CascadeMux I__8820 (
            .O(N__40301),
            .I(N__40298));
    InMux I__8819 (
            .O(N__40298),
            .I(N__40295));
    LocalMux I__8818 (
            .O(N__40295),
            .I(N__40292));
    Span4Mux_v I__8817 (
            .O(N__40292),
            .I(N__40289));
    Odrv4 I__8816 (
            .O(N__40289),
            .I(\phase_controller_inst1.stoper_tr.un6_running_14 ));
    InMux I__8815 (
            .O(N__40286),
            .I(N__40283));
    LocalMux I__8814 (
            .O(N__40283),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    InMux I__8813 (
            .O(N__40280),
            .I(N__40277));
    LocalMux I__8812 (
            .O(N__40277),
            .I(\phase_controller_inst1.stoper_tr.un6_running_15 ));
    CascadeMux I__8811 (
            .O(N__40274),
            .I(N__40271));
    InMux I__8810 (
            .O(N__40271),
            .I(N__40268));
    LocalMux I__8809 (
            .O(N__40268),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    InMux I__8808 (
            .O(N__40265),
            .I(N__40262));
    LocalMux I__8807 (
            .O(N__40262),
            .I(\phase_controller_inst1.stoper_tr.un6_running_16 ));
    CascadeMux I__8806 (
            .O(N__40259),
            .I(N__40256));
    InMux I__8805 (
            .O(N__40256),
            .I(N__40253));
    LocalMux I__8804 (
            .O(N__40253),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ));
    InMux I__8803 (
            .O(N__40250),
            .I(N__40247));
    LocalMux I__8802 (
            .O(N__40247),
            .I(N__40244));
    Span4Mux_h I__8801 (
            .O(N__40244),
            .I(N__40241));
    Odrv4 I__8800 (
            .O(N__40241),
            .I(\phase_controller_inst1.stoper_tr.un6_running_17 ));
    CascadeMux I__8799 (
            .O(N__40238),
            .I(N__40235));
    InMux I__8798 (
            .O(N__40235),
            .I(N__40232));
    LocalMux I__8797 (
            .O(N__40232),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ));
    CascadeMux I__8796 (
            .O(N__40229),
            .I(N__40226));
    InMux I__8795 (
            .O(N__40226),
            .I(N__40223));
    LocalMux I__8794 (
            .O(N__40223),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    InMux I__8793 (
            .O(N__40220),
            .I(N__40217));
    LocalMux I__8792 (
            .O(N__40217),
            .I(\phase_controller_inst1.stoper_tr.un6_running_3 ));
    CascadeMux I__8791 (
            .O(N__40214),
            .I(N__40211));
    InMux I__8790 (
            .O(N__40211),
            .I(N__40208));
    LocalMux I__8789 (
            .O(N__40208),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    CascadeMux I__8788 (
            .O(N__40205),
            .I(N__40202));
    InMux I__8787 (
            .O(N__40202),
            .I(N__40199));
    LocalMux I__8786 (
            .O(N__40199),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    InMux I__8785 (
            .O(N__40196),
            .I(N__40193));
    LocalMux I__8784 (
            .O(N__40193),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    InMux I__8783 (
            .O(N__40190),
            .I(N__40187));
    LocalMux I__8782 (
            .O(N__40187),
            .I(N__40184));
    Odrv4 I__8781 (
            .O(N__40184),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    CascadeMux I__8780 (
            .O(N__40181),
            .I(N__40178));
    InMux I__8779 (
            .O(N__40178),
            .I(N__40175));
    LocalMux I__8778 (
            .O(N__40175),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    InMux I__8777 (
            .O(N__40172),
            .I(N__40169));
    LocalMux I__8776 (
            .O(N__40169),
            .I(N__40166));
    Span4Mux_h I__8775 (
            .O(N__40166),
            .I(N__40163));
    Odrv4 I__8774 (
            .O(N__40163),
            .I(\phase_controller_inst1.stoper_tr.un6_running_8 ));
    CascadeMux I__8773 (
            .O(N__40160),
            .I(N__40157));
    InMux I__8772 (
            .O(N__40157),
            .I(N__40154));
    LocalMux I__8771 (
            .O(N__40154),
            .I(N__40151));
    Odrv4 I__8770 (
            .O(N__40151),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    InMux I__8769 (
            .O(N__40148),
            .I(N__40145));
    LocalMux I__8768 (
            .O(N__40145),
            .I(\phase_controller_inst1.stoper_tr.un6_running_9 ));
    CascadeMux I__8767 (
            .O(N__40142),
            .I(N__40139));
    InMux I__8766 (
            .O(N__40139),
            .I(N__40136));
    LocalMux I__8765 (
            .O(N__40136),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    InMux I__8764 (
            .O(N__40133),
            .I(N__40128));
    InMux I__8763 (
            .O(N__40132),
            .I(N__40124));
    InMux I__8762 (
            .O(N__40131),
            .I(N__40121));
    LocalMux I__8761 (
            .O(N__40128),
            .I(N__40118));
    InMux I__8760 (
            .O(N__40127),
            .I(N__40115));
    LocalMux I__8759 (
            .O(N__40124),
            .I(N__40110));
    LocalMux I__8758 (
            .O(N__40121),
            .I(N__40110));
    Odrv12 I__8757 (
            .O(N__40118),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ));
    LocalMux I__8756 (
            .O(N__40115),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ));
    Odrv4 I__8755 (
            .O(N__40110),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ));
    InMux I__8754 (
            .O(N__40103),
            .I(N__40100));
    LocalMux I__8753 (
            .O(N__40100),
            .I(N__40097));
    Span4Mux_v I__8752 (
            .O(N__40097),
            .I(N__40092));
    InMux I__8751 (
            .O(N__40096),
            .I(N__40089));
    InMux I__8750 (
            .O(N__40095),
            .I(N__40086));
    Odrv4 I__8749 (
            .O(N__40092),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto15 ));
    LocalMux I__8748 (
            .O(N__40089),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto15 ));
    LocalMux I__8747 (
            .O(N__40086),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto15 ));
    CascadeMux I__8746 (
            .O(N__40079),
            .I(N__40072));
    InMux I__8745 (
            .O(N__40078),
            .I(N__40069));
    InMux I__8744 (
            .O(N__40077),
            .I(N__40063));
    InMux I__8743 (
            .O(N__40076),
            .I(N__40063));
    InMux I__8742 (
            .O(N__40075),
            .I(N__40060));
    InMux I__8741 (
            .O(N__40072),
            .I(N__40053));
    LocalMux I__8740 (
            .O(N__40069),
            .I(N__40049));
    CascadeMux I__8739 (
            .O(N__40068),
            .I(N__40046));
    LocalMux I__8738 (
            .O(N__40063),
            .I(N__40040));
    LocalMux I__8737 (
            .O(N__40060),
            .I(N__40040));
    InMux I__8736 (
            .O(N__40059),
            .I(N__40023));
    InMux I__8735 (
            .O(N__40058),
            .I(N__40023));
    InMux I__8734 (
            .O(N__40057),
            .I(N__40023));
    InMux I__8733 (
            .O(N__40056),
            .I(N__40020));
    LocalMux I__8732 (
            .O(N__40053),
            .I(N__40017));
    InMux I__8731 (
            .O(N__40052),
            .I(N__40014));
    Span4Mux_v I__8730 (
            .O(N__40049),
            .I(N__40011));
    InMux I__8729 (
            .O(N__40046),
            .I(N__40008));
    InMux I__8728 (
            .O(N__40045),
            .I(N__40005));
    Span4Mux_h I__8727 (
            .O(N__40040),
            .I(N__40002));
    InMux I__8726 (
            .O(N__40039),
            .I(N__39995));
    InMux I__8725 (
            .O(N__40038),
            .I(N__39995));
    InMux I__8724 (
            .O(N__40037),
            .I(N__39995));
    InMux I__8723 (
            .O(N__40036),
            .I(N__39980));
    InMux I__8722 (
            .O(N__40035),
            .I(N__39980));
    InMux I__8721 (
            .O(N__40034),
            .I(N__39980));
    InMux I__8720 (
            .O(N__40033),
            .I(N__39980));
    InMux I__8719 (
            .O(N__40032),
            .I(N__39980));
    InMux I__8718 (
            .O(N__40031),
            .I(N__39980));
    InMux I__8717 (
            .O(N__40030),
            .I(N__39980));
    LocalMux I__8716 (
            .O(N__40023),
            .I(N__39975));
    LocalMux I__8715 (
            .O(N__40020),
            .I(N__39975));
    Span4Mux_v I__8714 (
            .O(N__40017),
            .I(N__39970));
    LocalMux I__8713 (
            .O(N__40014),
            .I(N__39970));
    Odrv4 I__8712 (
            .O(N__40011),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__8711 (
            .O(N__40008),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__8710 (
            .O(N__40005),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    Odrv4 I__8709 (
            .O(N__40002),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__8708 (
            .O(N__39995),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__8707 (
            .O(N__39980),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    Odrv4 I__8706 (
            .O(N__39975),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    Odrv4 I__8705 (
            .O(N__39970),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    CascadeMux I__8704 (
            .O(N__39953),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15_cascade_));
    InMux I__8703 (
            .O(N__39950),
            .I(N__39947));
    LocalMux I__8702 (
            .O(N__39947),
            .I(N__39943));
    InMux I__8701 (
            .O(N__39946),
            .I(N__39940));
    Span4Mux_v I__8700 (
            .O(N__39943),
            .I(N__39935));
    LocalMux I__8699 (
            .O(N__39940),
            .I(N__39935));
    Odrv4 I__8698 (
            .O(N__39935),
            .I(\phase_controller_inst1.stoper_tr.N_251 ));
    InMux I__8697 (
            .O(N__39932),
            .I(N__39929));
    LocalMux I__8696 (
            .O(N__39929),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9 ));
    InMux I__8695 (
            .O(N__39926),
            .I(N__39922));
    CascadeMux I__8694 (
            .O(N__39925),
            .I(N__39919));
    LocalMux I__8693 (
            .O(N__39922),
            .I(N__39913));
    InMux I__8692 (
            .O(N__39919),
            .I(N__39908));
    InMux I__8691 (
            .O(N__39918),
            .I(N__39908));
    InMux I__8690 (
            .O(N__39917),
            .I(N__39903));
    InMux I__8689 (
            .O(N__39916),
            .I(N__39903));
    Odrv4 I__8688 (
            .O(N__39913),
            .I(elapsed_time_ns_1_RNI1OL2M1_0_9));
    LocalMux I__8687 (
            .O(N__39908),
            .I(elapsed_time_ns_1_RNI1OL2M1_0_9));
    LocalMux I__8686 (
            .O(N__39903),
            .I(elapsed_time_ns_1_RNI1OL2M1_0_9));
    CascadeMux I__8685 (
            .O(N__39896),
            .I(N__39893));
    InMux I__8684 (
            .O(N__39893),
            .I(N__39886));
    InMux I__8683 (
            .O(N__39892),
            .I(N__39883));
    InMux I__8682 (
            .O(N__39891),
            .I(N__39880));
    InMux I__8681 (
            .O(N__39890),
            .I(N__39875));
    InMux I__8680 (
            .O(N__39889),
            .I(N__39875));
    LocalMux I__8679 (
            .O(N__39886),
            .I(elapsed_time_ns_1_RNIDE4DM1_0_14));
    LocalMux I__8678 (
            .O(N__39883),
            .I(elapsed_time_ns_1_RNIDE4DM1_0_14));
    LocalMux I__8677 (
            .O(N__39880),
            .I(elapsed_time_ns_1_RNIDE4DM1_0_14));
    LocalMux I__8676 (
            .O(N__39875),
            .I(elapsed_time_ns_1_RNIDE4DM1_0_14));
    CascadeMux I__8675 (
            .O(N__39866),
            .I(elapsed_time_ns_1_RNI1OL2M1_0_9_cascade_));
    InMux I__8674 (
            .O(N__39863),
            .I(N__39858));
    InMux I__8673 (
            .O(N__39862),
            .I(N__39855));
    InMux I__8672 (
            .O(N__39861),
            .I(N__39852));
    LocalMux I__8671 (
            .O(N__39858),
            .I(\phase_controller_inst1.stoper_tr.N_244 ));
    LocalMux I__8670 (
            .O(N__39855),
            .I(\phase_controller_inst1.stoper_tr.N_244 ));
    LocalMux I__8669 (
            .O(N__39852),
            .I(\phase_controller_inst1.stoper_tr.N_244 ));
    InMux I__8668 (
            .O(N__39845),
            .I(N__39841));
    InMux I__8667 (
            .O(N__39844),
            .I(N__39836));
    LocalMux I__8666 (
            .O(N__39841),
            .I(N__39833));
    InMux I__8665 (
            .O(N__39840),
            .I(N__39830));
    InMux I__8664 (
            .O(N__39839),
            .I(N__39827));
    LocalMux I__8663 (
            .O(N__39836),
            .I(N__39824));
    Odrv12 I__8662 (
            .O(N__39833),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2Z0Z_9 ));
    LocalMux I__8661 (
            .O(N__39830),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2Z0Z_9 ));
    LocalMux I__8660 (
            .O(N__39827),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2Z0Z_9 ));
    Odrv4 I__8659 (
            .O(N__39824),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2Z0Z_9 ));
    CascadeMux I__8658 (
            .O(N__39815),
            .I(N__39812));
    InMux I__8657 (
            .O(N__39812),
            .I(N__39808));
    CascadeMux I__8656 (
            .O(N__39811),
            .I(N__39803));
    LocalMux I__8655 (
            .O(N__39808),
            .I(N__39797));
    InMux I__8654 (
            .O(N__39807),
            .I(N__39794));
    InMux I__8653 (
            .O(N__39806),
            .I(N__39791));
    InMux I__8652 (
            .O(N__39803),
            .I(N__39786));
    InMux I__8651 (
            .O(N__39802),
            .I(N__39786));
    InMux I__8650 (
            .O(N__39801),
            .I(N__39781));
    InMux I__8649 (
            .O(N__39800),
            .I(N__39781));
    Odrv4 I__8648 (
            .O(N__39797),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    LocalMux I__8647 (
            .O(N__39794),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    LocalMux I__8646 (
            .O(N__39791),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    LocalMux I__8645 (
            .O(N__39786),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    LocalMux I__8644 (
            .O(N__39781),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    CascadeMux I__8643 (
            .O(N__39770),
            .I(\phase_controller_inst1.stoper_tr.N_211_cascade_ ));
    CascadeMux I__8642 (
            .O(N__39767),
            .I(N__39749));
    CascadeMux I__8641 (
            .O(N__39766),
            .I(N__39746));
    CascadeMux I__8640 (
            .O(N__39765),
            .I(N__39739));
    CascadeMux I__8639 (
            .O(N__39764),
            .I(N__39736));
    InMux I__8638 (
            .O(N__39763),
            .I(N__39725));
    InMux I__8637 (
            .O(N__39762),
            .I(N__39725));
    InMux I__8636 (
            .O(N__39761),
            .I(N__39725));
    InMux I__8635 (
            .O(N__39760),
            .I(N__39716));
    InMux I__8634 (
            .O(N__39759),
            .I(N__39716));
    InMux I__8633 (
            .O(N__39758),
            .I(N__39716));
    InMux I__8632 (
            .O(N__39757),
            .I(N__39716));
    CascadeMux I__8631 (
            .O(N__39756),
            .I(N__39710));
    InMux I__8630 (
            .O(N__39755),
            .I(N__39707));
    InMux I__8629 (
            .O(N__39754),
            .I(N__39696));
    InMux I__8628 (
            .O(N__39753),
            .I(N__39696));
    InMux I__8627 (
            .O(N__39752),
            .I(N__39696));
    InMux I__8626 (
            .O(N__39749),
            .I(N__39696));
    InMux I__8625 (
            .O(N__39746),
            .I(N__39696));
    InMux I__8624 (
            .O(N__39745),
            .I(N__39689));
    InMux I__8623 (
            .O(N__39744),
            .I(N__39689));
    InMux I__8622 (
            .O(N__39743),
            .I(N__39689));
    InMux I__8621 (
            .O(N__39742),
            .I(N__39678));
    InMux I__8620 (
            .O(N__39739),
            .I(N__39678));
    InMux I__8619 (
            .O(N__39736),
            .I(N__39678));
    InMux I__8618 (
            .O(N__39735),
            .I(N__39678));
    InMux I__8617 (
            .O(N__39734),
            .I(N__39678));
    InMux I__8616 (
            .O(N__39733),
            .I(N__39673));
    InMux I__8615 (
            .O(N__39732),
            .I(N__39673));
    LocalMux I__8614 (
            .O(N__39725),
            .I(N__39670));
    LocalMux I__8613 (
            .O(N__39716),
            .I(N__39667));
    InMux I__8612 (
            .O(N__39715),
            .I(N__39664));
    InMux I__8611 (
            .O(N__39714),
            .I(N__39659));
    InMux I__8610 (
            .O(N__39713),
            .I(N__39659));
    InMux I__8609 (
            .O(N__39710),
            .I(N__39656));
    LocalMux I__8608 (
            .O(N__39707),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    LocalMux I__8607 (
            .O(N__39696),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    LocalMux I__8606 (
            .O(N__39689),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    LocalMux I__8605 (
            .O(N__39678),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    LocalMux I__8604 (
            .O(N__39673),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    Odrv4 I__8603 (
            .O(N__39670),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    Odrv4 I__8602 (
            .O(N__39667),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    LocalMux I__8601 (
            .O(N__39664),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    LocalMux I__8600 (
            .O(N__39659),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    LocalMux I__8599 (
            .O(N__39656),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    CascadeMux I__8598 (
            .O(N__39635),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_0_6_cascade_ ));
    CascadeMux I__8597 (
            .O(N__39632),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1_cascade_ ));
    InMux I__8596 (
            .O(N__39629),
            .I(N__39626));
    LocalMux I__8595 (
            .O(N__39626),
            .I(N__39623));
    Span4Mux_h I__8594 (
            .O(N__39623),
            .I(N__39620));
    Odrv4 I__8593 (
            .O(N__39620),
            .I(\phase_controller_inst2.stoper_tr.un6_running_1 ));
    InMux I__8592 (
            .O(N__39617),
            .I(N__39614));
    LocalMux I__8591 (
            .O(N__39614),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    InMux I__8590 (
            .O(N__39611),
            .I(N__39608));
    LocalMux I__8589 (
            .O(N__39608),
            .I(N__39605));
    Span4Mux_h I__8588 (
            .O(N__39605),
            .I(N__39602));
    Odrv4 I__8587 (
            .O(N__39602),
            .I(\phase_controller_inst2.stoper_tr.un6_running_8 ));
    InMux I__8586 (
            .O(N__39599),
            .I(N__39596));
    LocalMux I__8585 (
            .O(N__39596),
            .I(N__39593));
    Span4Mux_h I__8584 (
            .O(N__39593),
            .I(N__39590));
    Odrv4 I__8583 (
            .O(N__39590),
            .I(\phase_controller_inst2.stoper_tr.un6_running_2 ));
    InMux I__8582 (
            .O(N__39587),
            .I(N__39584));
    LocalMux I__8581 (
            .O(N__39584),
            .I(N__39581));
    Span4Mux_h I__8580 (
            .O(N__39581),
            .I(N__39578));
    Odrv4 I__8579 (
            .O(N__39578),
            .I(\phase_controller_inst1.stoper_tr.N_219 ));
    InMux I__8578 (
            .O(N__39575),
            .I(N__39571));
    InMux I__8577 (
            .O(N__39574),
            .I(N__39568));
    LocalMux I__8576 (
            .O(N__39571),
            .I(N__39565));
    LocalMux I__8575 (
            .O(N__39568),
            .I(N__39559));
    Span12Mux_v I__8574 (
            .O(N__39565),
            .I(N__39559));
    InMux I__8573 (
            .O(N__39564),
            .I(N__39556));
    Odrv12 I__8572 (
            .O(N__39559),
            .I(elapsed_time_ns_1_RNIAE2591_0_2));
    LocalMux I__8571 (
            .O(N__39556),
            .I(elapsed_time_ns_1_RNIAE2591_0_2));
    InMux I__8570 (
            .O(N__39551),
            .I(N__39546));
    InMux I__8569 (
            .O(N__39550),
            .I(N__39541));
    InMux I__8568 (
            .O(N__39549),
            .I(N__39541));
    LocalMux I__8567 (
            .O(N__39546),
            .I(N__39538));
    LocalMux I__8566 (
            .O(N__39541),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_1Z0Z_2 ));
    Odrv4 I__8565 (
            .O(N__39538),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_1Z0Z_2 ));
    InMux I__8564 (
            .O(N__39533),
            .I(N__39530));
    LocalMux I__8563 (
            .O(N__39530),
            .I(N__39527));
    Span4Mux_v I__8562 (
            .O(N__39527),
            .I(N__39524));
    Odrv4 I__8561 (
            .O(N__39524),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6 ));
    InMux I__8560 (
            .O(N__39521),
            .I(N__39517));
    InMux I__8559 (
            .O(N__39520),
            .I(N__39514));
    LocalMux I__8558 (
            .O(N__39517),
            .I(N__39510));
    LocalMux I__8557 (
            .O(N__39514),
            .I(N__39506));
    InMux I__8556 (
            .O(N__39513),
            .I(N__39503));
    Span4Mux_v I__8555 (
            .O(N__39510),
            .I(N__39500));
    InMux I__8554 (
            .O(N__39509),
            .I(N__39497));
    Span4Mux_h I__8553 (
            .O(N__39506),
            .I(N__39494));
    LocalMux I__8552 (
            .O(N__39503),
            .I(elapsed_time_ns_1_RNIGK2591_0_8));
    Odrv4 I__8551 (
            .O(N__39500),
            .I(elapsed_time_ns_1_RNIGK2591_0_8));
    LocalMux I__8550 (
            .O(N__39497),
            .I(elapsed_time_ns_1_RNIGK2591_0_8));
    Odrv4 I__8549 (
            .O(N__39494),
            .I(elapsed_time_ns_1_RNIGK2591_0_8));
    CascadeMux I__8548 (
            .O(N__39485),
            .I(elapsed_time_ns_1_RNIUKL2M1_0_6_cascade_));
    CascadeMux I__8547 (
            .O(N__39482),
            .I(N__39479));
    InMux I__8546 (
            .O(N__39479),
            .I(N__39474));
    InMux I__8545 (
            .O(N__39478),
            .I(N__39471));
    InMux I__8544 (
            .O(N__39477),
            .I(N__39468));
    LocalMux I__8543 (
            .O(N__39474),
            .I(\phase_controller_inst1.stoper_tr.N_247 ));
    LocalMux I__8542 (
            .O(N__39471),
            .I(\phase_controller_inst1.stoper_tr.N_247 ));
    LocalMux I__8541 (
            .O(N__39468),
            .I(\phase_controller_inst1.stoper_tr.N_247 ));
    CascadeMux I__8540 (
            .O(N__39461),
            .I(\phase_controller_inst1.stoper_tr.N_247_cascade_ ));
    CascadeMux I__8539 (
            .O(N__39458),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6_cascade_ ));
    InMux I__8538 (
            .O(N__39455),
            .I(N__39452));
    LocalMux I__8537 (
            .O(N__39452),
            .I(N__39449));
    Span4Mux_v I__8536 (
            .O(N__39449),
            .I(N__39446));
    Odrv4 I__8535 (
            .O(N__39446),
            .I(\phase_controller_inst2.stoper_tr.un6_running_6 ));
    InMux I__8534 (
            .O(N__39443),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    InMux I__8533 (
            .O(N__39440),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    InMux I__8532 (
            .O(N__39437),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    InMux I__8531 (
            .O(N__39434),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    InMux I__8530 (
            .O(N__39431),
            .I(N__39393));
    InMux I__8529 (
            .O(N__39430),
            .I(N__39393));
    InMux I__8528 (
            .O(N__39429),
            .I(N__39393));
    InMux I__8527 (
            .O(N__39428),
            .I(N__39393));
    InMux I__8526 (
            .O(N__39427),
            .I(N__39388));
    InMux I__8525 (
            .O(N__39426),
            .I(N__39388));
    InMux I__8524 (
            .O(N__39425),
            .I(N__39379));
    InMux I__8523 (
            .O(N__39424),
            .I(N__39379));
    InMux I__8522 (
            .O(N__39423),
            .I(N__39379));
    InMux I__8521 (
            .O(N__39422),
            .I(N__39379));
    InMux I__8520 (
            .O(N__39421),
            .I(N__39370));
    InMux I__8519 (
            .O(N__39420),
            .I(N__39370));
    InMux I__8518 (
            .O(N__39419),
            .I(N__39370));
    InMux I__8517 (
            .O(N__39418),
            .I(N__39370));
    InMux I__8516 (
            .O(N__39417),
            .I(N__39361));
    InMux I__8515 (
            .O(N__39416),
            .I(N__39361));
    InMux I__8514 (
            .O(N__39415),
            .I(N__39361));
    InMux I__8513 (
            .O(N__39414),
            .I(N__39361));
    InMux I__8512 (
            .O(N__39413),
            .I(N__39352));
    InMux I__8511 (
            .O(N__39412),
            .I(N__39352));
    InMux I__8510 (
            .O(N__39411),
            .I(N__39352));
    InMux I__8509 (
            .O(N__39410),
            .I(N__39352));
    InMux I__8508 (
            .O(N__39409),
            .I(N__39343));
    InMux I__8507 (
            .O(N__39408),
            .I(N__39343));
    InMux I__8506 (
            .O(N__39407),
            .I(N__39343));
    InMux I__8505 (
            .O(N__39406),
            .I(N__39343));
    InMux I__8504 (
            .O(N__39405),
            .I(N__39334));
    InMux I__8503 (
            .O(N__39404),
            .I(N__39334));
    InMux I__8502 (
            .O(N__39403),
            .I(N__39334));
    InMux I__8501 (
            .O(N__39402),
            .I(N__39334));
    LocalMux I__8500 (
            .O(N__39393),
            .I(N__39321));
    LocalMux I__8499 (
            .O(N__39388),
            .I(N__39321));
    LocalMux I__8498 (
            .O(N__39379),
            .I(N__39321));
    LocalMux I__8497 (
            .O(N__39370),
            .I(N__39321));
    LocalMux I__8496 (
            .O(N__39361),
            .I(N__39321));
    LocalMux I__8495 (
            .O(N__39352),
            .I(N__39321));
    LocalMux I__8494 (
            .O(N__39343),
            .I(\current_shift_inst.timer_s1.running_i ));
    LocalMux I__8493 (
            .O(N__39334),
            .I(\current_shift_inst.timer_s1.running_i ));
    Odrv12 I__8492 (
            .O(N__39321),
            .I(\current_shift_inst.timer_s1.running_i ));
    InMux I__8491 (
            .O(N__39314),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    CEMux I__8490 (
            .O(N__39311),
            .I(N__39307));
    CEMux I__8489 (
            .O(N__39310),
            .I(N__39304));
    LocalMux I__8488 (
            .O(N__39307),
            .I(N__39299));
    LocalMux I__8487 (
            .O(N__39304),
            .I(N__39296));
    CEMux I__8486 (
            .O(N__39303),
            .I(N__39293));
    CEMux I__8485 (
            .O(N__39302),
            .I(N__39290));
    Span4Mux_v I__8484 (
            .O(N__39299),
            .I(N__39285));
    Span4Mux_v I__8483 (
            .O(N__39296),
            .I(N__39285));
    LocalMux I__8482 (
            .O(N__39293),
            .I(N__39280));
    LocalMux I__8481 (
            .O(N__39290),
            .I(N__39280));
    Odrv4 I__8480 (
            .O(N__39285),
            .I(\current_shift_inst.timer_s1.N_167_i ));
    Odrv4 I__8479 (
            .O(N__39280),
            .I(\current_shift_inst.timer_s1.N_167_i ));
    InMux I__8478 (
            .O(N__39275),
            .I(N__39272));
    LocalMux I__8477 (
            .O(N__39272),
            .I(N__39266));
    InMux I__8476 (
            .O(N__39271),
            .I(N__39263));
    InMux I__8475 (
            .O(N__39270),
            .I(N__39258));
    InMux I__8474 (
            .O(N__39269),
            .I(N__39258));
    Odrv4 I__8473 (
            .O(N__39266),
            .I(elapsed_time_ns_1_RNIIJ4DM1_0_19));
    LocalMux I__8472 (
            .O(N__39263),
            .I(elapsed_time_ns_1_RNIIJ4DM1_0_19));
    LocalMux I__8471 (
            .O(N__39258),
            .I(elapsed_time_ns_1_RNIIJ4DM1_0_19));
    InMux I__8470 (
            .O(N__39251),
            .I(N__39248));
    LocalMux I__8469 (
            .O(N__39248),
            .I(N__39245));
    Span4Mux_h I__8468 (
            .O(N__39245),
            .I(N__39242));
    Span4Mux_v I__8467 (
            .O(N__39242),
            .I(N__39239));
    Odrv4 I__8466 (
            .O(N__39239),
            .I(\phase_controller_inst2.stoper_tr.un6_running_19 ));
    InMux I__8465 (
            .O(N__39236),
            .I(N__39233));
    LocalMux I__8464 (
            .O(N__39233),
            .I(N__39230));
    Span4Mux_h I__8463 (
            .O(N__39230),
            .I(N__39227));
    Span4Mux_v I__8462 (
            .O(N__39227),
            .I(N__39224));
    Odrv4 I__8461 (
            .O(N__39224),
            .I(\phase_controller_inst2.stoper_tr.un6_running_16 ));
    InMux I__8460 (
            .O(N__39221),
            .I(N__39218));
    LocalMux I__8459 (
            .O(N__39218),
            .I(N__39215));
    Span4Mux_v I__8458 (
            .O(N__39215),
            .I(N__39212));
    Odrv4 I__8457 (
            .O(N__39212),
            .I(\phase_controller_inst2.stoper_tr.un6_running_15 ));
    InMux I__8456 (
            .O(N__39209),
            .I(N__39206));
    LocalMux I__8455 (
            .O(N__39206),
            .I(N__39203));
    Span4Mux_v I__8454 (
            .O(N__39203),
            .I(N__39200));
    Odrv4 I__8453 (
            .O(N__39200),
            .I(\phase_controller_inst2.stoper_tr.un6_running_7 ));
    InMux I__8452 (
            .O(N__39197),
            .I(bfn_16_23_0_));
    InMux I__8451 (
            .O(N__39194),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    InMux I__8450 (
            .O(N__39191),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    InMux I__8449 (
            .O(N__39188),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    InMux I__8448 (
            .O(N__39185),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    InMux I__8447 (
            .O(N__39182),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    InMux I__8446 (
            .O(N__39179),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    InMux I__8445 (
            .O(N__39176),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    InMux I__8444 (
            .O(N__39173),
            .I(bfn_16_24_0_));
    InMux I__8443 (
            .O(N__39170),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    InMux I__8442 (
            .O(N__39167),
            .I(bfn_16_22_0_));
    InMux I__8441 (
            .O(N__39164),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    InMux I__8440 (
            .O(N__39161),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    InMux I__8439 (
            .O(N__39158),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    InMux I__8438 (
            .O(N__39155),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    InMux I__8437 (
            .O(N__39152),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    InMux I__8436 (
            .O(N__39149),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    InMux I__8435 (
            .O(N__39146),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    InMux I__8434 (
            .O(N__39143),
            .I(N__39138));
    InMux I__8433 (
            .O(N__39142),
            .I(N__39135));
    InMux I__8432 (
            .O(N__39141),
            .I(N__39132));
    LocalMux I__8431 (
            .O(N__39138),
            .I(N__39127));
    LocalMux I__8430 (
            .O(N__39135),
            .I(N__39127));
    LocalMux I__8429 (
            .O(N__39132),
            .I(N__39121));
    Sp12to4 I__8428 (
            .O(N__39127),
            .I(N__39121));
    InMux I__8427 (
            .O(N__39126),
            .I(N__39118));
    Span12Mux_v I__8426 (
            .O(N__39121),
            .I(N__39115));
    LocalMux I__8425 (
            .O(N__39118),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    Odrv12 I__8424 (
            .O(N__39115),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    InMux I__8423 (
            .O(N__39110),
            .I(N__39107));
    LocalMux I__8422 (
            .O(N__39107),
            .I(N__39104));
    Span4Mux_h I__8421 (
            .O(N__39104),
            .I(N__39101));
    Odrv4 I__8420 (
            .O(N__39101),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ));
    InMux I__8419 (
            .O(N__39098),
            .I(N__39095));
    LocalMux I__8418 (
            .O(N__39095),
            .I(N__39092));
    Odrv4 I__8417 (
            .O(N__39092),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ));
    InMux I__8416 (
            .O(N__39089),
            .I(bfn_16_21_0_));
    InMux I__8415 (
            .O(N__39086),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    InMux I__8414 (
            .O(N__39083),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    InMux I__8413 (
            .O(N__39080),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    InMux I__8412 (
            .O(N__39077),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    InMux I__8411 (
            .O(N__39074),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    InMux I__8410 (
            .O(N__39071),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    InMux I__8409 (
            .O(N__39068),
            .I(N__39052));
    InMux I__8408 (
            .O(N__39067),
            .I(N__39049));
    CascadeMux I__8407 (
            .O(N__39066),
            .I(N__39044));
    CascadeMux I__8406 (
            .O(N__39065),
            .I(N__39040));
    CascadeMux I__8405 (
            .O(N__39064),
            .I(N__39036));
    CascadeMux I__8404 (
            .O(N__39063),
            .I(N__39024));
    CascadeMux I__8403 (
            .O(N__39062),
            .I(N__39020));
    CascadeMux I__8402 (
            .O(N__39061),
            .I(N__39016));
    CascadeMux I__8401 (
            .O(N__39060),
            .I(N__39012));
    InMux I__8400 (
            .O(N__39059),
            .I(N__38998));
    InMux I__8399 (
            .O(N__39058),
            .I(N__38998));
    InMux I__8398 (
            .O(N__39057),
            .I(N__38998));
    InMux I__8397 (
            .O(N__39056),
            .I(N__38998));
    CascadeMux I__8396 (
            .O(N__39055),
            .I(N__38986));
    LocalMux I__8395 (
            .O(N__39052),
            .I(N__38982));
    LocalMux I__8394 (
            .O(N__39049),
            .I(N__38979));
    InMux I__8393 (
            .O(N__39048),
            .I(N__38976));
    InMux I__8392 (
            .O(N__39047),
            .I(N__38960));
    InMux I__8391 (
            .O(N__39044),
            .I(N__38960));
    InMux I__8390 (
            .O(N__39043),
            .I(N__38960));
    InMux I__8389 (
            .O(N__39040),
            .I(N__38960));
    InMux I__8388 (
            .O(N__39039),
            .I(N__38960));
    InMux I__8387 (
            .O(N__39036),
            .I(N__38960));
    InMux I__8386 (
            .O(N__39035),
            .I(N__38960));
    InMux I__8385 (
            .O(N__39034),
            .I(N__38951));
    InMux I__8384 (
            .O(N__39033),
            .I(N__38951));
    InMux I__8383 (
            .O(N__39032),
            .I(N__38951));
    InMux I__8382 (
            .O(N__39031),
            .I(N__38951));
    InMux I__8381 (
            .O(N__39030),
            .I(N__38942));
    InMux I__8380 (
            .O(N__39029),
            .I(N__38942));
    InMux I__8379 (
            .O(N__39028),
            .I(N__38942));
    InMux I__8378 (
            .O(N__39027),
            .I(N__38942));
    InMux I__8377 (
            .O(N__39024),
            .I(N__38925));
    InMux I__8376 (
            .O(N__39023),
            .I(N__38925));
    InMux I__8375 (
            .O(N__39020),
            .I(N__38925));
    InMux I__8374 (
            .O(N__39019),
            .I(N__38925));
    InMux I__8373 (
            .O(N__39016),
            .I(N__38925));
    InMux I__8372 (
            .O(N__39015),
            .I(N__38925));
    InMux I__8371 (
            .O(N__39012),
            .I(N__38925));
    InMux I__8370 (
            .O(N__39011),
            .I(N__38925));
    InMux I__8369 (
            .O(N__39010),
            .I(N__38919));
    InMux I__8368 (
            .O(N__39009),
            .I(N__38912));
    InMux I__8367 (
            .O(N__39008),
            .I(N__38912));
    InMux I__8366 (
            .O(N__39007),
            .I(N__38912));
    LocalMux I__8365 (
            .O(N__38998),
            .I(N__38909));
    InMux I__8364 (
            .O(N__38997),
            .I(N__38906));
    InMux I__8363 (
            .O(N__38996),
            .I(N__38899));
    InMux I__8362 (
            .O(N__38995),
            .I(N__38899));
    InMux I__8361 (
            .O(N__38994),
            .I(N__38899));
    InMux I__8360 (
            .O(N__38993),
            .I(N__38890));
    InMux I__8359 (
            .O(N__38992),
            .I(N__38890));
    InMux I__8358 (
            .O(N__38991),
            .I(N__38890));
    InMux I__8357 (
            .O(N__38990),
            .I(N__38890));
    InMux I__8356 (
            .O(N__38989),
            .I(N__38883));
    InMux I__8355 (
            .O(N__38986),
            .I(N__38883));
    InMux I__8354 (
            .O(N__38985),
            .I(N__38883));
    Span4Mux_s1_h I__8353 (
            .O(N__38982),
            .I(N__38876));
    Span4Mux_s1_v I__8352 (
            .O(N__38979),
            .I(N__38876));
    LocalMux I__8351 (
            .O(N__38976),
            .I(N__38876));
    InMux I__8350 (
            .O(N__38975),
            .I(N__38873));
    LocalMux I__8349 (
            .O(N__38960),
            .I(N__38868));
    LocalMux I__8348 (
            .O(N__38951),
            .I(N__38868));
    LocalMux I__8347 (
            .O(N__38942),
            .I(N__38863));
    LocalMux I__8346 (
            .O(N__38925),
            .I(N__38863));
    CascadeMux I__8345 (
            .O(N__38924),
            .I(N__38859));
    CascadeMux I__8344 (
            .O(N__38923),
            .I(N__38855));
    CascadeMux I__8343 (
            .O(N__38922),
            .I(N__38851));
    LocalMux I__8342 (
            .O(N__38919),
            .I(N__38845));
    LocalMux I__8341 (
            .O(N__38912),
            .I(N__38845));
    Span4Mux_v I__8340 (
            .O(N__38909),
            .I(N__38840));
    LocalMux I__8339 (
            .O(N__38906),
            .I(N__38840));
    LocalMux I__8338 (
            .O(N__38899),
            .I(N__38835));
    LocalMux I__8337 (
            .O(N__38890),
            .I(N__38835));
    LocalMux I__8336 (
            .O(N__38883),
            .I(N__38832));
    Sp12to4 I__8335 (
            .O(N__38876),
            .I(N__38829));
    LocalMux I__8334 (
            .O(N__38873),
            .I(N__38826));
    Span4Mux_v I__8333 (
            .O(N__38868),
            .I(N__38821));
    Span4Mux_v I__8332 (
            .O(N__38863),
            .I(N__38821));
    InMux I__8331 (
            .O(N__38862),
            .I(N__38806));
    InMux I__8330 (
            .O(N__38859),
            .I(N__38806));
    InMux I__8329 (
            .O(N__38858),
            .I(N__38806));
    InMux I__8328 (
            .O(N__38855),
            .I(N__38806));
    InMux I__8327 (
            .O(N__38854),
            .I(N__38806));
    InMux I__8326 (
            .O(N__38851),
            .I(N__38806));
    InMux I__8325 (
            .O(N__38850),
            .I(N__38806));
    Sp12to4 I__8324 (
            .O(N__38845),
            .I(N__38803));
    Sp12to4 I__8323 (
            .O(N__38840),
            .I(N__38800));
    Span12Mux_s9_h I__8322 (
            .O(N__38835),
            .I(N__38795));
    Span12Mux_v I__8321 (
            .O(N__38832),
            .I(N__38790));
    Span12Mux_s11_v I__8320 (
            .O(N__38829),
            .I(N__38790));
    Span12Mux_s11_v I__8319 (
            .O(N__38826),
            .I(N__38783));
    Sp12to4 I__8318 (
            .O(N__38821),
            .I(N__38783));
    LocalMux I__8317 (
            .O(N__38806),
            .I(N__38783));
    Span12Mux_s10_v I__8316 (
            .O(N__38803),
            .I(N__38780));
    Span12Mux_v I__8315 (
            .O(N__38800),
            .I(N__38777));
    InMux I__8314 (
            .O(N__38799),
            .I(N__38772));
    InMux I__8313 (
            .O(N__38798),
            .I(N__38772));
    Span12Mux_v I__8312 (
            .O(N__38795),
            .I(N__38769));
    Span12Mux_h I__8311 (
            .O(N__38790),
            .I(N__38764));
    Span12Mux_h I__8310 (
            .O(N__38783),
            .I(N__38764));
    Span12Mux_h I__8309 (
            .O(N__38780),
            .I(N__38757));
    Span12Mux_h I__8308 (
            .O(N__38777),
            .I(N__38757));
    LocalMux I__8307 (
            .O(N__38772),
            .I(N__38757));
    Odrv12 I__8306 (
            .O(N__38769),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__8305 (
            .O(N__38764),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__8304 (
            .O(N__38757),
            .I(CONSTANT_ONE_NET));
    InMux I__8303 (
            .O(N__38750),
            .I(\current_shift_inst.un10_control_input_cry_30 ));
    CascadeMux I__8302 (
            .O(N__38747),
            .I(N__38744));
    InMux I__8301 (
            .O(N__38744),
            .I(N__38741));
    LocalMux I__8300 (
            .O(N__38741),
            .I(N__38737));
    InMux I__8299 (
            .O(N__38740),
            .I(N__38730));
    Span4Mux_h I__8298 (
            .O(N__38737),
            .I(N__38720));
    InMux I__8297 (
            .O(N__38736),
            .I(N__38711));
    InMux I__8296 (
            .O(N__38735),
            .I(N__38711));
    InMux I__8295 (
            .O(N__38734),
            .I(N__38711));
    InMux I__8294 (
            .O(N__38733),
            .I(N__38711));
    LocalMux I__8293 (
            .O(N__38730),
            .I(N__38708));
    InMux I__8292 (
            .O(N__38729),
            .I(N__38693));
    InMux I__8291 (
            .O(N__38728),
            .I(N__38693));
    InMux I__8290 (
            .O(N__38727),
            .I(N__38693));
    InMux I__8289 (
            .O(N__38726),
            .I(N__38693));
    InMux I__8288 (
            .O(N__38725),
            .I(N__38693));
    InMux I__8287 (
            .O(N__38724),
            .I(N__38693));
    InMux I__8286 (
            .O(N__38723),
            .I(N__38693));
    Odrv4 I__8285 (
            .O(N__38720),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    LocalMux I__8284 (
            .O(N__38711),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__8283 (
            .O(N__38708),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    LocalMux I__8282 (
            .O(N__38693),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    CascadeMux I__8281 (
            .O(N__38684),
            .I(N__38681));
    InMux I__8280 (
            .O(N__38681),
            .I(N__38678));
    LocalMux I__8279 (
            .O(N__38678),
            .I(N__38675));
    Odrv4 I__8278 (
            .O(N__38675),
            .I(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ));
    InMux I__8277 (
            .O(N__38672),
            .I(N__38669));
    LocalMux I__8276 (
            .O(N__38669),
            .I(N__38666));
    Span4Mux_v I__8275 (
            .O(N__38666),
            .I(N__38663));
    Span4Mux_h I__8274 (
            .O(N__38663),
            .I(N__38660));
    Odrv4 I__8273 (
            .O(N__38660),
            .I(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ));
    InMux I__8272 (
            .O(N__38657),
            .I(N__38654));
    LocalMux I__8271 (
            .O(N__38654),
            .I(N__38651));
    Span4Mux_h I__8270 (
            .O(N__38651),
            .I(N__38648));
    Odrv4 I__8269 (
            .O(N__38648),
            .I(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ));
    CascadeMux I__8268 (
            .O(N__38645),
            .I(N__38642));
    InMux I__8267 (
            .O(N__38642),
            .I(N__38639));
    LocalMux I__8266 (
            .O(N__38639),
            .I(N__38636));
    Odrv4 I__8265 (
            .O(N__38636),
            .I(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ));
    InMux I__8264 (
            .O(N__38633),
            .I(N__38630));
    LocalMux I__8263 (
            .O(N__38630),
            .I(N__38627));
    Odrv4 I__8262 (
            .O(N__38627),
            .I(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ));
    InMux I__8261 (
            .O(N__38624),
            .I(N__38621));
    LocalMux I__8260 (
            .O(N__38621),
            .I(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ));
    CascadeMux I__8259 (
            .O(N__38618),
            .I(N__38615));
    InMux I__8258 (
            .O(N__38615),
            .I(N__38612));
    LocalMux I__8257 (
            .O(N__38612),
            .I(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ));
    CascadeMux I__8256 (
            .O(N__38609),
            .I(N__38606));
    InMux I__8255 (
            .O(N__38606),
            .I(N__38603));
    LocalMux I__8254 (
            .O(N__38603),
            .I(N__38600));
    Odrv4 I__8253 (
            .O(N__38600),
            .I(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ));
    CascadeMux I__8252 (
            .O(N__38597),
            .I(N__38594));
    InMux I__8251 (
            .O(N__38594),
            .I(N__38591));
    LocalMux I__8250 (
            .O(N__38591),
            .I(N__38588));
    Span4Mux_h I__8249 (
            .O(N__38588),
            .I(N__38585));
    Odrv4 I__8248 (
            .O(N__38585),
            .I(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ));
    InMux I__8247 (
            .O(N__38582),
            .I(N__38579));
    LocalMux I__8246 (
            .O(N__38579),
            .I(N__38574));
    InMux I__8245 (
            .O(N__38578),
            .I(N__38569));
    InMux I__8244 (
            .O(N__38577),
            .I(N__38569));
    Span4Mux_h I__8243 (
            .O(N__38574),
            .I(N__38566));
    LocalMux I__8242 (
            .O(N__38569),
            .I(N__38563));
    Odrv4 I__8241 (
            .O(N__38566),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    Odrv4 I__8240 (
            .O(N__38563),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    CascadeMux I__8239 (
            .O(N__38558),
            .I(N__38554));
    InMux I__8238 (
            .O(N__38557),
            .I(N__38551));
    InMux I__8237 (
            .O(N__38554),
            .I(N__38548));
    LocalMux I__8236 (
            .O(N__38551),
            .I(N__38545));
    LocalMux I__8235 (
            .O(N__38548),
            .I(N__38542));
    Span4Mux_h I__8234 (
            .O(N__38545),
            .I(N__38537));
    Span4Mux_h I__8233 (
            .O(N__38542),
            .I(N__38537));
    Span4Mux_h I__8232 (
            .O(N__38537),
            .I(N__38534));
    Odrv4 I__8231 (
            .O(N__38534),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    InMux I__8230 (
            .O(N__38531),
            .I(N__38528));
    LocalMux I__8229 (
            .O(N__38528),
            .I(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ));
    CascadeMux I__8228 (
            .O(N__38525),
            .I(N__38522));
    InMux I__8227 (
            .O(N__38522),
            .I(N__38519));
    LocalMux I__8226 (
            .O(N__38519),
            .I(N__38516));
    Odrv4 I__8225 (
            .O(N__38516),
            .I(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ));
    InMux I__8224 (
            .O(N__38513),
            .I(N__38510));
    LocalMux I__8223 (
            .O(N__38510),
            .I(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ));
    CascadeMux I__8222 (
            .O(N__38507),
            .I(N__38504));
    InMux I__8221 (
            .O(N__38504),
            .I(N__38501));
    LocalMux I__8220 (
            .O(N__38501),
            .I(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ));
    InMux I__8219 (
            .O(N__38498),
            .I(N__38495));
    LocalMux I__8218 (
            .O(N__38495),
            .I(N__38492));
    Span4Mux_v I__8217 (
            .O(N__38492),
            .I(N__38489));
    Odrv4 I__8216 (
            .O(N__38489),
            .I(\current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ));
    InMux I__8215 (
            .O(N__38486),
            .I(N__38483));
    LocalMux I__8214 (
            .O(N__38483),
            .I(N__38480));
    Odrv12 I__8213 (
            .O(N__38480),
            .I(\current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ));
    CascadeMux I__8212 (
            .O(N__38477),
            .I(N__38474));
    InMux I__8211 (
            .O(N__38474),
            .I(N__38471));
    LocalMux I__8210 (
            .O(N__38471),
            .I(N__38468));
    Odrv4 I__8209 (
            .O(N__38468),
            .I(\current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ));
    CascadeMux I__8208 (
            .O(N__38465),
            .I(N__38462));
    InMux I__8207 (
            .O(N__38462),
            .I(N__38459));
    LocalMux I__8206 (
            .O(N__38459),
            .I(N__38456));
    Span4Mux_v I__8205 (
            .O(N__38456),
            .I(N__38453));
    Span4Mux_h I__8204 (
            .O(N__38453),
            .I(N__38450));
    Odrv4 I__8203 (
            .O(N__38450),
            .I(\current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ));
    InMux I__8202 (
            .O(N__38447),
            .I(N__38444));
    LocalMux I__8201 (
            .O(N__38444),
            .I(N__38441));
    Odrv4 I__8200 (
            .O(N__38441),
            .I(\current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ));
    InMux I__8199 (
            .O(N__38438),
            .I(N__38435));
    LocalMux I__8198 (
            .O(N__38435),
            .I(N__38432));
    Span4Mux_v I__8197 (
            .O(N__38432),
            .I(N__38429));
    Span4Mux_v I__8196 (
            .O(N__38429),
            .I(N__38424));
    InMux I__8195 (
            .O(N__38428),
            .I(N__38421));
    CascadeMux I__8194 (
            .O(N__38427),
            .I(N__38418));
    Span4Mux_v I__8193 (
            .O(N__38424),
            .I(N__38414));
    LocalMux I__8192 (
            .O(N__38421),
            .I(N__38411));
    InMux I__8191 (
            .O(N__38418),
            .I(N__38406));
    InMux I__8190 (
            .O(N__38417),
            .I(N__38406));
    Odrv4 I__8189 (
            .O(N__38414),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__8188 (
            .O(N__38411),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__8187 (
            .O(N__38406),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    InMux I__8186 (
            .O(N__38399),
            .I(N__38396));
    LocalMux I__8185 (
            .O(N__38396),
            .I(N__38391));
    InMux I__8184 (
            .O(N__38395),
            .I(N__38388));
    InMux I__8183 (
            .O(N__38394),
            .I(N__38385));
    Span4Mux_h I__8182 (
            .O(N__38391),
            .I(N__38378));
    LocalMux I__8181 (
            .O(N__38388),
            .I(N__38378));
    LocalMux I__8180 (
            .O(N__38385),
            .I(N__38378));
    Span4Mux_v I__8179 (
            .O(N__38378),
            .I(N__38375));
    Span4Mux_v I__8178 (
            .O(N__38375),
            .I(N__38372));
    Odrv4 I__8177 (
            .O(N__38372),
            .I(il_min_comp1_D2));
    CascadeMux I__8176 (
            .O(N__38369),
            .I(N__38366));
    InMux I__8175 (
            .O(N__38366),
            .I(N__38360));
    InMux I__8174 (
            .O(N__38365),
            .I(N__38360));
    LocalMux I__8173 (
            .O(N__38360),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    InMux I__8172 (
            .O(N__38357),
            .I(N__38354));
    LocalMux I__8171 (
            .O(N__38354),
            .I(N__38350));
    InMux I__8170 (
            .O(N__38353),
            .I(N__38347));
    Sp12to4 I__8169 (
            .O(N__38350),
            .I(N__38344));
    LocalMux I__8168 (
            .O(N__38347),
            .I(N__38341));
    Odrv12 I__8167 (
            .O(N__38344),
            .I(\phase_controller_inst1.N_56 ));
    Odrv4 I__8166 (
            .O(N__38341),
            .I(\phase_controller_inst1.N_56 ));
    InMux I__8165 (
            .O(N__38336),
            .I(N__38327));
    InMux I__8164 (
            .O(N__38335),
            .I(N__38327));
    InMux I__8163 (
            .O(N__38334),
            .I(N__38327));
    LocalMux I__8162 (
            .O(N__38327),
            .I(\phase_controller_inst1.tr_time_passed ));
    CascadeMux I__8161 (
            .O(N__38324),
            .I(N__38321));
    InMux I__8160 (
            .O(N__38321),
            .I(N__38318));
    LocalMux I__8159 (
            .O(N__38318),
            .I(N__38315));
    Span4Mux_h I__8158 (
            .O(N__38315),
            .I(N__38312));
    Odrv4 I__8157 (
            .O(N__38312),
            .I(\current_shift_inst.un38_control_input_cry_0_s0_sf ));
    CascadeMux I__8156 (
            .O(N__38309),
            .I(N__38306));
    InMux I__8155 (
            .O(N__38306),
            .I(N__38303));
    LocalMux I__8154 (
            .O(N__38303),
            .I(N__38300));
    Odrv4 I__8153 (
            .O(N__38300),
            .I(\current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ));
    InMux I__8152 (
            .O(N__38297),
            .I(N__38294));
    LocalMux I__8151 (
            .O(N__38294),
            .I(N__38291));
    Odrv4 I__8150 (
            .O(N__38291),
            .I(\current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ));
    CascadeMux I__8149 (
            .O(N__38288),
            .I(N__38285));
    InMux I__8148 (
            .O(N__38285),
            .I(N__38282));
    LocalMux I__8147 (
            .O(N__38282),
            .I(N__38279));
    Span4Mux_h I__8146 (
            .O(N__38279),
            .I(N__38276));
    Span4Mux_v I__8145 (
            .O(N__38276),
            .I(N__38273));
    Odrv4 I__8144 (
            .O(N__38273),
            .I(\current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ));
    InMux I__8143 (
            .O(N__38270),
            .I(N__38267));
    LocalMux I__8142 (
            .O(N__38267),
            .I(N__38264));
    Span4Mux_v I__8141 (
            .O(N__38264),
            .I(N__38261));
    Odrv4 I__8140 (
            .O(N__38261),
            .I(\current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ));
    InMux I__8139 (
            .O(N__38258),
            .I(N__38255));
    LocalMux I__8138 (
            .O(N__38255),
            .I(N__38252));
    Span4Mux_h I__8137 (
            .O(N__38252),
            .I(N__38249));
    Odrv4 I__8136 (
            .O(N__38249),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18 ));
    InMux I__8135 (
            .O(N__38246),
            .I(N__38242));
    InMux I__8134 (
            .O(N__38245),
            .I(N__38239));
    LocalMux I__8133 (
            .O(N__38242),
            .I(N__38234));
    LocalMux I__8132 (
            .O(N__38239),
            .I(N__38231));
    InMux I__8131 (
            .O(N__38238),
            .I(N__38226));
    InMux I__8130 (
            .O(N__38237),
            .I(N__38226));
    Span4Mux_v I__8129 (
            .O(N__38234),
            .I(N__38221));
    Span4Mux_v I__8128 (
            .O(N__38231),
            .I(N__38221));
    LocalMux I__8127 (
            .O(N__38226),
            .I(N__38218));
    Odrv4 I__8126 (
            .O(N__38221),
            .I(elapsed_time_ns_1_RNIHI4DM1_0_18));
    Odrv12 I__8125 (
            .O(N__38218),
            .I(elapsed_time_ns_1_RNIHI4DM1_0_18));
    CascadeMux I__8124 (
            .O(N__38213),
            .I(elapsed_time_ns_1_RNIHI4DM1_0_18_cascade_));
    InMux I__8123 (
            .O(N__38210),
            .I(N__38207));
    LocalMux I__8122 (
            .O(N__38207),
            .I(\phase_controller_inst2.stoper_tr.un6_running_18 ));
    InMux I__8121 (
            .O(N__38204),
            .I(N__38200));
    InMux I__8120 (
            .O(N__38203),
            .I(N__38197));
    LocalMux I__8119 (
            .O(N__38200),
            .I(N__38190));
    LocalMux I__8118 (
            .O(N__38197),
            .I(N__38190));
    InMux I__8117 (
            .O(N__38196),
            .I(N__38185));
    InMux I__8116 (
            .O(N__38195),
            .I(N__38185));
    Odrv12 I__8115 (
            .O(N__38190),
            .I(elapsed_time_ns_1_RNIGH4DM1_0_17));
    LocalMux I__8114 (
            .O(N__38185),
            .I(elapsed_time_ns_1_RNIGH4DM1_0_17));
    InMux I__8113 (
            .O(N__38180),
            .I(N__38177));
    LocalMux I__8112 (
            .O(N__38177),
            .I(\phase_controller_inst2.stoper_tr.un6_running_17 ));
    CascadeMux I__8111 (
            .O(N__38174),
            .I(N__38171));
    InMux I__8110 (
            .O(N__38171),
            .I(N__38164));
    InMux I__8109 (
            .O(N__38170),
            .I(N__38161));
    InMux I__8108 (
            .O(N__38169),
            .I(N__38158));
    InMux I__8107 (
            .O(N__38168),
            .I(N__38153));
    InMux I__8106 (
            .O(N__38167),
            .I(N__38153));
    LocalMux I__8105 (
            .O(N__38164),
            .I(N__38150));
    LocalMux I__8104 (
            .O(N__38161),
            .I(N__38147));
    LocalMux I__8103 (
            .O(N__38158),
            .I(N__38144));
    LocalMux I__8102 (
            .O(N__38153),
            .I(N__38139));
    Span4Mux_h I__8101 (
            .O(N__38150),
            .I(N__38139));
    Span4Mux_v I__8100 (
            .O(N__38147),
            .I(N__38136));
    Span4Mux_h I__8099 (
            .O(N__38144),
            .I(N__38131));
    Span4Mux_v I__8098 (
            .O(N__38139),
            .I(N__38131));
    Odrv4 I__8097 (
            .O(N__38136),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    Odrv4 I__8096 (
            .O(N__38131),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    InMux I__8095 (
            .O(N__38126),
            .I(N__38123));
    LocalMux I__8094 (
            .O(N__38123),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9 ));
    CascadeMux I__8093 (
            .O(N__38120),
            .I(elapsed_time_ns_1_RNISCJF91_0_31_cascade_));
    InMux I__8092 (
            .O(N__38117),
            .I(N__38114));
    LocalMux I__8091 (
            .O(N__38114),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9 ));
    InMux I__8090 (
            .O(N__38111),
            .I(N__38105));
    InMux I__8089 (
            .O(N__38110),
            .I(N__38102));
    CascadeMux I__8088 (
            .O(N__38109),
            .I(N__38099));
    CascadeMux I__8087 (
            .O(N__38108),
            .I(N__38096));
    LocalMux I__8086 (
            .O(N__38105),
            .I(N__38084));
    LocalMux I__8085 (
            .O(N__38102),
            .I(N__38084));
    InMux I__8084 (
            .O(N__38099),
            .I(N__38079));
    InMux I__8083 (
            .O(N__38096),
            .I(N__38079));
    InMux I__8082 (
            .O(N__38095),
            .I(N__38068));
    InMux I__8081 (
            .O(N__38094),
            .I(N__38068));
    InMux I__8080 (
            .O(N__38093),
            .I(N__38068));
    InMux I__8079 (
            .O(N__38092),
            .I(N__38068));
    InMux I__8078 (
            .O(N__38091),
            .I(N__38068));
    InMux I__8077 (
            .O(N__38090),
            .I(N__38063));
    InMux I__8076 (
            .O(N__38089),
            .I(N__38063));
    Span4Mux_v I__8075 (
            .O(N__38084),
            .I(N__38060));
    LocalMux I__8074 (
            .O(N__38079),
            .I(\phase_controller_inst1.stoper_tr.N_241 ));
    LocalMux I__8073 (
            .O(N__38068),
            .I(\phase_controller_inst1.stoper_tr.N_241 ));
    LocalMux I__8072 (
            .O(N__38063),
            .I(\phase_controller_inst1.stoper_tr.N_241 ));
    Odrv4 I__8071 (
            .O(N__38060),
            .I(\phase_controller_inst1.stoper_tr.N_241 ));
    CascadeMux I__8070 (
            .O(N__38051),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_ ));
    InMux I__8069 (
            .O(N__38048),
            .I(N__38045));
    LocalMux I__8068 (
            .O(N__38045),
            .I(\phase_controller_inst2.stoper_tr.un6_running_9 ));
    CascadeMux I__8067 (
            .O(N__38042),
            .I(N__38039));
    InMux I__8066 (
            .O(N__38039),
            .I(N__38036));
    LocalMux I__8065 (
            .O(N__38036),
            .I(N__38033));
    Span4Mux_v I__8064 (
            .O(N__38033),
            .I(N__38029));
    InMux I__8063 (
            .O(N__38032),
            .I(N__38026));
    Odrv4 I__8062 (
            .O(N__38029),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    LocalMux I__8061 (
            .O(N__38026),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__8060 (
            .O(N__38021),
            .I(N__38018));
    LocalMux I__8059 (
            .O(N__38018),
            .I(N__38015));
    Span4Mux_v I__8058 (
            .O(N__38015),
            .I(N__38011));
    InMux I__8057 (
            .O(N__38014),
            .I(N__38008));
    Odrv4 I__8056 (
            .O(N__38011),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    LocalMux I__8055 (
            .O(N__38008),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    InMux I__8054 (
            .O(N__38003),
            .I(N__38000));
    LocalMux I__8053 (
            .O(N__38000),
            .I(elapsed_time_ns_1_RNIRAIF91_0_21));
    InMux I__8052 (
            .O(N__37997),
            .I(N__37993));
    InMux I__8051 (
            .O(N__37996),
            .I(N__37990));
    LocalMux I__8050 (
            .O(N__37993),
            .I(N__37987));
    LocalMux I__8049 (
            .O(N__37990),
            .I(elapsed_time_ns_1_RNIRBJF91_0_30));
    Odrv4 I__8048 (
            .O(N__37987),
            .I(elapsed_time_ns_1_RNIRBJF91_0_30));
    InMux I__8047 (
            .O(N__37982),
            .I(N__37978));
    InMux I__8046 (
            .O(N__37981),
            .I(N__37975));
    LocalMux I__8045 (
            .O(N__37978),
            .I(elapsed_time_ns_1_RNI3JIF91_0_29));
    LocalMux I__8044 (
            .O(N__37975),
            .I(elapsed_time_ns_1_RNI3JIF91_0_29));
    CascadeMux I__8043 (
            .O(N__37970),
            .I(elapsed_time_ns_1_RNIRAIF91_0_21_cascade_));
    InMux I__8042 (
            .O(N__37967),
            .I(N__37964));
    LocalMux I__8041 (
            .O(N__37964),
            .I(N__37960));
    InMux I__8040 (
            .O(N__37963),
            .I(N__37957));
    Span4Mux_h I__8039 (
            .O(N__37960),
            .I(N__37954));
    LocalMux I__8038 (
            .O(N__37957),
            .I(elapsed_time_ns_1_RNIQ9IF91_0_20));
    Odrv4 I__8037 (
            .O(N__37954),
            .I(elapsed_time_ns_1_RNIQ9IF91_0_20));
    InMux I__8036 (
            .O(N__37949),
            .I(N__37943));
    InMux I__8035 (
            .O(N__37948),
            .I(N__37943));
    LocalMux I__8034 (
            .O(N__37943),
            .I(elapsed_time_ns_1_RNISBIF91_0_22));
    InMux I__8033 (
            .O(N__37940),
            .I(N__37937));
    LocalMux I__8032 (
            .O(N__37937),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15 ));
    CascadeMux I__8031 (
            .O(N__37934),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15_cascade_ ));
    InMux I__8030 (
            .O(N__37931),
            .I(N__37928));
    LocalMux I__8029 (
            .O(N__37928),
            .I(N__37925));
    Span4Mux_h I__8028 (
            .O(N__37925),
            .I(N__37922));
    Odrv4 I__8027 (
            .O(N__37922),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15 ));
    CascadeMux I__8026 (
            .O(N__37919),
            .I(\phase_controller_inst1.stoper_tr.N_241_cascade_ ));
    InMux I__8025 (
            .O(N__37916),
            .I(N__37913));
    LocalMux I__8024 (
            .O(N__37913),
            .I(N__37910));
    Odrv4 I__8023 (
            .O(N__37910),
            .I(\phase_controller_inst2.stoper_tr.un6_running_14 ));
    CascadeMux I__8022 (
            .O(N__37907),
            .I(N__37904));
    InMux I__8021 (
            .O(N__37904),
            .I(N__37899));
    CascadeMux I__8020 (
            .O(N__37903),
            .I(N__37896));
    CascadeMux I__8019 (
            .O(N__37902),
            .I(N__37893));
    LocalMux I__8018 (
            .O(N__37899),
            .I(N__37890));
    InMux I__8017 (
            .O(N__37896),
            .I(N__37884));
    InMux I__8016 (
            .O(N__37893),
            .I(N__37884));
    Span4Mux_v I__8015 (
            .O(N__37890),
            .I(N__37881));
    InMux I__8014 (
            .O(N__37889),
            .I(N__37878));
    LocalMux I__8013 (
            .O(N__37884),
            .I(N__37875));
    Odrv4 I__8012 (
            .O(N__37881),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ));
    LocalMux I__8011 (
            .O(N__37878),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ));
    Odrv4 I__8010 (
            .O(N__37875),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ));
    InMux I__8009 (
            .O(N__37868),
            .I(N__37865));
    LocalMux I__8008 (
            .O(N__37865),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14 ));
    InMux I__8007 (
            .O(N__37862),
            .I(N__37859));
    LocalMux I__8006 (
            .O(N__37859),
            .I(N__37856));
    Span4Mux_h I__8005 (
            .O(N__37856),
            .I(N__37853));
    Odrv4 I__8004 (
            .O(N__37853),
            .I(\phase_controller_inst2.stoper_tr.un6_running_10 ));
    CascadeMux I__8003 (
            .O(N__37850),
            .I(N__37847));
    InMux I__8002 (
            .O(N__37847),
            .I(N__37844));
    LocalMux I__8001 (
            .O(N__37844),
            .I(N__37841));
    Odrv4 I__8000 (
            .O(N__37841),
            .I(\phase_controller_inst2.stoper_tr.un6_running_11 ));
    CascadeMux I__7999 (
            .O(N__37838),
            .I(N__37835));
    InMux I__7998 (
            .O(N__37835),
            .I(N__37832));
    LocalMux I__7997 (
            .O(N__37832),
            .I(N__37829));
    Odrv4 I__7996 (
            .O(N__37829),
            .I(\phase_controller_inst2.stoper_tr.un6_running_12 ));
    InMux I__7995 (
            .O(N__37826),
            .I(N__37823));
    LocalMux I__7994 (
            .O(N__37823),
            .I(N__37820));
    Odrv4 I__7993 (
            .O(N__37820),
            .I(\phase_controller_inst2.stoper_tr.un6_running_13 ));
    InMux I__7992 (
            .O(N__37817),
            .I(N__37812));
    InMux I__7991 (
            .O(N__37816),
            .I(N__37809));
    InMux I__7990 (
            .O(N__37815),
            .I(N__37806));
    LocalMux I__7989 (
            .O(N__37812),
            .I(elapsed_time_ns_1_RNISAHF91_0_13));
    LocalMux I__7988 (
            .O(N__37809),
            .I(elapsed_time_ns_1_RNISAHF91_0_13));
    LocalMux I__7987 (
            .O(N__37806),
            .I(elapsed_time_ns_1_RNISAHF91_0_13));
    CascadeMux I__7986 (
            .O(N__37799),
            .I(N__37794));
    InMux I__7985 (
            .O(N__37798),
            .I(N__37790));
    InMux I__7984 (
            .O(N__37797),
            .I(N__37787));
    InMux I__7983 (
            .O(N__37794),
            .I(N__37784));
    InMux I__7982 (
            .O(N__37793),
            .I(N__37781));
    LocalMux I__7981 (
            .O(N__37790),
            .I(elapsed_time_ns_1_RNIQ8HF91_0_11));
    LocalMux I__7980 (
            .O(N__37787),
            .I(elapsed_time_ns_1_RNIQ8HF91_0_11));
    LocalMux I__7979 (
            .O(N__37784),
            .I(elapsed_time_ns_1_RNIQ8HF91_0_11));
    LocalMux I__7978 (
            .O(N__37781),
            .I(elapsed_time_ns_1_RNIQ8HF91_0_11));
    CascadeMux I__7977 (
            .O(N__37772),
            .I(N__37766));
    InMux I__7976 (
            .O(N__37771),
            .I(N__37763));
    InMux I__7975 (
            .O(N__37770),
            .I(N__37760));
    InMux I__7974 (
            .O(N__37769),
            .I(N__37757));
    InMux I__7973 (
            .O(N__37766),
            .I(N__37754));
    LocalMux I__7972 (
            .O(N__37763),
            .I(elapsed_time_ns_1_RNIP7HF91_0_10));
    LocalMux I__7971 (
            .O(N__37760),
            .I(elapsed_time_ns_1_RNIP7HF91_0_10));
    LocalMux I__7970 (
            .O(N__37757),
            .I(elapsed_time_ns_1_RNIP7HF91_0_10));
    LocalMux I__7969 (
            .O(N__37754),
            .I(elapsed_time_ns_1_RNIP7HF91_0_10));
    InMux I__7968 (
            .O(N__37745),
            .I(N__37739));
    InMux I__7967 (
            .O(N__37744),
            .I(N__37736));
    InMux I__7966 (
            .O(N__37743),
            .I(N__37733));
    InMux I__7965 (
            .O(N__37742),
            .I(N__37730));
    LocalMux I__7964 (
            .O(N__37739),
            .I(elapsed_time_ns_1_RNIR9HF91_0_12));
    LocalMux I__7963 (
            .O(N__37736),
            .I(elapsed_time_ns_1_RNIR9HF91_0_12));
    LocalMux I__7962 (
            .O(N__37733),
            .I(elapsed_time_ns_1_RNIR9HF91_0_12));
    LocalMux I__7961 (
            .O(N__37730),
            .I(elapsed_time_ns_1_RNIR9HF91_0_12));
    InMux I__7960 (
            .O(N__37721),
            .I(N__37717));
    InMux I__7959 (
            .O(N__37720),
            .I(N__37713));
    LocalMux I__7958 (
            .O(N__37717),
            .I(N__37710));
    InMux I__7957 (
            .O(N__37716),
            .I(N__37707));
    LocalMux I__7956 (
            .O(N__37713),
            .I(N__37704));
    Odrv4 I__7955 (
            .O(N__37710),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    LocalMux I__7954 (
            .O(N__37707),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    Odrv4 I__7953 (
            .O(N__37704),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    CascadeMux I__7952 (
            .O(N__37697),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_ ));
    CascadeMux I__7951 (
            .O(N__37694),
            .I(N__37691));
    InMux I__7950 (
            .O(N__37691),
            .I(N__37688));
    LocalMux I__7949 (
            .O(N__37688),
            .I(N__37683));
    InMux I__7948 (
            .O(N__37687),
            .I(N__37678));
    InMux I__7947 (
            .O(N__37686),
            .I(N__37678));
    Span4Mux_h I__7946 (
            .O(N__37683),
            .I(N__37673));
    LocalMux I__7945 (
            .O(N__37678),
            .I(N__37673));
    Odrv4 I__7944 (
            .O(N__37673),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    CascadeMux I__7943 (
            .O(N__37670),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17_cascade_ ));
    CascadeMux I__7942 (
            .O(N__37667),
            .I(elapsed_time_ns_1_RNIGH4DM1_0_17_cascade_));
    InMux I__7941 (
            .O(N__37664),
            .I(N__37661));
    LocalMux I__7940 (
            .O(N__37661),
            .I(N__37658));
    Span4Mux_h I__7939 (
            .O(N__37658),
            .I(N__37654));
    InMux I__7938 (
            .O(N__37657),
            .I(N__37651));
    Odrv4 I__7937 (
            .O(N__37654),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    LocalMux I__7936 (
            .O(N__37651),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    CascadeMux I__7935 (
            .O(N__37646),
            .I(elapsed_time_ns_1_RNICG2591_0_4_cascade_));
    CascadeMux I__7934 (
            .O(N__37643),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2_cascade_ ));
    CascadeMux I__7933 (
            .O(N__37640),
            .I(elapsed_time_ns_1_RNIDE4DM1_0_14_cascade_));
    CascadeMux I__7932 (
            .O(N__37637),
            .I(N__37634));
    InMux I__7931 (
            .O(N__37634),
            .I(N__37631));
    LocalMux I__7930 (
            .O(N__37631),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ));
    IoInMux I__7929 (
            .O(N__37628),
            .I(N__37625));
    LocalMux I__7928 (
            .O(N__37625),
            .I(N__37622));
    IoSpan4Mux I__7927 (
            .O(N__37622),
            .I(N__37619));
    Sp12to4 I__7926 (
            .O(N__37619),
            .I(N__37616));
    Odrv12 I__7925 (
            .O(N__37616),
            .I(\current_shift_inst.timer_s1.N_166_i ));
    IoInMux I__7924 (
            .O(N__37613),
            .I(N__37610));
    LocalMux I__7923 (
            .O(N__37610),
            .I(N__37607));
    IoSpan4Mux I__7922 (
            .O(N__37607),
            .I(N__37604));
    Span4Mux_s1_v I__7921 (
            .O(N__37604),
            .I(N__37601));
    Span4Mux_v I__7920 (
            .O(N__37601),
            .I(N__37596));
    InMux I__7919 (
            .O(N__37600),
            .I(N__37591));
    InMux I__7918 (
            .O(N__37599),
            .I(N__37591));
    Odrv4 I__7917 (
            .O(N__37596),
            .I(s1_phy_c));
    LocalMux I__7916 (
            .O(N__37591),
            .I(s1_phy_c));
    InMux I__7915 (
            .O(N__37586),
            .I(N__37582));
    InMux I__7914 (
            .O(N__37585),
            .I(N__37579));
    LocalMux I__7913 (
            .O(N__37582),
            .I(N__37576));
    LocalMux I__7912 (
            .O(N__37579),
            .I(N__37573));
    Span4Mux_h I__7911 (
            .O(N__37576),
            .I(N__37568));
    Span4Mux_h I__7910 (
            .O(N__37573),
            .I(N__37568));
    Odrv4 I__7909 (
            .O(N__37568),
            .I(state_ns_i_a3_1));
    CascadeMux I__7908 (
            .O(N__37565),
            .I(N__37562));
    InMux I__7907 (
            .O(N__37562),
            .I(N__37559));
    LocalMux I__7906 (
            .O(N__37559),
            .I(N__37556));
    Span4Mux_v I__7905 (
            .O(N__37556),
            .I(N__37553));
    Span4Mux_v I__7904 (
            .O(N__37553),
            .I(N__37548));
    CascadeMux I__7903 (
            .O(N__37552),
            .I(N__37544));
    InMux I__7902 (
            .O(N__37551),
            .I(N__37539));
    Span4Mux_h I__7901 (
            .O(N__37548),
            .I(N__37536));
    InMux I__7900 (
            .O(N__37547),
            .I(N__37527));
    InMux I__7899 (
            .O(N__37544),
            .I(N__37527));
    InMux I__7898 (
            .O(N__37543),
            .I(N__37527));
    InMux I__7897 (
            .O(N__37542),
            .I(N__37527));
    LocalMux I__7896 (
            .O(N__37539),
            .I(state_3));
    Odrv4 I__7895 (
            .O(N__37536),
            .I(state_3));
    LocalMux I__7894 (
            .O(N__37527),
            .I(state_3));
    InMux I__7893 (
            .O(N__37520),
            .I(N__37515));
    InMux I__7892 (
            .O(N__37519),
            .I(N__37512));
    InMux I__7891 (
            .O(N__37518),
            .I(N__37509));
    LocalMux I__7890 (
            .O(N__37515),
            .I(N__37506));
    LocalMux I__7889 (
            .O(N__37512),
            .I(N__37501));
    LocalMux I__7888 (
            .O(N__37509),
            .I(N__37501));
    Span4Mux_v I__7887 (
            .O(N__37506),
            .I(N__37496));
    Span4Mux_v I__7886 (
            .O(N__37501),
            .I(N__37496));
    Span4Mux_v I__7885 (
            .O(N__37496),
            .I(N__37493));
    Span4Mux_v I__7884 (
            .O(N__37493),
            .I(N__37490));
    Span4Mux_v I__7883 (
            .O(N__37490),
            .I(N__37487));
    Odrv4 I__7882 (
            .O(N__37487),
            .I(il_max_comp1_D2));
    InMux I__7881 (
            .O(N__37484),
            .I(N__37481));
    LocalMux I__7880 (
            .O(N__37481),
            .I(N__37478));
    Span4Mux_v I__7879 (
            .O(N__37478),
            .I(N__37475));
    Span4Mux_v I__7878 (
            .O(N__37475),
            .I(N__37472));
    Odrv4 I__7877 (
            .O(N__37472),
            .I(\phase_controller_inst1.start_timer_hc_0_sqmuxa ));
    InMux I__7876 (
            .O(N__37469),
            .I(N__37466));
    LocalMux I__7875 (
            .O(N__37466),
            .I(N__37463));
    Span4Mux_v I__7874 (
            .O(N__37463),
            .I(N__37460));
    Span4Mux_v I__7873 (
            .O(N__37460),
            .I(N__37456));
    CascadeMux I__7872 (
            .O(N__37459),
            .I(N__37453));
    Span4Mux_v I__7871 (
            .O(N__37456),
            .I(N__37448));
    InMux I__7870 (
            .O(N__37453),
            .I(N__37443));
    InMux I__7869 (
            .O(N__37452),
            .I(N__37443));
    InMux I__7868 (
            .O(N__37451),
            .I(N__37440));
    Odrv4 I__7867 (
            .O(N__37448),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__7866 (
            .O(N__37443),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__7865 (
            .O(N__37440),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    InMux I__7864 (
            .O(N__37433),
            .I(N__37430));
    LocalMux I__7863 (
            .O(N__37430),
            .I(N__37427));
    Span4Mux_v I__7862 (
            .O(N__37427),
            .I(N__37424));
    Span4Mux_v I__7861 (
            .O(N__37424),
            .I(N__37420));
    InMux I__7860 (
            .O(N__37423),
            .I(N__37415));
    Span4Mux_v I__7859 (
            .O(N__37420),
            .I(N__37412));
    InMux I__7858 (
            .O(N__37419),
            .I(N__37409));
    InMux I__7857 (
            .O(N__37418),
            .I(N__37406));
    LocalMux I__7856 (
            .O(N__37415),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    Odrv4 I__7855 (
            .O(N__37412),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__7854 (
            .O(N__37409),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__7853 (
            .O(N__37406),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    InMux I__7852 (
            .O(N__37397),
            .I(N__37394));
    LocalMux I__7851 (
            .O(N__37394),
            .I(N__37389));
    CascadeMux I__7850 (
            .O(N__37393),
            .I(N__37386));
    InMux I__7849 (
            .O(N__37392),
            .I(N__37383));
    Span4Mux_h I__7848 (
            .O(N__37389),
            .I(N__37380));
    InMux I__7847 (
            .O(N__37386),
            .I(N__37377));
    LocalMux I__7846 (
            .O(N__37383),
            .I(N__37374));
    Odrv4 I__7845 (
            .O(N__37380),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    LocalMux I__7844 (
            .O(N__37377),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    Odrv4 I__7843 (
            .O(N__37374),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    InMux I__7842 (
            .O(N__37367),
            .I(N__37364));
    LocalMux I__7841 (
            .O(N__37364),
            .I(N__37361));
    Odrv4 I__7840 (
            .O(N__37361),
            .I(\current_shift_inst.un38_control_input_0_s1_24 ));
    InMux I__7839 (
            .O(N__37358),
            .I(N__37355));
    LocalMux I__7838 (
            .O(N__37355),
            .I(N__37352));
    Odrv4 I__7837 (
            .O(N__37352),
            .I(\current_shift_inst.un38_control_input_0_s0_24 ));
    InMux I__7836 (
            .O(N__37349),
            .I(N__37346));
    LocalMux I__7835 (
            .O(N__37346),
            .I(N__37343));
    Odrv4 I__7834 (
            .O(N__37343),
            .I(\current_shift_inst.control_input_1_axb_4 ));
    InMux I__7833 (
            .O(N__37340),
            .I(N__37337));
    LocalMux I__7832 (
            .O(N__37337),
            .I(N__37334));
    Odrv4 I__7831 (
            .O(N__37334),
            .I(\current_shift_inst.un38_control_input_0_s1_25 ));
    InMux I__7830 (
            .O(N__37331),
            .I(N__37328));
    LocalMux I__7829 (
            .O(N__37328),
            .I(N__37325));
    Odrv4 I__7828 (
            .O(N__37325),
            .I(\current_shift_inst.un38_control_input_0_s0_25 ));
    InMux I__7827 (
            .O(N__37322),
            .I(N__37319));
    LocalMux I__7826 (
            .O(N__37319),
            .I(N__37316));
    Odrv12 I__7825 (
            .O(N__37316),
            .I(\current_shift_inst.control_input_1_axb_5 ));
    CascadeMux I__7824 (
            .O(N__37313),
            .I(N__37310));
    InMux I__7823 (
            .O(N__37310),
            .I(N__37307));
    LocalMux I__7822 (
            .O(N__37307),
            .I(N__37304));
    Odrv4 I__7821 (
            .O(N__37304),
            .I(\current_shift_inst.un38_control_input_0_s0_26 ));
    InMux I__7820 (
            .O(N__37301),
            .I(N__37298));
    LocalMux I__7819 (
            .O(N__37298),
            .I(N__37295));
    Odrv4 I__7818 (
            .O(N__37295),
            .I(\current_shift_inst.un38_control_input_0_s1_26 ));
    InMux I__7817 (
            .O(N__37292),
            .I(N__37289));
    LocalMux I__7816 (
            .O(N__37289),
            .I(N__37286));
    Odrv12 I__7815 (
            .O(N__37286),
            .I(\current_shift_inst.control_input_1_axb_6 ));
    InMux I__7814 (
            .O(N__37283),
            .I(N__37280));
    LocalMux I__7813 (
            .O(N__37280),
            .I(\current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ));
    InMux I__7812 (
            .O(N__37277),
            .I(N__37274));
    LocalMux I__7811 (
            .O(N__37274),
            .I(\current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ));
    CascadeMux I__7810 (
            .O(N__37271),
            .I(N__37268));
    InMux I__7809 (
            .O(N__37268),
            .I(N__37265));
    LocalMux I__7808 (
            .O(N__37265),
            .I(\current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ));
    InMux I__7807 (
            .O(N__37262),
            .I(N__37259));
    LocalMux I__7806 (
            .O(N__37259),
            .I(\current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ));
    CascadeMux I__7805 (
            .O(N__37256),
            .I(N__37253));
    InMux I__7804 (
            .O(N__37253),
            .I(N__37247));
    InMux I__7803 (
            .O(N__37252),
            .I(N__37247));
    LocalMux I__7802 (
            .O(N__37247),
            .I(N__37244));
    Span4Mux_h I__7801 (
            .O(N__37244),
            .I(N__37240));
    InMux I__7800 (
            .O(N__37243),
            .I(N__37237));
    Span4Mux_h I__7799 (
            .O(N__37240),
            .I(N__37234));
    LocalMux I__7798 (
            .O(N__37237),
            .I(elapsed_time_ns_1_RNI81DJ11_0_2));
    Odrv4 I__7797 (
            .O(N__37234),
            .I(elapsed_time_ns_1_RNI81DJ11_0_2));
    InMux I__7796 (
            .O(N__37229),
            .I(N__37226));
    LocalMux I__7795 (
            .O(N__37226),
            .I(N__37222));
    InMux I__7794 (
            .O(N__37225),
            .I(N__37219));
    Span4Mux_v I__7793 (
            .O(N__37222),
            .I(N__37215));
    LocalMux I__7792 (
            .O(N__37219),
            .I(N__37212));
    InMux I__7791 (
            .O(N__37218),
            .I(N__37209));
    Odrv4 I__7790 (
            .O(N__37215),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    Odrv12 I__7789 (
            .O(N__37212),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__7788 (
            .O(N__37209),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    InMux I__7787 (
            .O(N__37202),
            .I(N__37195));
    InMux I__7786 (
            .O(N__37201),
            .I(N__37195));
    CascadeMux I__7785 (
            .O(N__37200),
            .I(N__37192));
    LocalMux I__7784 (
            .O(N__37195),
            .I(N__37189));
    InMux I__7783 (
            .O(N__37192),
            .I(N__37186));
    Span4Mux_h I__7782 (
            .O(N__37189),
            .I(N__37183));
    LocalMux I__7781 (
            .O(N__37186),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    Odrv4 I__7780 (
            .O(N__37183),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    CEMux I__7779 (
            .O(N__37178),
            .I(N__37163));
    CEMux I__7778 (
            .O(N__37177),
            .I(N__37163));
    CEMux I__7777 (
            .O(N__37176),
            .I(N__37163));
    CEMux I__7776 (
            .O(N__37175),
            .I(N__37163));
    CEMux I__7775 (
            .O(N__37174),
            .I(N__37163));
    GlobalMux I__7774 (
            .O(N__37163),
            .I(N__37160));
    gio2CtrlBuf I__7773 (
            .O(N__37160),
            .I(\delay_measurement_inst.delay_hc_timer.N_432_i_g ));
    InMux I__7772 (
            .O(N__37157),
            .I(N__37148));
    InMux I__7771 (
            .O(N__37156),
            .I(N__37148));
    CascadeMux I__7770 (
            .O(N__37155),
            .I(N__37138));
    InMux I__7769 (
            .O(N__37154),
            .I(N__37135));
    CascadeMux I__7768 (
            .O(N__37153),
            .I(N__37132));
    LocalMux I__7767 (
            .O(N__37148),
            .I(N__37128));
    InMux I__7766 (
            .O(N__37147),
            .I(N__37125));
    InMux I__7765 (
            .O(N__37146),
            .I(N__37122));
    InMux I__7764 (
            .O(N__37145),
            .I(N__37119));
    InMux I__7763 (
            .O(N__37144),
            .I(N__37116));
    InMux I__7762 (
            .O(N__37143),
            .I(N__37107));
    InMux I__7761 (
            .O(N__37142),
            .I(N__37107));
    InMux I__7760 (
            .O(N__37141),
            .I(N__37107));
    InMux I__7759 (
            .O(N__37138),
            .I(N__37107));
    LocalMux I__7758 (
            .O(N__37135),
            .I(N__37099));
    InMux I__7757 (
            .O(N__37132),
            .I(N__37096));
    InMux I__7756 (
            .O(N__37131),
            .I(N__37093));
    Span4Mux_h I__7755 (
            .O(N__37128),
            .I(N__37090));
    LocalMux I__7754 (
            .O(N__37125),
            .I(N__37079));
    LocalMux I__7753 (
            .O(N__37122),
            .I(N__37079));
    LocalMux I__7752 (
            .O(N__37119),
            .I(N__37079));
    LocalMux I__7751 (
            .O(N__37116),
            .I(N__37079));
    LocalMux I__7750 (
            .O(N__37107),
            .I(N__37079));
    InMux I__7749 (
            .O(N__37106),
            .I(N__37072));
    InMux I__7748 (
            .O(N__37105),
            .I(N__37069));
    InMux I__7747 (
            .O(N__37104),
            .I(N__37066));
    InMux I__7746 (
            .O(N__37103),
            .I(N__37061));
    InMux I__7745 (
            .O(N__37102),
            .I(N__37061));
    Span4Mux_h I__7744 (
            .O(N__37099),
            .I(N__37058));
    LocalMux I__7743 (
            .O(N__37096),
            .I(N__37049));
    LocalMux I__7742 (
            .O(N__37093),
            .I(N__37049));
    Span4Mux_v I__7741 (
            .O(N__37090),
            .I(N__37049));
    Span4Mux_v I__7740 (
            .O(N__37079),
            .I(N__37049));
    InMux I__7739 (
            .O(N__37078),
            .I(N__37040));
    InMux I__7738 (
            .O(N__37077),
            .I(N__37040));
    InMux I__7737 (
            .O(N__37076),
            .I(N__37040));
    InMux I__7736 (
            .O(N__37075),
            .I(N__37040));
    LocalMux I__7735 (
            .O(N__37072),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    LocalMux I__7734 (
            .O(N__37069),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    LocalMux I__7733 (
            .O(N__37066),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    LocalMux I__7732 (
            .O(N__37061),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    Odrv4 I__7731 (
            .O(N__37058),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    Odrv4 I__7730 (
            .O(N__37049),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    LocalMux I__7729 (
            .O(N__37040),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    CascadeMux I__7728 (
            .O(N__37025),
            .I(N__37022));
    InMux I__7727 (
            .O(N__37022),
            .I(N__37019));
    LocalMux I__7726 (
            .O(N__37019),
            .I(N__37015));
    CascadeMux I__7725 (
            .O(N__37018),
            .I(N__37012));
    Span12Mux_h I__7724 (
            .O(N__37015),
            .I(N__37009));
    InMux I__7723 (
            .O(N__37012),
            .I(N__37006));
    Odrv12 I__7722 (
            .O(N__37009),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    LocalMux I__7721 (
            .O(N__37006),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    InMux I__7720 (
            .O(N__37001),
            .I(N__36991));
    CascadeMux I__7719 (
            .O(N__37000),
            .I(N__36988));
    CascadeMux I__7718 (
            .O(N__36999),
            .I(N__36985));
    InMux I__7717 (
            .O(N__36998),
            .I(N__36975));
    InMux I__7716 (
            .O(N__36997),
            .I(N__36975));
    CascadeMux I__7715 (
            .O(N__36996),
            .I(N__36971));
    CascadeMux I__7714 (
            .O(N__36995),
            .I(N__36966));
    CascadeMux I__7713 (
            .O(N__36994),
            .I(N__36963));
    LocalMux I__7712 (
            .O(N__36991),
            .I(N__36958));
    InMux I__7711 (
            .O(N__36988),
            .I(N__36953));
    InMux I__7710 (
            .O(N__36985),
            .I(N__36953));
    InMux I__7709 (
            .O(N__36984),
            .I(N__36948));
    InMux I__7708 (
            .O(N__36983),
            .I(N__36948));
    CascadeMux I__7707 (
            .O(N__36982),
            .I(N__36945));
    InMux I__7706 (
            .O(N__36981),
            .I(N__36941));
    InMux I__7705 (
            .O(N__36980),
            .I(N__36938));
    LocalMux I__7704 (
            .O(N__36975),
            .I(N__36935));
    InMux I__7703 (
            .O(N__36974),
            .I(N__36929));
    InMux I__7702 (
            .O(N__36971),
            .I(N__36929));
    InMux I__7701 (
            .O(N__36970),
            .I(N__36926));
    InMux I__7700 (
            .O(N__36969),
            .I(N__36921));
    InMux I__7699 (
            .O(N__36966),
            .I(N__36921));
    InMux I__7698 (
            .O(N__36963),
            .I(N__36918));
    InMux I__7697 (
            .O(N__36962),
            .I(N__36913));
    InMux I__7696 (
            .O(N__36961),
            .I(N__36913));
    Span4Mux_h I__7695 (
            .O(N__36958),
            .I(N__36906));
    LocalMux I__7694 (
            .O(N__36953),
            .I(N__36906));
    LocalMux I__7693 (
            .O(N__36948),
            .I(N__36906));
    InMux I__7692 (
            .O(N__36945),
            .I(N__36903));
    InMux I__7691 (
            .O(N__36944),
            .I(N__36900));
    LocalMux I__7690 (
            .O(N__36941),
            .I(N__36892));
    LocalMux I__7689 (
            .O(N__36938),
            .I(N__36887));
    Span4Mux_h I__7688 (
            .O(N__36935),
            .I(N__36887));
    InMux I__7687 (
            .O(N__36934),
            .I(N__36884));
    LocalMux I__7686 (
            .O(N__36929),
            .I(N__36869));
    LocalMux I__7685 (
            .O(N__36926),
            .I(N__36869));
    LocalMux I__7684 (
            .O(N__36921),
            .I(N__36869));
    LocalMux I__7683 (
            .O(N__36918),
            .I(N__36869));
    LocalMux I__7682 (
            .O(N__36913),
            .I(N__36869));
    Span4Mux_h I__7681 (
            .O(N__36906),
            .I(N__36869));
    LocalMux I__7680 (
            .O(N__36903),
            .I(N__36869));
    LocalMux I__7679 (
            .O(N__36900),
            .I(N__36861));
    InMux I__7678 (
            .O(N__36899),
            .I(N__36856));
    InMux I__7677 (
            .O(N__36898),
            .I(N__36856));
    InMux I__7676 (
            .O(N__36897),
            .I(N__36849));
    InMux I__7675 (
            .O(N__36896),
            .I(N__36849));
    InMux I__7674 (
            .O(N__36895),
            .I(N__36849));
    Span4Mux_v I__7673 (
            .O(N__36892),
            .I(N__36840));
    Span4Mux_v I__7672 (
            .O(N__36887),
            .I(N__36840));
    LocalMux I__7671 (
            .O(N__36884),
            .I(N__36840));
    Span4Mux_v I__7670 (
            .O(N__36869),
            .I(N__36840));
    InMux I__7669 (
            .O(N__36868),
            .I(N__36829));
    InMux I__7668 (
            .O(N__36867),
            .I(N__36829));
    InMux I__7667 (
            .O(N__36866),
            .I(N__36829));
    InMux I__7666 (
            .O(N__36865),
            .I(N__36829));
    InMux I__7665 (
            .O(N__36864),
            .I(N__36829));
    Span4Mux_h I__7664 (
            .O(N__36861),
            .I(N__36826));
    LocalMux I__7663 (
            .O(N__36856),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    LocalMux I__7662 (
            .O(N__36849),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    Odrv4 I__7661 (
            .O(N__36840),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    LocalMux I__7660 (
            .O(N__36829),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    Odrv4 I__7659 (
            .O(N__36826),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    InMux I__7658 (
            .O(N__36815),
            .I(N__36812));
    LocalMux I__7657 (
            .O(N__36812),
            .I(N__36809));
    Span4Mux_h I__7656 (
            .O(N__36809),
            .I(N__36805));
    InMux I__7655 (
            .O(N__36808),
            .I(N__36802));
    Span4Mux_h I__7654 (
            .O(N__36805),
            .I(N__36799));
    LocalMux I__7653 (
            .O(N__36802),
            .I(elapsed_time_ns_1_RNIO1ND11_0_20));
    Odrv4 I__7652 (
            .O(N__36799),
            .I(elapsed_time_ns_1_RNIO1ND11_0_20));
    InMux I__7651 (
            .O(N__36794),
            .I(N__36791));
    LocalMux I__7650 (
            .O(N__36791),
            .I(N__36788));
    Odrv4 I__7649 (
            .O(N__36788),
            .I(\current_shift_inst.un38_control_input_0_s0_20 ));
    InMux I__7648 (
            .O(N__36785),
            .I(N__36782));
    LocalMux I__7647 (
            .O(N__36782),
            .I(\current_shift_inst.un38_control_input_0_s1_20 ));
    InMux I__7646 (
            .O(N__36779),
            .I(N__36776));
    LocalMux I__7645 (
            .O(N__36776),
            .I(N__36773));
    Span4Mux_h I__7644 (
            .O(N__36773),
            .I(N__36770));
    Odrv4 I__7643 (
            .O(N__36770),
            .I(\current_shift_inst.control_input_1_axb_0 ));
    InMux I__7642 (
            .O(N__36767),
            .I(N__36764));
    LocalMux I__7641 (
            .O(N__36764),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ));
    InMux I__7640 (
            .O(N__36761),
            .I(N__36758));
    LocalMux I__7639 (
            .O(N__36758),
            .I(N__36755));
    Odrv4 I__7638 (
            .O(N__36755),
            .I(\current_shift_inst.un38_control_input_0_s0_21 ));
    InMux I__7637 (
            .O(N__36752),
            .I(N__36749));
    LocalMux I__7636 (
            .O(N__36749),
            .I(\current_shift_inst.un38_control_input_0_s1_21 ));
    CascadeMux I__7635 (
            .O(N__36746),
            .I(N__36743));
    InMux I__7634 (
            .O(N__36743),
            .I(N__36740));
    LocalMux I__7633 (
            .O(N__36740),
            .I(N__36737));
    Odrv4 I__7632 (
            .O(N__36737),
            .I(\current_shift_inst.control_input_1_axb_1 ));
    InMux I__7631 (
            .O(N__36734),
            .I(N__36731));
    LocalMux I__7630 (
            .O(N__36731),
            .I(N__36728));
    Odrv4 I__7629 (
            .O(N__36728),
            .I(\current_shift_inst.un38_control_input_0_s0_22 ));
    InMux I__7628 (
            .O(N__36725),
            .I(N__36722));
    LocalMux I__7627 (
            .O(N__36722),
            .I(\current_shift_inst.un38_control_input_0_s1_22 ));
    InMux I__7626 (
            .O(N__36719),
            .I(N__36716));
    LocalMux I__7625 (
            .O(N__36716),
            .I(N__36713));
    Span4Mux_h I__7624 (
            .O(N__36713),
            .I(N__36710));
    Odrv4 I__7623 (
            .O(N__36710),
            .I(\current_shift_inst.control_input_1_axb_2 ));
    InMux I__7622 (
            .O(N__36707),
            .I(N__36704));
    LocalMux I__7621 (
            .O(N__36704),
            .I(\current_shift_inst.un38_control_input_0_s1_23 ));
    InMux I__7620 (
            .O(N__36701),
            .I(N__36698));
    LocalMux I__7619 (
            .O(N__36698),
            .I(N__36695));
    Odrv4 I__7618 (
            .O(N__36695),
            .I(\current_shift_inst.un38_control_input_0_s0_23 ));
    InMux I__7617 (
            .O(N__36692),
            .I(N__36689));
    LocalMux I__7616 (
            .O(N__36689),
            .I(N__36686));
    Odrv12 I__7615 (
            .O(N__36686),
            .I(\current_shift_inst.control_input_1_axb_3 ));
    InMux I__7614 (
            .O(N__36683),
            .I(N__36680));
    LocalMux I__7613 (
            .O(N__36680),
            .I(N__36677));
    Odrv4 I__7612 (
            .O(N__36677),
            .I(\current_shift_inst.control_input_1_axb_11 ));
    InMux I__7611 (
            .O(N__36674),
            .I(\current_shift_inst.control_input_1_cry_10 ));
    InMux I__7610 (
            .O(N__36671),
            .I(N__36668));
    LocalMux I__7609 (
            .O(N__36668),
            .I(N__36665));
    Span4Mux_v I__7608 (
            .O(N__36665),
            .I(N__36661));
    InMux I__7607 (
            .O(N__36664),
            .I(N__36658));
    Span4Mux_v I__7606 (
            .O(N__36661),
            .I(N__36653));
    LocalMux I__7605 (
            .O(N__36658),
            .I(N__36653));
    Odrv4 I__7604 (
            .O(N__36653),
            .I(\current_shift_inst.control_inputZ0Z_11 ));
    CascadeMux I__7603 (
            .O(N__36650),
            .I(N__36647));
    InMux I__7602 (
            .O(N__36647),
            .I(N__36644));
    LocalMux I__7601 (
            .O(N__36644),
            .I(N__36641));
    Odrv4 I__7600 (
            .O(N__36641),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ));
    CascadeMux I__7599 (
            .O(N__36638),
            .I(N__36634));
    InMux I__7598 (
            .O(N__36637),
            .I(N__36631));
    InMux I__7597 (
            .O(N__36634),
            .I(N__36628));
    LocalMux I__7596 (
            .O(N__36631),
            .I(\current_shift_inst.N_1609_i ));
    LocalMux I__7595 (
            .O(N__36628),
            .I(\current_shift_inst.N_1609_i ));
    CascadeMux I__7594 (
            .O(N__36623),
            .I(N__36620));
    InMux I__7593 (
            .O(N__36620),
            .I(N__36617));
    LocalMux I__7592 (
            .O(N__36617),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ));
    InMux I__7591 (
            .O(N__36614),
            .I(N__36611));
    LocalMux I__7590 (
            .O(N__36611),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ));
    InMux I__7589 (
            .O(N__36608),
            .I(N__36605));
    LocalMux I__7588 (
            .O(N__36605),
            .I(\current_shift_inst.un38_control_input_0_s0_27 ));
    InMux I__7587 (
            .O(N__36602),
            .I(N__36599));
    LocalMux I__7586 (
            .O(N__36599),
            .I(N__36596));
    Odrv4 I__7585 (
            .O(N__36596),
            .I(\current_shift_inst.un38_control_input_0_s1_27 ));
    InMux I__7584 (
            .O(N__36593),
            .I(N__36590));
    LocalMux I__7583 (
            .O(N__36590),
            .I(N__36587));
    Odrv4 I__7582 (
            .O(N__36587),
            .I(\current_shift_inst.control_input_1_axb_7 ));
    InMux I__7581 (
            .O(N__36584),
            .I(N__36581));
    LocalMux I__7580 (
            .O(N__36581),
            .I(N__36578));
    Span4Mux_v I__7579 (
            .O(N__36578),
            .I(N__36575));
    Odrv4 I__7578 (
            .O(N__36575),
            .I(\current_shift_inst.un38_control_input_0_s1_28 ));
    InMux I__7577 (
            .O(N__36572),
            .I(N__36569));
    LocalMux I__7576 (
            .O(N__36569),
            .I(\current_shift_inst.un38_control_input_0_s0_28 ));
    InMux I__7575 (
            .O(N__36566),
            .I(N__36563));
    LocalMux I__7574 (
            .O(N__36563),
            .I(\current_shift_inst.control_input_1_axb_8 ));
    InMux I__7573 (
            .O(N__36560),
            .I(N__36557));
    LocalMux I__7572 (
            .O(N__36557),
            .I(\current_shift_inst.un38_control_input_0_s0_29 ));
    InMux I__7571 (
            .O(N__36554),
            .I(N__36551));
    LocalMux I__7570 (
            .O(N__36551),
            .I(N__36548));
    Span4Mux_v I__7569 (
            .O(N__36548),
            .I(N__36545));
    Odrv4 I__7568 (
            .O(N__36545),
            .I(\current_shift_inst.un38_control_input_0_s1_29 ));
    InMux I__7567 (
            .O(N__36542),
            .I(N__36539));
    LocalMux I__7566 (
            .O(N__36539),
            .I(\current_shift_inst.control_input_1_axb_9 ));
    InMux I__7565 (
            .O(N__36536),
            .I(N__36533));
    LocalMux I__7564 (
            .O(N__36533),
            .I(N__36530));
    Span4Mux_h I__7563 (
            .O(N__36530),
            .I(N__36527));
    Odrv4 I__7562 (
            .O(N__36527),
            .I(\current_shift_inst.un38_control_input_0_s1_30 ));
    InMux I__7561 (
            .O(N__36524),
            .I(N__36521));
    LocalMux I__7560 (
            .O(N__36521),
            .I(\current_shift_inst.un38_control_input_0_s0_30 ));
    InMux I__7559 (
            .O(N__36518),
            .I(N__36515));
    LocalMux I__7558 (
            .O(N__36515),
            .I(\current_shift_inst.control_input_1_axb_10 ));
    InMux I__7557 (
            .O(N__36512),
            .I(N__36509));
    LocalMux I__7556 (
            .O(N__36509),
            .I(N__36506));
    Span4Mux_v I__7555 (
            .O(N__36506),
            .I(N__36503));
    Odrv4 I__7554 (
            .O(N__36503),
            .I(\current_shift_inst.control_inputZ0Z_3 ));
    InMux I__7553 (
            .O(N__36500),
            .I(\current_shift_inst.control_input_1_cry_2 ));
    InMux I__7552 (
            .O(N__36497),
            .I(N__36494));
    LocalMux I__7551 (
            .O(N__36494),
            .I(N__36491));
    Span4Mux_h I__7550 (
            .O(N__36491),
            .I(N__36488));
    Odrv4 I__7549 (
            .O(N__36488),
            .I(\current_shift_inst.control_inputZ0Z_4 ));
    InMux I__7548 (
            .O(N__36485),
            .I(\current_shift_inst.control_input_1_cry_3 ));
    InMux I__7547 (
            .O(N__36482),
            .I(N__36479));
    LocalMux I__7546 (
            .O(N__36479),
            .I(N__36476));
    Span4Mux_v I__7545 (
            .O(N__36476),
            .I(N__36473));
    Odrv4 I__7544 (
            .O(N__36473),
            .I(\current_shift_inst.control_inputZ0Z_5 ));
    InMux I__7543 (
            .O(N__36470),
            .I(\current_shift_inst.control_input_1_cry_4 ));
    InMux I__7542 (
            .O(N__36467),
            .I(N__36464));
    LocalMux I__7541 (
            .O(N__36464),
            .I(N__36461));
    Span4Mux_h I__7540 (
            .O(N__36461),
            .I(N__36458));
    Odrv4 I__7539 (
            .O(N__36458),
            .I(\current_shift_inst.control_inputZ0Z_6 ));
    InMux I__7538 (
            .O(N__36455),
            .I(\current_shift_inst.control_input_1_cry_5 ));
    InMux I__7537 (
            .O(N__36452),
            .I(N__36449));
    LocalMux I__7536 (
            .O(N__36449),
            .I(N__36446));
    Span4Mux_v I__7535 (
            .O(N__36446),
            .I(N__36443));
    Odrv4 I__7534 (
            .O(N__36443),
            .I(\current_shift_inst.control_inputZ0Z_7 ));
    InMux I__7533 (
            .O(N__36440),
            .I(\current_shift_inst.control_input_1_cry_6 ));
    InMux I__7532 (
            .O(N__36437),
            .I(N__36434));
    LocalMux I__7531 (
            .O(N__36434),
            .I(N__36431));
    Span4Mux_h I__7530 (
            .O(N__36431),
            .I(N__36428));
    Odrv4 I__7529 (
            .O(N__36428),
            .I(\current_shift_inst.control_inputZ0Z_8 ));
    InMux I__7528 (
            .O(N__36425),
            .I(bfn_15_17_0_));
    InMux I__7527 (
            .O(N__36422),
            .I(N__36419));
    LocalMux I__7526 (
            .O(N__36419),
            .I(N__36416));
    Span4Mux_v I__7525 (
            .O(N__36416),
            .I(N__36413));
    Odrv4 I__7524 (
            .O(N__36413),
            .I(\current_shift_inst.control_inputZ0Z_9 ));
    InMux I__7523 (
            .O(N__36410),
            .I(\current_shift_inst.control_input_1_cry_8 ));
    InMux I__7522 (
            .O(N__36407),
            .I(N__36404));
    LocalMux I__7521 (
            .O(N__36404),
            .I(N__36401));
    Span4Mux_v I__7520 (
            .O(N__36401),
            .I(N__36398));
    Odrv4 I__7519 (
            .O(N__36398),
            .I(\current_shift_inst.control_inputZ0Z_10 ));
    InMux I__7518 (
            .O(N__36395),
            .I(\current_shift_inst.control_input_1_cry_9 ));
    InMux I__7517 (
            .O(N__36392),
            .I(N__36388));
    InMux I__7516 (
            .O(N__36391),
            .I(N__36385));
    LocalMux I__7515 (
            .O(N__36388),
            .I(N__36382));
    LocalMux I__7514 (
            .O(N__36385),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv12 I__7513 (
            .O(N__36382),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__7512 (
            .O(N__36377),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__7511 (
            .O(N__36374),
            .I(N__36370));
    InMux I__7510 (
            .O(N__36373),
            .I(N__36367));
    LocalMux I__7509 (
            .O(N__36370),
            .I(N__36364));
    LocalMux I__7508 (
            .O(N__36367),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__7507 (
            .O(N__36364),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__7506 (
            .O(N__36359),
            .I(bfn_15_15_0_));
    InMux I__7505 (
            .O(N__36356),
            .I(N__36352));
    InMux I__7504 (
            .O(N__36355),
            .I(N__36349));
    LocalMux I__7503 (
            .O(N__36352),
            .I(N__36346));
    LocalMux I__7502 (
            .O(N__36349),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__7501 (
            .O(N__36346),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__7500 (
            .O(N__36341),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ));
    InMux I__7499 (
            .O(N__36338),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ));
    InMux I__7498 (
            .O(N__36335),
            .I(N__36331));
    InMux I__7497 (
            .O(N__36334),
            .I(N__36328));
    LocalMux I__7496 (
            .O(N__36331),
            .I(N__36325));
    LocalMux I__7495 (
            .O(N__36328),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__7494 (
            .O(N__36325),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__7493 (
            .O(N__36320),
            .I(N__36317));
    LocalMux I__7492 (
            .O(N__36317),
            .I(N__36314));
    Span12Mux_v I__7491 (
            .O(N__36314),
            .I(N__36311));
    Odrv12 I__7490 (
            .O(N__36311),
            .I(\phase_controller_inst1.stoper_hc.un1_start_latched2_0 ));
    InMux I__7489 (
            .O(N__36308),
            .I(N__36305));
    LocalMux I__7488 (
            .O(N__36305),
            .I(N__36302));
    Span4Mux_v I__7487 (
            .O(N__36302),
            .I(N__36297));
    InMux I__7486 (
            .O(N__36301),
            .I(N__36294));
    CascadeMux I__7485 (
            .O(N__36300),
            .I(N__36290));
    Span4Mux_h I__7484 (
            .O(N__36297),
            .I(N__36285));
    LocalMux I__7483 (
            .O(N__36294),
            .I(N__36285));
    CascadeMux I__7482 (
            .O(N__36293),
            .I(N__36281));
    InMux I__7481 (
            .O(N__36290),
            .I(N__36276));
    Span4Mux_h I__7480 (
            .O(N__36285),
            .I(N__36273));
    InMux I__7479 (
            .O(N__36284),
            .I(N__36270));
    InMux I__7478 (
            .O(N__36281),
            .I(N__36263));
    InMux I__7477 (
            .O(N__36280),
            .I(N__36263));
    InMux I__7476 (
            .O(N__36279),
            .I(N__36263));
    LocalMux I__7475 (
            .O(N__36276),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    Odrv4 I__7474 (
            .O(N__36273),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    LocalMux I__7473 (
            .O(N__36270),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    LocalMux I__7472 (
            .O(N__36263),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    InMux I__7471 (
            .O(N__36254),
            .I(N__36248));
    InMux I__7470 (
            .O(N__36253),
            .I(N__36245));
    InMux I__7469 (
            .O(N__36252),
            .I(N__36242));
    CascadeMux I__7468 (
            .O(N__36251),
            .I(N__36236));
    LocalMux I__7467 (
            .O(N__36248),
            .I(N__36233));
    LocalMux I__7466 (
            .O(N__36245),
            .I(N__36228));
    LocalMux I__7465 (
            .O(N__36242),
            .I(N__36228));
    InMux I__7464 (
            .O(N__36241),
            .I(N__36221));
    InMux I__7463 (
            .O(N__36240),
            .I(N__36221));
    InMux I__7462 (
            .O(N__36239),
            .I(N__36221));
    InMux I__7461 (
            .O(N__36236),
            .I(N__36217));
    Span4Mux_v I__7460 (
            .O(N__36233),
            .I(N__36214));
    Sp12to4 I__7459 (
            .O(N__36228),
            .I(N__36209));
    LocalMux I__7458 (
            .O(N__36221),
            .I(N__36209));
    InMux I__7457 (
            .O(N__36220),
            .I(N__36206));
    LocalMux I__7456 (
            .O(N__36217),
            .I(N__36203));
    Sp12to4 I__7455 (
            .O(N__36214),
            .I(N__36198));
    Span12Mux_v I__7454 (
            .O(N__36209),
            .I(N__36198));
    LocalMux I__7453 (
            .O(N__36206),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__7452 (
            .O(N__36203),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv12 I__7451 (
            .O(N__36198),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    InMux I__7450 (
            .O(N__36191),
            .I(N__36186));
    InMux I__7449 (
            .O(N__36190),
            .I(N__36181));
    InMux I__7448 (
            .O(N__36189),
            .I(N__36181));
    LocalMux I__7447 (
            .O(N__36186),
            .I(N__36177));
    LocalMux I__7446 (
            .O(N__36181),
            .I(N__36174));
    InMux I__7445 (
            .O(N__36180),
            .I(N__36171));
    Span4Mux_v I__7444 (
            .O(N__36177),
            .I(N__36166));
    Span4Mux_h I__7443 (
            .O(N__36174),
            .I(N__36166));
    LocalMux I__7442 (
            .O(N__36171),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv4 I__7441 (
            .O(N__36166),
            .I(\phase_controller_inst1.hc_time_passed ));
    InMux I__7440 (
            .O(N__36161),
            .I(N__36158));
    LocalMux I__7439 (
            .O(N__36158),
            .I(N__36154));
    InMux I__7438 (
            .O(N__36157),
            .I(N__36151));
    Span4Mux_v I__7437 (
            .O(N__36154),
            .I(N__36146));
    LocalMux I__7436 (
            .O(N__36151),
            .I(N__36146));
    Span4Mux_v I__7435 (
            .O(N__36146),
            .I(N__36143));
    Span4Mux_h I__7434 (
            .O(N__36143),
            .I(N__36140));
    Odrv4 I__7433 (
            .O(N__36140),
            .I(\current_shift_inst.control_inputZ0Z_0 ));
    InMux I__7432 (
            .O(N__36137),
            .I(N__36134));
    LocalMux I__7431 (
            .O(N__36134),
            .I(N__36131));
    Odrv12 I__7430 (
            .O(N__36131),
            .I(\current_shift_inst.control_inputZ0Z_1 ));
    InMux I__7429 (
            .O(N__36128),
            .I(\current_shift_inst.control_input_1_cry_0 ));
    InMux I__7428 (
            .O(N__36125),
            .I(N__36122));
    LocalMux I__7427 (
            .O(N__36122),
            .I(N__36119));
    Span4Mux_h I__7426 (
            .O(N__36119),
            .I(N__36116));
    Odrv4 I__7425 (
            .O(N__36116),
            .I(\current_shift_inst.control_inputZ0Z_2 ));
    InMux I__7424 (
            .O(N__36113),
            .I(\current_shift_inst.control_input_1_cry_1 ));
    InMux I__7423 (
            .O(N__36110),
            .I(N__36106));
    InMux I__7422 (
            .O(N__36109),
            .I(N__36103));
    LocalMux I__7421 (
            .O(N__36106),
            .I(N__36100));
    LocalMux I__7420 (
            .O(N__36103),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv12 I__7419 (
            .O(N__36100),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__7418 (
            .O(N__36095),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__7417 (
            .O(N__36092),
            .I(N__36088));
    InMux I__7416 (
            .O(N__36091),
            .I(N__36085));
    LocalMux I__7415 (
            .O(N__36088),
            .I(N__36082));
    LocalMux I__7414 (
            .O(N__36085),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    Odrv12 I__7413 (
            .O(N__36082),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__7412 (
            .O(N__36077),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__7411 (
            .O(N__36074),
            .I(N__36070));
    InMux I__7410 (
            .O(N__36073),
            .I(N__36067));
    LocalMux I__7409 (
            .O(N__36070),
            .I(N__36064));
    LocalMux I__7408 (
            .O(N__36067),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__7407 (
            .O(N__36064),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__7406 (
            .O(N__36059),
            .I(bfn_15_14_0_));
    InMux I__7405 (
            .O(N__36056),
            .I(N__36052));
    InMux I__7404 (
            .O(N__36055),
            .I(N__36049));
    LocalMux I__7403 (
            .O(N__36052),
            .I(N__36046));
    LocalMux I__7402 (
            .O(N__36049),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv4 I__7401 (
            .O(N__36046),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__7400 (
            .O(N__36041),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__7399 (
            .O(N__36038),
            .I(N__36034));
    InMux I__7398 (
            .O(N__36037),
            .I(N__36031));
    LocalMux I__7397 (
            .O(N__36034),
            .I(N__36028));
    LocalMux I__7396 (
            .O(N__36031),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv4 I__7395 (
            .O(N__36028),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__7394 (
            .O(N__36023),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__7393 (
            .O(N__36020),
            .I(N__36016));
    InMux I__7392 (
            .O(N__36019),
            .I(N__36013));
    LocalMux I__7391 (
            .O(N__36016),
            .I(N__36010));
    LocalMux I__7390 (
            .O(N__36013),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__7389 (
            .O(N__36010),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__7388 (
            .O(N__36005),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__7387 (
            .O(N__36002),
            .I(N__35999));
    LocalMux I__7386 (
            .O(N__35999),
            .I(N__35995));
    InMux I__7385 (
            .O(N__35998),
            .I(N__35992));
    Span4Mux_v I__7384 (
            .O(N__35995),
            .I(N__35989));
    LocalMux I__7383 (
            .O(N__35992),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__7382 (
            .O(N__35989),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__7381 (
            .O(N__35984),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__7380 (
            .O(N__35981),
            .I(N__35977));
    InMux I__7379 (
            .O(N__35980),
            .I(N__35974));
    LocalMux I__7378 (
            .O(N__35977),
            .I(N__35971));
    LocalMux I__7377 (
            .O(N__35974),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__7376 (
            .O(N__35971),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__7375 (
            .O(N__35966),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__7374 (
            .O(N__35963),
            .I(N__35960));
    LocalMux I__7373 (
            .O(N__35960),
            .I(N__35956));
    InMux I__7372 (
            .O(N__35959),
            .I(N__35953));
    Span4Mux_v I__7371 (
            .O(N__35956),
            .I(N__35950));
    LocalMux I__7370 (
            .O(N__35953),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv4 I__7369 (
            .O(N__35950),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__7368 (
            .O(N__35945),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ));
    InMux I__7367 (
            .O(N__35942),
            .I(N__35939));
    LocalMux I__7366 (
            .O(N__35939),
            .I(N__35936));
    Span4Mux_h I__7365 (
            .O(N__35936),
            .I(N__35933));
    Odrv4 I__7364 (
            .O(N__35933),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ));
    InMux I__7363 (
            .O(N__35930),
            .I(N__35923));
    InMux I__7362 (
            .O(N__35929),
            .I(N__35919));
    InMux I__7361 (
            .O(N__35928),
            .I(N__35914));
    InMux I__7360 (
            .O(N__35927),
            .I(N__35911));
    InMux I__7359 (
            .O(N__35926),
            .I(N__35908));
    LocalMux I__7358 (
            .O(N__35923),
            .I(N__35905));
    CascadeMux I__7357 (
            .O(N__35922),
            .I(N__35902));
    LocalMux I__7356 (
            .O(N__35919),
            .I(N__35899));
    InMux I__7355 (
            .O(N__35918),
            .I(N__35894));
    InMux I__7354 (
            .O(N__35917),
            .I(N__35894));
    LocalMux I__7353 (
            .O(N__35914),
            .I(N__35891));
    LocalMux I__7352 (
            .O(N__35911),
            .I(N__35886));
    LocalMux I__7351 (
            .O(N__35908),
            .I(N__35886));
    Span4Mux_v I__7350 (
            .O(N__35905),
            .I(N__35883));
    InMux I__7349 (
            .O(N__35902),
            .I(N__35880));
    Span4Mux_v I__7348 (
            .O(N__35899),
            .I(N__35877));
    LocalMux I__7347 (
            .O(N__35894),
            .I(N__35874));
    Span4Mux_v I__7346 (
            .O(N__35891),
            .I(N__35867));
    Span4Mux_v I__7345 (
            .O(N__35886),
            .I(N__35867));
    Span4Mux_h I__7344 (
            .O(N__35883),
            .I(N__35867));
    LocalMux I__7343 (
            .O(N__35880),
            .I(N__35862));
    Span4Mux_h I__7342 (
            .O(N__35877),
            .I(N__35862));
    Odrv12 I__7341 (
            .O(N__35874),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5 ));
    Odrv4 I__7340 (
            .O(N__35867),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5 ));
    Odrv4 I__7339 (
            .O(N__35862),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5 ));
    CascadeMux I__7338 (
            .O(N__35855),
            .I(N__35852));
    InMux I__7337 (
            .O(N__35852),
            .I(N__35849));
    LocalMux I__7336 (
            .O(N__35849),
            .I(N__35846));
    Span4Mux_h I__7335 (
            .O(N__35846),
            .I(N__35840));
    InMux I__7334 (
            .O(N__35845),
            .I(N__35837));
    InMux I__7333 (
            .O(N__35844),
            .I(N__35834));
    InMux I__7332 (
            .O(N__35843),
            .I(N__35831));
    Odrv4 I__7331 (
            .O(N__35840),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto9 ));
    LocalMux I__7330 (
            .O(N__35837),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto9 ));
    LocalMux I__7329 (
            .O(N__35834),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto9 ));
    LocalMux I__7328 (
            .O(N__35831),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto9 ));
    InMux I__7327 (
            .O(N__35822),
            .I(N__35817));
    InMux I__7326 (
            .O(N__35821),
            .I(N__35810));
    InMux I__7325 (
            .O(N__35820),
            .I(N__35810));
    LocalMux I__7324 (
            .O(N__35817),
            .I(N__35807));
    CascadeMux I__7323 (
            .O(N__35816),
            .I(N__35804));
    InMux I__7322 (
            .O(N__35815),
            .I(N__35801));
    LocalMux I__7321 (
            .O(N__35810),
            .I(N__35798));
    Span4Mux_h I__7320 (
            .O(N__35807),
            .I(N__35795));
    InMux I__7319 (
            .O(N__35804),
            .I(N__35792));
    LocalMux I__7318 (
            .O(N__35801),
            .I(N__35785));
    Span4Mux_v I__7317 (
            .O(N__35798),
            .I(N__35785));
    Span4Mux_h I__7316 (
            .O(N__35795),
            .I(N__35785));
    LocalMux I__7315 (
            .O(N__35792),
            .I(elapsed_time_ns_1_RNIL13KD1_0_9));
    Odrv4 I__7314 (
            .O(N__35785),
            .I(elapsed_time_ns_1_RNIL13KD1_0_9));
    InMux I__7313 (
            .O(N__35780),
            .I(N__35777));
    LocalMux I__7312 (
            .O(N__35777),
            .I(N__35774));
    Span4Mux_v I__7311 (
            .O(N__35774),
            .I(N__35771));
    Span4Mux_h I__7310 (
            .O(N__35771),
            .I(N__35768));
    Odrv4 I__7309 (
            .O(N__35768),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9 ));
    InMux I__7308 (
            .O(N__35765),
            .I(N__35762));
    LocalMux I__7307 (
            .O(N__35762),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ));
    CascadeMux I__7306 (
            .O(N__35759),
            .I(N__35756));
    InMux I__7305 (
            .O(N__35756),
            .I(N__35752));
    InMux I__7304 (
            .O(N__35755),
            .I(N__35749));
    LocalMux I__7303 (
            .O(N__35752),
            .I(N__35746));
    LocalMux I__7302 (
            .O(N__35749),
            .I(N__35743));
    Span4Mux_v I__7301 (
            .O(N__35746),
            .I(N__35739));
    Span4Mux_h I__7300 (
            .O(N__35743),
            .I(N__35736));
    CascadeMux I__7299 (
            .O(N__35742),
            .I(N__35733));
    Span4Mux_h I__7298 (
            .O(N__35739),
            .I(N__35728));
    Span4Mux_v I__7297 (
            .O(N__35736),
            .I(N__35728));
    InMux I__7296 (
            .O(N__35733),
            .I(N__35725));
    Span4Mux_h I__7295 (
            .O(N__35728),
            .I(N__35722));
    LocalMux I__7294 (
            .O(N__35725),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__7293 (
            .O(N__35722),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__7292 (
            .O(N__35717),
            .I(N__35713));
    InMux I__7291 (
            .O(N__35716),
            .I(N__35710));
    LocalMux I__7290 (
            .O(N__35713),
            .I(N__35707));
    LocalMux I__7289 (
            .O(N__35710),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    Odrv4 I__7288 (
            .O(N__35707),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__7287 (
            .O(N__35702),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ));
    CascadeMux I__7286 (
            .O(N__35699),
            .I(N__35696));
    InMux I__7285 (
            .O(N__35696),
            .I(N__35693));
    LocalMux I__7284 (
            .O(N__35693),
            .I(N__35690));
    Odrv4 I__7283 (
            .O(N__35690),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNI2FGQZ0Z1 ));
    InMux I__7282 (
            .O(N__35687),
            .I(N__35683));
    InMux I__7281 (
            .O(N__35686),
            .I(N__35680));
    LocalMux I__7280 (
            .O(N__35683),
            .I(N__35677));
    LocalMux I__7279 (
            .O(N__35680),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    Odrv4 I__7278 (
            .O(N__35677),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__7277 (
            .O(N__35672),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__7276 (
            .O(N__35669),
            .I(N__35665));
    InMux I__7275 (
            .O(N__35668),
            .I(N__35662));
    LocalMux I__7274 (
            .O(N__35665),
            .I(N__35659));
    LocalMux I__7273 (
            .O(N__35662),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    Odrv4 I__7272 (
            .O(N__35659),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__7271 (
            .O(N__35654),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__7270 (
            .O(N__35651),
            .I(N__35647));
    InMux I__7269 (
            .O(N__35650),
            .I(N__35644));
    LocalMux I__7268 (
            .O(N__35647),
            .I(N__35641));
    LocalMux I__7267 (
            .O(N__35644),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    Odrv4 I__7266 (
            .O(N__35641),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__7265 (
            .O(N__35636),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ));
    InMux I__7264 (
            .O(N__35633),
            .I(N__35629));
    InMux I__7263 (
            .O(N__35632),
            .I(N__35626));
    LocalMux I__7262 (
            .O(N__35629),
            .I(N__35623));
    LocalMux I__7261 (
            .O(N__35626),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    Odrv4 I__7260 (
            .O(N__35623),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__7259 (
            .O(N__35618),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ));
    CascadeMux I__7258 (
            .O(N__35615),
            .I(N__35612));
    InMux I__7257 (
            .O(N__35612),
            .I(N__35609));
    LocalMux I__7256 (
            .O(N__35609),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ));
    CascadeMux I__7255 (
            .O(N__35606),
            .I(N__35603));
    InMux I__7254 (
            .O(N__35603),
            .I(N__35600));
    LocalMux I__7253 (
            .O(N__35600),
            .I(N__35597));
    Odrv4 I__7252 (
            .O(N__35597),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ));
    CascadeMux I__7251 (
            .O(N__35594),
            .I(N__35591));
    InMux I__7250 (
            .O(N__35591),
            .I(N__35588));
    LocalMux I__7249 (
            .O(N__35588),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ));
    CascadeMux I__7248 (
            .O(N__35585),
            .I(N__35582));
    InMux I__7247 (
            .O(N__35582),
            .I(N__35579));
    LocalMux I__7246 (
            .O(N__35579),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_16 ));
    CascadeMux I__7245 (
            .O(N__35576),
            .I(N__35573));
    InMux I__7244 (
            .O(N__35573),
            .I(N__35570));
    LocalMux I__7243 (
            .O(N__35570),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_17 ));
    CascadeMux I__7242 (
            .O(N__35567),
            .I(N__35564));
    InMux I__7241 (
            .O(N__35564),
            .I(N__35561));
    LocalMux I__7240 (
            .O(N__35561),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_18 ));
    CascadeMux I__7239 (
            .O(N__35558),
            .I(N__35555));
    InMux I__7238 (
            .O(N__35555),
            .I(N__35552));
    LocalMux I__7237 (
            .O(N__35552),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_19 ));
    InMux I__7236 (
            .O(N__35549),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_19 ));
    InMux I__7235 (
            .O(N__35546),
            .I(N__35543));
    LocalMux I__7234 (
            .O(N__35543),
            .I(N__35540));
    Span4Mux_h I__7233 (
            .O(N__35540),
            .I(N__35536));
    InMux I__7232 (
            .O(N__35539),
            .I(N__35533));
    Odrv4 I__7231 (
            .O(N__35536),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_CO ));
    LocalMux I__7230 (
            .O(N__35533),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_CO ));
    InMux I__7229 (
            .O(N__35528),
            .I(N__35525));
    LocalMux I__7228 (
            .O(N__35525),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ));
    CascadeMux I__7227 (
            .O(N__35522),
            .I(N__35519));
    InMux I__7226 (
            .O(N__35519),
            .I(N__35516));
    LocalMux I__7225 (
            .O(N__35516),
            .I(N__35513));
    Odrv4 I__7224 (
            .O(N__35513),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ));
    CascadeMux I__7223 (
            .O(N__35510),
            .I(N__35507));
    InMux I__7222 (
            .O(N__35507),
            .I(N__35504));
    LocalMux I__7221 (
            .O(N__35504),
            .I(N__35501));
    Odrv4 I__7220 (
            .O(N__35501),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ));
    CascadeMux I__7219 (
            .O(N__35498),
            .I(N__35495));
    InMux I__7218 (
            .O(N__35495),
            .I(N__35492));
    LocalMux I__7217 (
            .O(N__35492),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ));
    CascadeMux I__7216 (
            .O(N__35489),
            .I(N__35486));
    InMux I__7215 (
            .O(N__35486),
            .I(N__35483));
    LocalMux I__7214 (
            .O(N__35483),
            .I(N__35480));
    Odrv4 I__7213 (
            .O(N__35480),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ));
    CascadeMux I__7212 (
            .O(N__35477),
            .I(N__35474));
    InMux I__7211 (
            .O(N__35474),
            .I(N__35471));
    LocalMux I__7210 (
            .O(N__35471),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ));
    CascadeMux I__7209 (
            .O(N__35468),
            .I(N__35465));
    InMux I__7208 (
            .O(N__35465),
            .I(N__35462));
    LocalMux I__7207 (
            .O(N__35462),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ));
    InMux I__7206 (
            .O(N__35459),
            .I(N__35456));
    LocalMux I__7205 (
            .O(N__35456),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ));
    InMux I__7204 (
            .O(N__35453),
            .I(N__35450));
    LocalMux I__7203 (
            .O(N__35450),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ));
    InMux I__7202 (
            .O(N__35447),
            .I(N__35443));
    InMux I__7201 (
            .O(N__35446),
            .I(N__35440));
    LocalMux I__7200 (
            .O(N__35443),
            .I(elapsed_time_ns_1_RNI0GIF91_0_26));
    LocalMux I__7199 (
            .O(N__35440),
            .I(elapsed_time_ns_1_RNI0GIF91_0_26));
    CascadeMux I__7198 (
            .O(N__35435),
            .I(N__35432));
    InMux I__7197 (
            .O(N__35432),
            .I(N__35429));
    LocalMux I__7196 (
            .O(N__35429),
            .I(N__35426));
    Span4Mux_h I__7195 (
            .O(N__35426),
            .I(N__35422));
    InMux I__7194 (
            .O(N__35425),
            .I(N__35419));
    Odrv4 I__7193 (
            .O(N__35422),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    LocalMux I__7192 (
            .O(N__35419),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__7191 (
            .O(N__35414),
            .I(N__35408));
    InMux I__7190 (
            .O(N__35413),
            .I(N__35408));
    LocalMux I__7189 (
            .O(N__35408),
            .I(elapsed_time_ns_1_RNI2IIF91_0_28));
    CascadeMux I__7188 (
            .O(N__35405),
            .I(N__35402));
    InMux I__7187 (
            .O(N__35402),
            .I(N__35399));
    LocalMux I__7186 (
            .O(N__35399),
            .I(N__35395));
    InMux I__7185 (
            .O(N__35398),
            .I(N__35392));
    Odrv4 I__7184 (
            .O(N__35395),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    LocalMux I__7183 (
            .O(N__35392),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    InMux I__7182 (
            .O(N__35387),
            .I(N__35383));
    InMux I__7181 (
            .O(N__35386),
            .I(N__35379));
    LocalMux I__7180 (
            .O(N__35383),
            .I(N__35376));
    InMux I__7179 (
            .O(N__35382),
            .I(N__35373));
    LocalMux I__7178 (
            .O(N__35379),
            .I(N__35370));
    Odrv4 I__7177 (
            .O(N__35376),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    LocalMux I__7176 (
            .O(N__35373),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    Odrv4 I__7175 (
            .O(N__35370),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    CascadeMux I__7174 (
            .O(N__35363),
            .I(N__35360));
    InMux I__7173 (
            .O(N__35360),
            .I(N__35357));
    LocalMux I__7172 (
            .O(N__35357),
            .I(N__35353));
    InMux I__7171 (
            .O(N__35356),
            .I(N__35350));
    Span4Mux_v I__7170 (
            .O(N__35353),
            .I(N__35347));
    LocalMux I__7169 (
            .O(N__35350),
            .I(N__35344));
    Odrv4 I__7168 (
            .O(N__35347),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    Odrv4 I__7167 (
            .O(N__35344),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    InMux I__7166 (
            .O(N__35339),
            .I(N__35336));
    LocalMux I__7165 (
            .O(N__35336),
            .I(N__35332));
    CascadeMux I__7164 (
            .O(N__35335),
            .I(N__35329));
    Span4Mux_v I__7163 (
            .O(N__35332),
            .I(N__35326));
    InMux I__7162 (
            .O(N__35329),
            .I(N__35323));
    Odrv4 I__7161 (
            .O(N__35326),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    LocalMux I__7160 (
            .O(N__35323),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    CascadeMux I__7159 (
            .O(N__35318),
            .I(N__35315));
    InMux I__7158 (
            .O(N__35315),
            .I(N__35312));
    LocalMux I__7157 (
            .O(N__35312),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ));
    CascadeMux I__7156 (
            .O(N__35309),
            .I(N__35306));
    InMux I__7155 (
            .O(N__35306),
            .I(N__35303));
    LocalMux I__7154 (
            .O(N__35303),
            .I(N__35300));
    Odrv4 I__7153 (
            .O(N__35300),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ));
    CascadeMux I__7152 (
            .O(N__35297),
            .I(N__35294));
    InMux I__7151 (
            .O(N__35294),
            .I(N__35291));
    LocalMux I__7150 (
            .O(N__35291),
            .I(N__35288));
    Odrv4 I__7149 (
            .O(N__35288),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ));
    InMux I__7148 (
            .O(N__35285),
            .I(N__35282));
    LocalMux I__7147 (
            .O(N__35282),
            .I(N__35279));
    Span4Mux_v I__7146 (
            .O(N__35279),
            .I(N__35275));
    InMux I__7145 (
            .O(N__35278),
            .I(N__35272));
    Odrv4 I__7144 (
            .O(N__35275),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    LocalMux I__7143 (
            .O(N__35272),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    CascadeMux I__7142 (
            .O(N__35267),
            .I(elapsed_time_ns_1_RNISAHF91_0_13_cascade_));
    InMux I__7141 (
            .O(N__35264),
            .I(N__35261));
    LocalMux I__7140 (
            .O(N__35261),
            .I(N__35258));
    Span4Mux_h I__7139 (
            .O(N__35258),
            .I(N__35254));
    InMux I__7138 (
            .O(N__35257),
            .I(N__35251));
    Odrv4 I__7137 (
            .O(N__35254),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    LocalMux I__7136 (
            .O(N__35251),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__7135 (
            .O(N__35246),
            .I(N__35243));
    LocalMux I__7134 (
            .O(N__35243),
            .I(N__35240));
    Span4Mux_h I__7133 (
            .O(N__35240),
            .I(N__35236));
    InMux I__7132 (
            .O(N__35239),
            .I(N__35233));
    Odrv4 I__7131 (
            .O(N__35236),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    LocalMux I__7130 (
            .O(N__35233),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__7129 (
            .O(N__35228),
            .I(N__35225));
    LocalMux I__7128 (
            .O(N__35225),
            .I(elapsed_time_ns_1_RNIVEIF91_0_25));
    InMux I__7127 (
            .O(N__35222),
            .I(N__35218));
    InMux I__7126 (
            .O(N__35221),
            .I(N__35215));
    LocalMux I__7125 (
            .O(N__35218),
            .I(elapsed_time_ns_1_RNI1HIF91_0_27));
    LocalMux I__7124 (
            .O(N__35215),
            .I(elapsed_time_ns_1_RNI1HIF91_0_27));
    CascadeMux I__7123 (
            .O(N__35210),
            .I(elapsed_time_ns_1_RNIVEIF91_0_25_cascade_));
    InMux I__7122 (
            .O(N__35207),
            .I(N__35204));
    LocalMux I__7121 (
            .O(N__35204),
            .I(N__35201));
    Span4Mux_h I__7120 (
            .O(N__35201),
            .I(N__35197));
    InMux I__7119 (
            .O(N__35200),
            .I(N__35194));
    Span4Mux_v I__7118 (
            .O(N__35197),
            .I(N__35189));
    LocalMux I__7117 (
            .O(N__35194),
            .I(N__35186));
    InMux I__7116 (
            .O(N__35193),
            .I(N__35181));
    InMux I__7115 (
            .O(N__35192),
            .I(N__35181));
    Odrv4 I__7114 (
            .O(N__35189),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ));
    Odrv4 I__7113 (
            .O(N__35186),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ));
    LocalMux I__7112 (
            .O(N__35181),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ));
    InMux I__7111 (
            .O(N__35174),
            .I(N__35171));
    LocalMux I__7110 (
            .O(N__35171),
            .I(N__35168));
    Span4Mux_h I__7109 (
            .O(N__35168),
            .I(N__35165));
    Span4Mux_v I__7108 (
            .O(N__35165),
            .I(N__35161));
    InMux I__7107 (
            .O(N__35164),
            .I(N__35158));
    Odrv4 I__7106 (
            .O(N__35161),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    LocalMux I__7105 (
            .O(N__35158),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    CascadeMux I__7104 (
            .O(N__35153),
            .I(N__35150));
    InMux I__7103 (
            .O(N__35150),
            .I(N__35147));
    LocalMux I__7102 (
            .O(N__35147),
            .I(N__35143));
    InMux I__7101 (
            .O(N__35146),
            .I(N__35140));
    Odrv12 I__7100 (
            .O(N__35143),
            .I(\delay_measurement_inst.delay_tr_timer.N_381 ));
    LocalMux I__7099 (
            .O(N__35140),
            .I(\delay_measurement_inst.delay_tr_timer.N_381 ));
    InMux I__7098 (
            .O(N__35135),
            .I(N__35132));
    LocalMux I__7097 (
            .O(N__35132),
            .I(\delay_measurement_inst.delay_tr_timer.N_358 ));
    CascadeMux I__7096 (
            .O(N__35129),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_ ));
    InMux I__7095 (
            .O(N__35126),
            .I(N__35123));
    LocalMux I__7094 (
            .O(N__35123),
            .I(N__35120));
    Span4Mux_v I__7093 (
            .O(N__35120),
            .I(N__35116));
    InMux I__7092 (
            .O(N__35119),
            .I(N__35113));
    Odrv4 I__7091 (
            .O(N__35116),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    LocalMux I__7090 (
            .O(N__35113),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    InMux I__7089 (
            .O(N__35108),
            .I(N__35104));
    CascadeMux I__7088 (
            .O(N__35107),
            .I(N__35100));
    LocalMux I__7087 (
            .O(N__35104),
            .I(N__35097));
    InMux I__7086 (
            .O(N__35103),
            .I(N__35094));
    InMux I__7085 (
            .O(N__35100),
            .I(N__35091));
    Span4Mux_h I__7084 (
            .O(N__35097),
            .I(N__35088));
    LocalMux I__7083 (
            .O(N__35094),
            .I(N__35083));
    LocalMux I__7082 (
            .O(N__35091),
            .I(N__35083));
    Odrv4 I__7081 (
            .O(N__35088),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    Odrv4 I__7080 (
            .O(N__35083),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    CascadeMux I__7079 (
            .O(N__35078),
            .I(elapsed_time_ns_1_RNIIJ4DM1_0_19_cascade_));
    InMux I__7078 (
            .O(N__35075),
            .I(N__35072));
    LocalMux I__7077 (
            .O(N__35072),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19 ));
    InMux I__7076 (
            .O(N__35069),
            .I(bfn_14_21_0_));
    InMux I__7075 (
            .O(N__35066),
            .I(\current_shift_inst.un38_control_input_cry_24_s1 ));
    CascadeMux I__7074 (
            .O(N__35063),
            .I(N__35060));
    InMux I__7073 (
            .O(N__35060),
            .I(N__35057));
    LocalMux I__7072 (
            .O(N__35057),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ));
    InMux I__7071 (
            .O(N__35054),
            .I(\current_shift_inst.un38_control_input_cry_25_s1 ));
    InMux I__7070 (
            .O(N__35051),
            .I(\current_shift_inst.un38_control_input_cry_26_s1 ));
    CascadeMux I__7069 (
            .O(N__35048),
            .I(N__35045));
    InMux I__7068 (
            .O(N__35045),
            .I(N__35042));
    LocalMux I__7067 (
            .O(N__35042),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ));
    InMux I__7066 (
            .O(N__35039),
            .I(\current_shift_inst.un38_control_input_cry_27_s1 ));
    InMux I__7065 (
            .O(N__35036),
            .I(\current_shift_inst.un38_control_input_cry_28_s1 ));
    InMux I__7064 (
            .O(N__35033),
            .I(\current_shift_inst.un38_control_input_cry_29_s1 ));
    InMux I__7063 (
            .O(N__35030),
            .I(\current_shift_inst.un38_control_input_cry_30_s1 ));
    InMux I__7062 (
            .O(N__35027),
            .I(N__35024));
    LocalMux I__7061 (
            .O(N__35024),
            .I(N__35021));
    Odrv12 I__7060 (
            .O(N__35021),
            .I(\current_shift_inst.un38_control_input_0_s1_31 ));
    CascadeMux I__7059 (
            .O(N__35018),
            .I(N__35015));
    InMux I__7058 (
            .O(N__35015),
            .I(N__35012));
    LocalMux I__7057 (
            .O(N__35012),
            .I(N__35009));
    Span4Mux_h I__7056 (
            .O(N__35009),
            .I(N__35006));
    Odrv4 I__7055 (
            .O(N__35006),
            .I(\current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ));
    InMux I__7054 (
            .O(N__35003),
            .I(\current_shift_inst.un38_control_input_cry_19_s1 ));
    CascadeMux I__7053 (
            .O(N__35000),
            .I(N__34997));
    InMux I__7052 (
            .O(N__34997),
            .I(N__34994));
    LocalMux I__7051 (
            .O(N__34994),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ));
    InMux I__7050 (
            .O(N__34991),
            .I(\current_shift_inst.un38_control_input_cry_20_s1 ));
    InMux I__7049 (
            .O(N__34988),
            .I(\current_shift_inst.un38_control_input_cry_21_s1 ));
    InMux I__7048 (
            .O(N__34985),
            .I(\current_shift_inst.un38_control_input_cry_22_s1 ));
    InMux I__7047 (
            .O(N__34982),
            .I(\current_shift_inst.un38_control_input_cry_28_s0 ));
    InMux I__7046 (
            .O(N__34979),
            .I(\current_shift_inst.un38_control_input_cry_29_s0 ));
    InMux I__7045 (
            .O(N__34976),
            .I(N__34973));
    LocalMux I__7044 (
            .O(N__34973),
            .I(N__34970));
    Odrv4 I__7043 (
            .O(N__34970),
            .I(\current_shift_inst.un38_control_input_axb_31_s0 ));
    InMux I__7042 (
            .O(N__34967),
            .I(\current_shift_inst.un38_control_input_cry_30_s0 ));
    InMux I__7041 (
            .O(N__34964),
            .I(N__34960));
    InMux I__7040 (
            .O(N__34963),
            .I(N__34957));
    LocalMux I__7039 (
            .O(N__34960),
            .I(N__34954));
    LocalMux I__7038 (
            .O(N__34957),
            .I(N__34951));
    Odrv4 I__7037 (
            .O(N__34954),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    Odrv4 I__7036 (
            .O(N__34951),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    InMux I__7035 (
            .O(N__34946),
            .I(N__34943));
    LocalMux I__7034 (
            .O(N__34943),
            .I(\current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ));
    InMux I__7033 (
            .O(N__34940),
            .I(\current_shift_inst.un38_control_input_cry_19_s0 ));
    InMux I__7032 (
            .O(N__34937),
            .I(N__34934));
    LocalMux I__7031 (
            .O(N__34934),
            .I(N__34931));
    Odrv4 I__7030 (
            .O(N__34931),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ));
    InMux I__7029 (
            .O(N__34928),
            .I(\current_shift_inst.un38_control_input_cry_20_s0 ));
    InMux I__7028 (
            .O(N__34925),
            .I(\current_shift_inst.un38_control_input_cry_21_s0 ));
    InMux I__7027 (
            .O(N__34922),
            .I(\current_shift_inst.un38_control_input_cry_22_s0 ));
    InMux I__7026 (
            .O(N__34919),
            .I(bfn_14_17_0_));
    InMux I__7025 (
            .O(N__34916),
            .I(N__34913));
    LocalMux I__7024 (
            .O(N__34913),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ));
    InMux I__7023 (
            .O(N__34910),
            .I(\current_shift_inst.un38_control_input_cry_24_s0 ));
    InMux I__7022 (
            .O(N__34907),
            .I(\current_shift_inst.un38_control_input_cry_25_s0 ));
    InMux I__7021 (
            .O(N__34904),
            .I(N__34901));
    LocalMux I__7020 (
            .O(N__34901),
            .I(N__34898));
    Odrv4 I__7019 (
            .O(N__34898),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ));
    InMux I__7018 (
            .O(N__34895),
            .I(\current_shift_inst.un38_control_input_cry_26_s0 ));
    CascadeMux I__7017 (
            .O(N__34892),
            .I(N__34889));
    InMux I__7016 (
            .O(N__34889),
            .I(N__34886));
    LocalMux I__7015 (
            .O(N__34886),
            .I(N__34883));
    Odrv4 I__7014 (
            .O(N__34883),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ));
    InMux I__7013 (
            .O(N__34880),
            .I(\current_shift_inst.un38_control_input_cry_27_s0 ));
    InMux I__7012 (
            .O(N__34877),
            .I(N__34874));
    LocalMux I__7011 (
            .O(N__34874),
            .I(\current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ));
    InMux I__7010 (
            .O(N__34871),
            .I(N__34868));
    LocalMux I__7009 (
            .O(N__34868),
            .I(\current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ));
    InMux I__7008 (
            .O(N__34865),
            .I(N__34862));
    LocalMux I__7007 (
            .O(N__34862),
            .I(\current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ));
    InMux I__7006 (
            .O(N__34859),
            .I(N__34856));
    LocalMux I__7005 (
            .O(N__34856),
            .I(N__34853));
    Odrv4 I__7004 (
            .O(N__34853),
            .I(\current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ));
    CascadeMux I__7003 (
            .O(N__34850),
            .I(N__34847));
    InMux I__7002 (
            .O(N__34847),
            .I(N__34844));
    LocalMux I__7001 (
            .O(N__34844),
            .I(\current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ));
    CascadeMux I__7000 (
            .O(N__34841),
            .I(N__34838));
    InMux I__6999 (
            .O(N__34838),
            .I(N__34835));
    LocalMux I__6998 (
            .O(N__34835),
            .I(\current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ));
    CascadeMux I__6997 (
            .O(N__34832),
            .I(\phase_controller_inst1.start_timer_tr_0_sqmuxa_cascade_ ));
    InMux I__6996 (
            .O(N__34829),
            .I(N__34822));
    InMux I__6995 (
            .O(N__34828),
            .I(N__34822));
    InMux I__6994 (
            .O(N__34827),
            .I(N__34819));
    LocalMux I__6993 (
            .O(N__34822),
            .I(N__34816));
    LocalMux I__6992 (
            .O(N__34819),
            .I(N__34813));
    Span4Mux_h I__6991 (
            .O(N__34816),
            .I(N__34809));
    Span4Mux_v I__6990 (
            .O(N__34813),
            .I(N__34806));
    InMux I__6989 (
            .O(N__34812),
            .I(N__34803));
    Span4Mux_v I__6988 (
            .O(N__34809),
            .I(N__34798));
    Span4Mux_h I__6987 (
            .O(N__34806),
            .I(N__34793));
    LocalMux I__6986 (
            .O(N__34803),
            .I(N__34793));
    InMux I__6985 (
            .O(N__34802),
            .I(N__34790));
    InMux I__6984 (
            .O(N__34801),
            .I(N__34787));
    Odrv4 I__6983 (
            .O(N__34798),
            .I(phase_controller_inst1_state_4));
    Odrv4 I__6982 (
            .O(N__34793),
            .I(phase_controller_inst1_state_4));
    LocalMux I__6981 (
            .O(N__34790),
            .I(phase_controller_inst1_state_4));
    LocalMux I__6980 (
            .O(N__34787),
            .I(phase_controller_inst1_state_4));
    CascadeMux I__6979 (
            .O(N__34778),
            .I(N__34775));
    InMux I__6978 (
            .O(N__34775),
            .I(N__34772));
    LocalMux I__6977 (
            .O(N__34772),
            .I(\phase_controller_inst2.stoper_tr.un1_start_latched2_0 ));
    InMux I__6976 (
            .O(N__34769),
            .I(N__34765));
    InMux I__6975 (
            .O(N__34768),
            .I(N__34762));
    LocalMux I__6974 (
            .O(N__34765),
            .I(N__34756));
    LocalMux I__6973 (
            .O(N__34762),
            .I(N__34756));
    InMux I__6972 (
            .O(N__34761),
            .I(N__34753));
    Span4Mux_v I__6971 (
            .O(N__34756),
            .I(N__34750));
    LocalMux I__6970 (
            .O(N__34753),
            .I(\phase_controller_inst2.tr_time_passed ));
    Odrv4 I__6969 (
            .O(N__34750),
            .I(\phase_controller_inst2.tr_time_passed ));
    CascadeMux I__6968 (
            .O(N__34745),
            .I(N__34742));
    InMux I__6967 (
            .O(N__34742),
            .I(N__34739));
    LocalMux I__6966 (
            .O(N__34739),
            .I(\phase_controller_inst2.stoper_tr.running_1_sqmuxa ));
    InMux I__6965 (
            .O(N__34736),
            .I(N__34731));
    InMux I__6964 (
            .O(N__34735),
            .I(N__34726));
    InMux I__6963 (
            .O(N__34734),
            .I(N__34726));
    LocalMux I__6962 (
            .O(N__34731),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    LocalMux I__6961 (
            .O(N__34726),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    InMux I__6960 (
            .O(N__34721),
            .I(N__34709));
    InMux I__6959 (
            .O(N__34720),
            .I(N__34709));
    InMux I__6958 (
            .O(N__34719),
            .I(N__34709));
    InMux I__6957 (
            .O(N__34718),
            .I(N__34702));
    InMux I__6956 (
            .O(N__34717),
            .I(N__34702));
    InMux I__6955 (
            .O(N__34716),
            .I(N__34702));
    LocalMux I__6954 (
            .O(N__34709),
            .I(N__34697));
    LocalMux I__6953 (
            .O(N__34702),
            .I(N__34697));
    Span4Mux_h I__6952 (
            .O(N__34697),
            .I(N__34693));
    InMux I__6951 (
            .O(N__34696),
            .I(N__34690));
    Span4Mux_v I__6950 (
            .O(N__34693),
            .I(N__34687));
    LocalMux I__6949 (
            .O(N__34690),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    Odrv4 I__6948 (
            .O(N__34687),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    InMux I__6947 (
            .O(N__34682),
            .I(N__34672));
    InMux I__6946 (
            .O(N__34681),
            .I(N__34672));
    InMux I__6945 (
            .O(N__34680),
            .I(N__34669));
    InMux I__6944 (
            .O(N__34679),
            .I(N__34664));
    InMux I__6943 (
            .O(N__34678),
            .I(N__34664));
    CascadeMux I__6942 (
            .O(N__34677),
            .I(N__34661));
    LocalMux I__6941 (
            .O(N__34672),
            .I(N__34657));
    LocalMux I__6940 (
            .O(N__34669),
            .I(N__34651));
    LocalMux I__6939 (
            .O(N__34664),
            .I(N__34651));
    InMux I__6938 (
            .O(N__34661),
            .I(N__34646));
    InMux I__6937 (
            .O(N__34660),
            .I(N__34646));
    Span4Mux_v I__6936 (
            .O(N__34657),
            .I(N__34643));
    InMux I__6935 (
            .O(N__34656),
            .I(N__34640));
    Span4Mux_v I__6934 (
            .O(N__34651),
            .I(N__34637));
    LocalMux I__6933 (
            .O(N__34646),
            .I(N__34632));
    Span4Mux_v I__6932 (
            .O(N__34643),
            .I(N__34632));
    LocalMux I__6931 (
            .O(N__34640),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv4 I__6930 (
            .O(N__34637),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv4 I__6929 (
            .O(N__34632),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    InMux I__6928 (
            .O(N__34625),
            .I(N__34622));
    LocalMux I__6927 (
            .O(N__34622),
            .I(N__34619));
    Span4Mux_v I__6926 (
            .O(N__34619),
            .I(N__34616));
    Span4Mux_h I__6925 (
            .O(N__34616),
            .I(N__34613));
    Span4Mux_h I__6924 (
            .O(N__34613),
            .I(N__34609));
    InMux I__6923 (
            .O(N__34612),
            .I(N__34606));
    Odrv4 I__6922 (
            .O(N__34609),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    LocalMux I__6921 (
            .O(N__34606),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    CascadeMux I__6920 (
            .O(N__34601),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ));
    InMux I__6919 (
            .O(N__34598),
            .I(N__34595));
    LocalMux I__6918 (
            .O(N__34595),
            .I(N__34592));
    Span4Mux_v I__6917 (
            .O(N__34592),
            .I(N__34589));
    Span4Mux_h I__6916 (
            .O(N__34589),
            .I(N__34586));
    Span4Mux_v I__6915 (
            .O(N__34586),
            .I(N__34581));
    InMux I__6914 (
            .O(N__34585),
            .I(N__34576));
    InMux I__6913 (
            .O(N__34584),
            .I(N__34576));
    Odrv4 I__6912 (
            .O(N__34581),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    LocalMux I__6911 (
            .O(N__34576),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    InMux I__6910 (
            .O(N__34571),
            .I(N__34568));
    LocalMux I__6909 (
            .O(N__34568),
            .I(N__34565));
    Odrv12 I__6908 (
            .O(N__34565),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ));
    CascadeMux I__6907 (
            .O(N__34562),
            .I(N__34558));
    InMux I__6906 (
            .O(N__34561),
            .I(N__34555));
    InMux I__6905 (
            .O(N__34558),
            .I(N__34552));
    LocalMux I__6904 (
            .O(N__34555),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    LocalMux I__6903 (
            .O(N__34552),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    CascadeMux I__6902 (
            .O(N__34547),
            .I(N__34544));
    InMux I__6901 (
            .O(N__34544),
            .I(N__34541));
    LocalMux I__6900 (
            .O(N__34541),
            .I(elapsed_time_ns_1_RNITCIF91_0_23));
    CascadeMux I__6899 (
            .O(N__34538),
            .I(elapsed_time_ns_1_RNITCIF91_0_23_cascade_));
    InMux I__6898 (
            .O(N__34535),
            .I(N__34531));
    InMux I__6897 (
            .O(N__34534),
            .I(N__34528));
    LocalMux I__6896 (
            .O(N__34531),
            .I(elapsed_time_ns_1_RNIUDIF91_0_24));
    LocalMux I__6895 (
            .O(N__34528),
            .I(elapsed_time_ns_1_RNIUDIF91_0_24));
    InMux I__6894 (
            .O(N__34523),
            .I(N__34520));
    LocalMux I__6893 (
            .O(N__34520),
            .I(N__34517));
    Odrv4 I__6892 (
            .O(N__34517),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ));
    CascadeMux I__6891 (
            .O(N__34514),
            .I(\phase_controller_inst1.N_55_cascade_ ));
    InMux I__6890 (
            .O(N__34511),
            .I(N__34502));
    InMux I__6889 (
            .O(N__34510),
            .I(N__34502));
    InMux I__6888 (
            .O(N__34509),
            .I(N__34502));
    LocalMux I__6887 (
            .O(N__34502),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    CascadeMux I__6886 (
            .O(N__34499),
            .I(N__34495));
    InMux I__6885 (
            .O(N__34498),
            .I(N__34490));
    InMux I__6884 (
            .O(N__34495),
            .I(N__34490));
    LocalMux I__6883 (
            .O(N__34490),
            .I(N__34487));
    Odrv4 I__6882 (
            .O(N__34487),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__6881 (
            .O(N__34484),
            .I(N__34478));
    InMux I__6880 (
            .O(N__34483),
            .I(N__34478));
    LocalMux I__6879 (
            .O(N__34478),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__6878 (
            .O(N__34475),
            .I(N__34468));
    InMux I__6877 (
            .O(N__34474),
            .I(N__34468));
    InMux I__6876 (
            .O(N__34473),
            .I(N__34465));
    LocalMux I__6875 (
            .O(N__34468),
            .I(N__34462));
    LocalMux I__6874 (
            .O(N__34465),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8 ));
    Odrv4 I__6873 (
            .O(N__34462),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8 ));
    InMux I__6872 (
            .O(N__34457),
            .I(N__34454));
    LocalMux I__6871 (
            .O(N__34454),
            .I(\delay_measurement_inst.delay_tr_timer.N_347 ));
    CascadeMux I__6870 (
            .O(N__34451),
            .I(\delay_measurement_inst.delay_tr_timer.N_347_cascade_ ));
    CascadeMux I__6869 (
            .O(N__34448),
            .I(N__34443));
    InMux I__6868 (
            .O(N__34447),
            .I(N__34440));
    InMux I__6867 (
            .O(N__34446),
            .I(N__34435));
    InMux I__6866 (
            .O(N__34443),
            .I(N__34435));
    LocalMux I__6865 (
            .O(N__34440),
            .I(N__34432));
    LocalMux I__6864 (
            .O(N__34435),
            .I(N__34429));
    Odrv4 I__6863 (
            .O(N__34432),
            .I(\delay_measurement_inst.delay_tr_timer.N_365 ));
    Odrv12 I__6862 (
            .O(N__34429),
            .I(\delay_measurement_inst.delay_tr_timer.N_365 ));
    InMux I__6861 (
            .O(N__34424),
            .I(N__34420));
    CascadeMux I__6860 (
            .O(N__34423),
            .I(N__34417));
    LocalMux I__6859 (
            .O(N__34420),
            .I(N__34414));
    InMux I__6858 (
            .O(N__34417),
            .I(N__34411));
    Odrv4 I__6857 (
            .O(N__34414),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    LocalMux I__6856 (
            .O(N__34411),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__6855 (
            .O(N__34406),
            .I(N__34401));
    InMux I__6854 (
            .O(N__34405),
            .I(N__34396));
    InMux I__6853 (
            .O(N__34404),
            .I(N__34396));
    LocalMux I__6852 (
            .O(N__34401),
            .I(N__34393));
    LocalMux I__6851 (
            .O(N__34396),
            .I(N__34390));
    Odrv4 I__6850 (
            .O(N__34393),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_7 ));
    Odrv12 I__6849 (
            .O(N__34390),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_7 ));
    InMux I__6848 (
            .O(N__34385),
            .I(N__34381));
    InMux I__6847 (
            .O(N__34384),
            .I(N__34378));
    LocalMux I__6846 (
            .O(N__34381),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    LocalMux I__6845 (
            .O(N__34378),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__6844 (
            .O(N__34373),
            .I(N__34370));
    LocalMux I__6843 (
            .O(N__34370),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_6 ));
    CascadeMux I__6842 (
            .O(N__34367),
            .I(N__34363));
    InMux I__6841 (
            .O(N__34366),
            .I(N__34360));
    InMux I__6840 (
            .O(N__34363),
            .I(N__34357));
    LocalMux I__6839 (
            .O(N__34360),
            .I(\delay_measurement_inst.delay_tr_timer.N_341 ));
    LocalMux I__6838 (
            .O(N__34357),
            .I(\delay_measurement_inst.delay_tr_timer.N_341 ));
    CascadeMux I__6837 (
            .O(N__34352),
            .I(N__34348));
    InMux I__6836 (
            .O(N__34351),
            .I(N__34345));
    InMux I__6835 (
            .O(N__34348),
            .I(N__34342));
    LocalMux I__6834 (
            .O(N__34345),
            .I(N__34339));
    LocalMux I__6833 (
            .O(N__34342),
            .I(N__34335));
    Span4Mux_v I__6832 (
            .O(N__34339),
            .I(N__34332));
    InMux I__6831 (
            .O(N__34338),
            .I(N__34329));
    Span4Mux_v I__6830 (
            .O(N__34335),
            .I(N__34326));
    Odrv4 I__6829 (
            .O(N__34332),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__6828 (
            .O(N__34329),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    Odrv4 I__6827 (
            .O(N__34326),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    InMux I__6826 (
            .O(N__34319),
            .I(N__34312));
    InMux I__6825 (
            .O(N__34318),
            .I(N__34312));
    InMux I__6824 (
            .O(N__34317),
            .I(N__34309));
    LocalMux I__6823 (
            .O(N__34312),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    LocalMux I__6822 (
            .O(N__34309),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    CEMux I__6821 (
            .O(N__34304),
            .I(N__34286));
    CEMux I__6820 (
            .O(N__34303),
            .I(N__34286));
    CEMux I__6819 (
            .O(N__34302),
            .I(N__34286));
    CEMux I__6818 (
            .O(N__34301),
            .I(N__34286));
    CEMux I__6817 (
            .O(N__34300),
            .I(N__34286));
    CEMux I__6816 (
            .O(N__34299),
            .I(N__34286));
    GlobalMux I__6815 (
            .O(N__34286),
            .I(N__34283));
    gio2CtrlBuf I__6814 (
            .O(N__34283),
            .I(\delay_measurement_inst.delay_tr_timer.N_434_i_g ));
    InMux I__6813 (
            .O(N__34280),
            .I(N__34277));
    LocalMux I__6812 (
            .O(N__34277),
            .I(N__34274));
    Odrv4 I__6811 (
            .O(N__34274),
            .I(\delay_measurement_inst.delay_tr_timer.N_348 ));
    InMux I__6810 (
            .O(N__34271),
            .I(N__34267));
    InMux I__6809 (
            .O(N__34270),
            .I(N__34264));
    LocalMux I__6808 (
            .O(N__34267),
            .I(\delay_measurement_inst.delay_tr_timer.N_367 ));
    LocalMux I__6807 (
            .O(N__34264),
            .I(\delay_measurement_inst.delay_tr_timer.N_367 ));
    CascadeMux I__6806 (
            .O(N__34259),
            .I(\delay_measurement_inst.delay_tr_timer.N_349_cascade_ ));
    CascadeMux I__6805 (
            .O(N__34256),
            .I(\delay_measurement_inst.delay_tr_timer.N_363_cascade_ ));
    CascadeMux I__6804 (
            .O(N__34253),
            .I(N__34249));
    InMux I__6803 (
            .O(N__34252),
            .I(N__34246));
    InMux I__6802 (
            .O(N__34249),
            .I(N__34243));
    LocalMux I__6801 (
            .O(N__34246),
            .I(\delay_measurement_inst.delay_tr_timer.N_380 ));
    LocalMux I__6800 (
            .O(N__34243),
            .I(\delay_measurement_inst.delay_tr_timer.N_380 ));
    CascadeMux I__6799 (
            .O(N__34238),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9_cascade_ ));
    CascadeMux I__6798 (
            .O(N__34235),
            .I(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0_cascade_ ));
    InMux I__6797 (
            .O(N__34232),
            .I(N__34225));
    InMux I__6796 (
            .O(N__34231),
            .I(N__34225));
    InMux I__6795 (
            .O(N__34230),
            .I(N__34222));
    LocalMux I__6794 (
            .O(N__34225),
            .I(\delay_measurement_inst.delay_tr_timer.N_378 ));
    LocalMux I__6793 (
            .O(N__34222),
            .I(\delay_measurement_inst.delay_tr_timer.N_378 ));
    InMux I__6792 (
            .O(N__34217),
            .I(N__34214));
    LocalMux I__6791 (
            .O(N__34214),
            .I(N__34211));
    Odrv4 I__6790 (
            .O(N__34211),
            .I(\delay_measurement_inst.delay_tr_timer.N_359_1 ));
    InMux I__6789 (
            .O(N__34208),
            .I(N__34202));
    InMux I__6788 (
            .O(N__34207),
            .I(N__34202));
    LocalMux I__6787 (
            .O(N__34202),
            .I(N__34198));
    InMux I__6786 (
            .O(N__34201),
            .I(N__34195));
    Span4Mux_v I__6785 (
            .O(N__34198),
            .I(N__34192));
    LocalMux I__6784 (
            .O(N__34195),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    Odrv4 I__6783 (
            .O(N__34192),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    CascadeMux I__6782 (
            .O(N__34187),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_ ));
    CascadeMux I__6781 (
            .O(N__34184),
            .I(\delay_measurement_inst.delay_tr_timer.N_359_1_cascade_ ));
    InMux I__6780 (
            .O(N__34181),
            .I(N__34178));
    LocalMux I__6779 (
            .O(N__34178),
            .I(\delay_measurement_inst.delay_tr_timer.N_345 ));
    CascadeMux I__6778 (
            .O(N__34175),
            .I(\delay_measurement_inst.delay_tr_timer.N_345_cascade_ ));
    CascadeMux I__6777 (
            .O(N__34172),
            .I(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_ ));
    InMux I__6776 (
            .O(N__34169),
            .I(N__34166));
    LocalMux I__6775 (
            .O(N__34166),
            .I(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5 ));
    InMux I__6774 (
            .O(N__34163),
            .I(N__34160));
    LocalMux I__6773 (
            .O(N__34160),
            .I(N__34156));
    InMux I__6772 (
            .O(N__34159),
            .I(N__34153));
    Span4Mux_s1_v I__6771 (
            .O(N__34156),
            .I(N__34148));
    LocalMux I__6770 (
            .O(N__34153),
            .I(N__34148));
    Span4Mux_v I__6769 (
            .O(N__34148),
            .I(N__34143));
    InMux I__6768 (
            .O(N__34147),
            .I(N__34140));
    InMux I__6767 (
            .O(N__34146),
            .I(N__34137));
    Span4Mux_h I__6766 (
            .O(N__34143),
            .I(N__34134));
    LocalMux I__6765 (
            .O(N__34140),
            .I(N__34131));
    LocalMux I__6764 (
            .O(N__34137),
            .I(N__34128));
    Sp12to4 I__6763 (
            .O(N__34134),
            .I(N__34125));
    Span4Mux_v I__6762 (
            .O(N__34131),
            .I(N__34122));
    Span4Mux_v I__6761 (
            .O(N__34128),
            .I(N__34119));
    Span12Mux_v I__6760 (
            .O(N__34125),
            .I(N__34116));
    Sp12to4 I__6759 (
            .O(N__34122),
            .I(N__34113));
    Span4Mux_h I__6758 (
            .O(N__34119),
            .I(N__34110));
    Span12Mux_v I__6757 (
            .O(N__34116),
            .I(N__34107));
    Span12Mux_h I__6756 (
            .O(N__34113),
            .I(N__34102));
    Sp12to4 I__6755 (
            .O(N__34110),
            .I(N__34102));
    Span12Mux_h I__6754 (
            .O(N__34107),
            .I(N__34099));
    Span12Mux_v I__6753 (
            .O(N__34102),
            .I(N__34096));
    Odrv12 I__6752 (
            .O(N__34099),
            .I(start_stop_c));
    Odrv12 I__6751 (
            .O(N__34096),
            .I(start_stop_c));
    InMux I__6750 (
            .O(N__34091),
            .I(N__34088));
    LocalMux I__6749 (
            .O(N__34088),
            .I(N__34085));
    Span4Mux_v I__6748 (
            .O(N__34085),
            .I(N__34082));
    Span4Mux_v I__6747 (
            .O(N__34082),
            .I(N__34079));
    Odrv4 I__6746 (
            .O(N__34079),
            .I(\current_shift_inst.elapsed_time_ns_s1_fast_31 ));
    IoInMux I__6745 (
            .O(N__34076),
            .I(N__34073));
    LocalMux I__6744 (
            .O(N__34073),
            .I(N__34070));
    Span4Mux_s2_v I__6743 (
            .O(N__34070),
            .I(N__34067));
    Odrv4 I__6742 (
            .O(N__34067),
            .I(s2_phy_c));
    InMux I__6741 (
            .O(N__34064),
            .I(N__34060));
    InMux I__6740 (
            .O(N__34063),
            .I(N__34056));
    LocalMux I__6739 (
            .O(N__34060),
            .I(N__34053));
    InMux I__6738 (
            .O(N__34059),
            .I(N__34050));
    LocalMux I__6737 (
            .O(N__34056),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    Odrv12 I__6736 (
            .O(N__34053),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__6735 (
            .O(N__34050),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    InMux I__6734 (
            .O(N__34043),
            .I(N__34040));
    LocalMux I__6733 (
            .O(N__34040),
            .I(N__34037));
    Span4Mux_h I__6732 (
            .O(N__34037),
            .I(N__34033));
    InMux I__6731 (
            .O(N__34036),
            .I(N__34030));
    Span4Mux_v I__6730 (
            .O(N__34033),
            .I(N__34021));
    LocalMux I__6729 (
            .O(N__34030),
            .I(N__34021));
    InMux I__6728 (
            .O(N__34029),
            .I(N__34018));
    InMux I__6727 (
            .O(N__34028),
            .I(N__34013));
    InMux I__6726 (
            .O(N__34027),
            .I(N__34013));
    InMux I__6725 (
            .O(N__34026),
            .I(N__34010));
    Odrv4 I__6724 (
            .O(N__34021),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    LocalMux I__6723 (
            .O(N__34018),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    LocalMux I__6722 (
            .O(N__34013),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    LocalMux I__6721 (
            .O(N__34010),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    CascadeMux I__6720 (
            .O(N__34001),
            .I(N__33997));
    InMux I__6719 (
            .O(N__34000),
            .I(N__33993));
    InMux I__6718 (
            .O(N__33997),
            .I(N__33988));
    InMux I__6717 (
            .O(N__33996),
            .I(N__33988));
    LocalMux I__6716 (
            .O(N__33993),
            .I(N__33985));
    LocalMux I__6715 (
            .O(N__33988),
            .I(N__33982));
    Sp12to4 I__6714 (
            .O(N__33985),
            .I(N__33979));
    Span4Mux_v I__6713 (
            .O(N__33982),
            .I(N__33976));
    Span12Mux_h I__6712 (
            .O(N__33979),
            .I(N__33973));
    Span4Mux_v I__6711 (
            .O(N__33976),
            .I(N__33970));
    Span12Mux_v I__6710 (
            .O(N__33973),
            .I(N__33967));
    Odrv4 I__6709 (
            .O(N__33970),
            .I(il_min_comp2_D2));
    Odrv12 I__6708 (
            .O(N__33967),
            .I(il_min_comp2_D2));
    InMux I__6707 (
            .O(N__33962),
            .I(N__33959));
    LocalMux I__6706 (
            .O(N__33959),
            .I(\phase_controller_inst2.start_timer_tr_0_sqmuxa ));
    CascadeMux I__6705 (
            .O(N__33956),
            .I(N__33953));
    InMux I__6704 (
            .O(N__33953),
            .I(N__33950));
    LocalMux I__6703 (
            .O(N__33950),
            .I(N__33947));
    Sp12to4 I__6702 (
            .O(N__33947),
            .I(N__33944));
    Odrv12 I__6701 (
            .O(N__33944),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ));
    CascadeMux I__6700 (
            .O(N__33941),
            .I(N__33936));
    InMux I__6699 (
            .O(N__33940),
            .I(N__33933));
    InMux I__6698 (
            .O(N__33939),
            .I(N__33930));
    InMux I__6697 (
            .O(N__33936),
            .I(N__33926));
    LocalMux I__6696 (
            .O(N__33933),
            .I(N__33923));
    LocalMux I__6695 (
            .O(N__33930),
            .I(N__33920));
    InMux I__6694 (
            .O(N__33929),
            .I(N__33917));
    LocalMux I__6693 (
            .O(N__33926),
            .I(N__33914));
    Span4Mux_v I__6692 (
            .O(N__33923),
            .I(N__33905));
    Span4Mux_v I__6691 (
            .O(N__33920),
            .I(N__33905));
    LocalMux I__6690 (
            .O(N__33917),
            .I(N__33905));
    Span4Mux_v I__6689 (
            .O(N__33914),
            .I(N__33905));
    Odrv4 I__6688 (
            .O(N__33905),
            .I(elapsed_time_ns_1_RNI3VBED1_0_16));
    InMux I__6687 (
            .O(N__33902),
            .I(N__33899));
    LocalMux I__6686 (
            .O(N__33899),
            .I(N__33895));
    CascadeMux I__6685 (
            .O(N__33898),
            .I(N__33892));
    Span4Mux_h I__6684 (
            .O(N__33895),
            .I(N__33888));
    InMux I__6683 (
            .O(N__33892),
            .I(N__33883));
    InMux I__6682 (
            .O(N__33891),
            .I(N__33883));
    Odrv4 I__6681 (
            .O(N__33888),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    LocalMux I__6680 (
            .O(N__33883),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    InMux I__6679 (
            .O(N__33878),
            .I(N__33875));
    LocalMux I__6678 (
            .O(N__33875),
            .I(N__33872));
    Span4Mux_h I__6677 (
            .O(N__33872),
            .I(N__33869));
    Odrv4 I__6676 (
            .O(N__33869),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16 ));
    CascadeMux I__6675 (
            .O(N__33866),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ));
    InMux I__6674 (
            .O(N__33863),
            .I(N__33860));
    LocalMux I__6673 (
            .O(N__33860),
            .I(N__33857));
    Span4Mux_v I__6672 (
            .O(N__33857),
            .I(N__33854));
    Odrv4 I__6671 (
            .O(N__33854),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ));
    InMux I__6670 (
            .O(N__33851),
            .I(N__33848));
    LocalMux I__6669 (
            .O(N__33848),
            .I(N__33844));
    InMux I__6668 (
            .O(N__33847),
            .I(N__33841));
    Span4Mux_h I__6667 (
            .O(N__33844),
            .I(N__33837));
    LocalMux I__6666 (
            .O(N__33841),
            .I(N__33834));
    InMux I__6665 (
            .O(N__33840),
            .I(N__33831));
    Span4Mux_v I__6664 (
            .O(N__33837),
            .I(N__33828));
    Odrv4 I__6663 (
            .O(N__33834),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    LocalMux I__6662 (
            .O(N__33831),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    Odrv4 I__6661 (
            .O(N__33828),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    InMux I__6660 (
            .O(N__33821),
            .I(N__33816));
    InMux I__6659 (
            .O(N__33820),
            .I(N__33810));
    InMux I__6658 (
            .O(N__33819),
            .I(N__33810));
    LocalMux I__6657 (
            .O(N__33816),
            .I(N__33807));
    InMux I__6656 (
            .O(N__33815),
            .I(N__33804));
    LocalMux I__6655 (
            .O(N__33810),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    Odrv4 I__6654 (
            .O(N__33807),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    LocalMux I__6653 (
            .O(N__33804),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    ClkMux I__6652 (
            .O(N__33797),
            .I(N__33794));
    GlobalMux I__6651 (
            .O(N__33794),
            .I(N__33791));
    gio2CtrlBuf I__6650 (
            .O(N__33791),
            .I(delay_tr_input_c_g));
    InMux I__6649 (
            .O(N__33788),
            .I(N__33785));
    LocalMux I__6648 (
            .O(N__33785),
            .I(N__33782));
    Span4Mux_v I__6647 (
            .O(N__33782),
            .I(N__33779));
    Odrv4 I__6646 (
            .O(N__33779),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ));
    CascadeMux I__6645 (
            .O(N__33776),
            .I(N__33770));
    CascadeMux I__6644 (
            .O(N__33775),
            .I(N__33767));
    InMux I__6643 (
            .O(N__33774),
            .I(N__33752));
    InMux I__6642 (
            .O(N__33773),
            .I(N__33749));
    InMux I__6641 (
            .O(N__33770),
            .I(N__33746));
    InMux I__6640 (
            .O(N__33767),
            .I(N__33738));
    InMux I__6639 (
            .O(N__33766),
            .I(N__33735));
    InMux I__6638 (
            .O(N__33765),
            .I(N__33728));
    InMux I__6637 (
            .O(N__33764),
            .I(N__33728));
    InMux I__6636 (
            .O(N__33763),
            .I(N__33728));
    CascadeMux I__6635 (
            .O(N__33762),
            .I(N__33722));
    CascadeMux I__6634 (
            .O(N__33761),
            .I(N__33719));
    CascadeMux I__6633 (
            .O(N__33760),
            .I(N__33713));
    CascadeMux I__6632 (
            .O(N__33759),
            .I(N__33709));
    CascadeMux I__6631 (
            .O(N__33758),
            .I(N__33704));
    CascadeMux I__6630 (
            .O(N__33757),
            .I(N__33699));
    CascadeMux I__6629 (
            .O(N__33756),
            .I(N__33696));
    InMux I__6628 (
            .O(N__33755),
            .I(N__33688));
    LocalMux I__6627 (
            .O(N__33752),
            .I(N__33685));
    LocalMux I__6626 (
            .O(N__33749),
            .I(N__33680));
    LocalMux I__6625 (
            .O(N__33746),
            .I(N__33680));
    CascadeMux I__6624 (
            .O(N__33745),
            .I(N__33673));
    InMux I__6623 (
            .O(N__33744),
            .I(N__33666));
    InMux I__6622 (
            .O(N__33743),
            .I(N__33661));
    InMux I__6621 (
            .O(N__33742),
            .I(N__33661));
    InMux I__6620 (
            .O(N__33741),
            .I(N__33658));
    LocalMux I__6619 (
            .O(N__33738),
            .I(N__33651));
    LocalMux I__6618 (
            .O(N__33735),
            .I(N__33651));
    LocalMux I__6617 (
            .O(N__33728),
            .I(N__33651));
    InMux I__6616 (
            .O(N__33727),
            .I(N__33644));
    InMux I__6615 (
            .O(N__33726),
            .I(N__33644));
    InMux I__6614 (
            .O(N__33725),
            .I(N__33644));
    InMux I__6613 (
            .O(N__33722),
            .I(N__33631));
    InMux I__6612 (
            .O(N__33719),
            .I(N__33631));
    InMux I__6611 (
            .O(N__33718),
            .I(N__33631));
    InMux I__6610 (
            .O(N__33717),
            .I(N__33631));
    InMux I__6609 (
            .O(N__33716),
            .I(N__33631));
    InMux I__6608 (
            .O(N__33713),
            .I(N__33631));
    InMux I__6607 (
            .O(N__33712),
            .I(N__33616));
    InMux I__6606 (
            .O(N__33709),
            .I(N__33616));
    InMux I__6605 (
            .O(N__33708),
            .I(N__33616));
    InMux I__6604 (
            .O(N__33707),
            .I(N__33616));
    InMux I__6603 (
            .O(N__33704),
            .I(N__33616));
    InMux I__6602 (
            .O(N__33703),
            .I(N__33616));
    InMux I__6601 (
            .O(N__33702),
            .I(N__33616));
    InMux I__6600 (
            .O(N__33699),
            .I(N__33603));
    InMux I__6599 (
            .O(N__33696),
            .I(N__33603));
    InMux I__6598 (
            .O(N__33695),
            .I(N__33603));
    InMux I__6597 (
            .O(N__33694),
            .I(N__33603));
    InMux I__6596 (
            .O(N__33693),
            .I(N__33603));
    InMux I__6595 (
            .O(N__33692),
            .I(N__33603));
    InMux I__6594 (
            .O(N__33691),
            .I(N__33594));
    LocalMux I__6593 (
            .O(N__33688),
            .I(N__33587));
    Span4Mux_v I__6592 (
            .O(N__33685),
            .I(N__33587));
    Span4Mux_v I__6591 (
            .O(N__33680),
            .I(N__33587));
    InMux I__6590 (
            .O(N__33679),
            .I(N__33584));
    InMux I__6589 (
            .O(N__33678),
            .I(N__33579));
    InMux I__6588 (
            .O(N__33677),
            .I(N__33579));
    InMux I__6587 (
            .O(N__33676),
            .I(N__33566));
    InMux I__6586 (
            .O(N__33673),
            .I(N__33566));
    InMux I__6585 (
            .O(N__33672),
            .I(N__33566));
    InMux I__6584 (
            .O(N__33671),
            .I(N__33566));
    InMux I__6583 (
            .O(N__33670),
            .I(N__33566));
    InMux I__6582 (
            .O(N__33669),
            .I(N__33566));
    LocalMux I__6581 (
            .O(N__33666),
            .I(N__33561));
    LocalMux I__6580 (
            .O(N__33661),
            .I(N__33561));
    LocalMux I__6579 (
            .O(N__33658),
            .I(N__33548));
    Span4Mux_h I__6578 (
            .O(N__33651),
            .I(N__33548));
    LocalMux I__6577 (
            .O(N__33644),
            .I(N__33548));
    LocalMux I__6576 (
            .O(N__33631),
            .I(N__33548));
    LocalMux I__6575 (
            .O(N__33616),
            .I(N__33548));
    LocalMux I__6574 (
            .O(N__33603),
            .I(N__33548));
    InMux I__6573 (
            .O(N__33602),
            .I(N__33545));
    InMux I__6572 (
            .O(N__33601),
            .I(N__33534));
    InMux I__6571 (
            .O(N__33600),
            .I(N__33534));
    InMux I__6570 (
            .O(N__33599),
            .I(N__33534));
    InMux I__6569 (
            .O(N__33598),
            .I(N__33534));
    InMux I__6568 (
            .O(N__33597),
            .I(N__33534));
    LocalMux I__6567 (
            .O(N__33594),
            .I(N__33529));
    Span4Mux_h I__6566 (
            .O(N__33587),
            .I(N__33529));
    LocalMux I__6565 (
            .O(N__33584),
            .I(N__33526));
    LocalMux I__6564 (
            .O(N__33579),
            .I(N__33523));
    LocalMux I__6563 (
            .O(N__33566),
            .I(N__33516));
    Span4Mux_v I__6562 (
            .O(N__33561),
            .I(N__33516));
    Span4Mux_v I__6561 (
            .O(N__33548),
            .I(N__33516));
    LocalMux I__6560 (
            .O(N__33545),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    LocalMux I__6559 (
            .O(N__33534),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv4 I__6558 (
            .O(N__33529),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv4 I__6557 (
            .O(N__33526),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv12 I__6556 (
            .O(N__33523),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv4 I__6555 (
            .O(N__33516),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    CascadeMux I__6554 (
            .O(N__33503),
            .I(N__33498));
    InMux I__6553 (
            .O(N__33502),
            .I(N__33495));
    InMux I__6552 (
            .O(N__33501),
            .I(N__33490));
    InMux I__6551 (
            .O(N__33498),
            .I(N__33490));
    LocalMux I__6550 (
            .O(N__33495),
            .I(N__33485));
    LocalMux I__6549 (
            .O(N__33490),
            .I(N__33485));
    Span4Mux_h I__6548 (
            .O(N__33485),
            .I(N__33482));
    Span4Mux_h I__6547 (
            .O(N__33482),
            .I(N__33479));
    Odrv4 I__6546 (
            .O(N__33479),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_i_0_12 ));
    InMux I__6545 (
            .O(N__33476),
            .I(N__33473));
    LocalMux I__6544 (
            .O(N__33473),
            .I(N__33470));
    Span4Mux_h I__6543 (
            .O(N__33470),
            .I(N__33467));
    Odrv4 I__6542 (
            .O(N__33467),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ));
    InMux I__6541 (
            .O(N__33464),
            .I(N__33457));
    InMux I__6540 (
            .O(N__33463),
            .I(N__33457));
    InMux I__6539 (
            .O(N__33462),
            .I(N__33454));
    LocalMux I__6538 (
            .O(N__33457),
            .I(N__33451));
    LocalMux I__6537 (
            .O(N__33454),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    Odrv12 I__6536 (
            .O(N__33451),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    CascadeMux I__6535 (
            .O(N__33446),
            .I(N__33443));
    InMux I__6534 (
            .O(N__33443),
            .I(N__33439));
    InMux I__6533 (
            .O(N__33442),
            .I(N__33436));
    LocalMux I__6532 (
            .O(N__33439),
            .I(N__33433));
    LocalMux I__6531 (
            .O(N__33436),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    Odrv12 I__6530 (
            .O(N__33433),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    InMux I__6529 (
            .O(N__33428),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__6528 (
            .O(N__33425),
            .I(N__33421));
    InMux I__6527 (
            .O(N__33424),
            .I(N__33418));
    LocalMux I__6526 (
            .O(N__33421),
            .I(N__33415));
    LocalMux I__6525 (
            .O(N__33418),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    Odrv12 I__6524 (
            .O(N__33415),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CascadeMux I__6523 (
            .O(N__33410),
            .I(N__33407));
    InMux I__6522 (
            .O(N__33407),
            .I(N__33403));
    InMux I__6521 (
            .O(N__33406),
            .I(N__33400));
    LocalMux I__6520 (
            .O(N__33403),
            .I(N__33394));
    LocalMux I__6519 (
            .O(N__33400),
            .I(N__33394));
    InMux I__6518 (
            .O(N__33399),
            .I(N__33391));
    Span4Mux_v I__6517 (
            .O(N__33394),
            .I(N__33388));
    LocalMux I__6516 (
            .O(N__33391),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    Odrv4 I__6515 (
            .O(N__33388),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__6514 (
            .O(N__33383),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__6513 (
            .O(N__33380),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__6512 (
            .O(N__33377),
            .I(N__33373));
    InMux I__6511 (
            .O(N__33376),
            .I(N__33370));
    LocalMux I__6510 (
            .O(N__33373),
            .I(N__33367));
    LocalMux I__6509 (
            .O(N__33370),
            .I(N__33361));
    Span4Mux_h I__6508 (
            .O(N__33367),
            .I(N__33361));
    InMux I__6507 (
            .O(N__33366),
            .I(N__33357));
    Span4Mux_v I__6506 (
            .O(N__33361),
            .I(N__33354));
    InMux I__6505 (
            .O(N__33360),
            .I(N__33351));
    LocalMux I__6504 (
            .O(N__33357),
            .I(N__33348));
    Span4Mux_v I__6503 (
            .O(N__33354),
            .I(N__33345));
    LocalMux I__6502 (
            .O(N__33351),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv4 I__6501 (
            .O(N__33348),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv4 I__6500 (
            .O(N__33345),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    CEMux I__6499 (
            .O(N__33338),
            .I(N__33332));
    CEMux I__6498 (
            .O(N__33337),
            .I(N__33329));
    CEMux I__6497 (
            .O(N__33336),
            .I(N__33326));
    CEMux I__6496 (
            .O(N__33335),
            .I(N__33323));
    LocalMux I__6495 (
            .O(N__33332),
            .I(N__33320));
    LocalMux I__6494 (
            .O(N__33329),
            .I(N__33317));
    LocalMux I__6493 (
            .O(N__33326),
            .I(N__33314));
    LocalMux I__6492 (
            .O(N__33323),
            .I(N__33311));
    Span4Mux_v I__6491 (
            .O(N__33320),
            .I(N__33308));
    Span4Mux_v I__6490 (
            .O(N__33317),
            .I(N__33305));
    Span4Mux_v I__6489 (
            .O(N__33314),
            .I(N__33302));
    Odrv12 I__6488 (
            .O(N__33311),
            .I(\delay_measurement_inst.delay_tr_timer.N_435_i ));
    Odrv4 I__6487 (
            .O(N__33308),
            .I(\delay_measurement_inst.delay_tr_timer.N_435_i ));
    Odrv4 I__6486 (
            .O(N__33305),
            .I(\delay_measurement_inst.delay_tr_timer.N_435_i ));
    Odrv4 I__6485 (
            .O(N__33302),
            .I(\delay_measurement_inst.delay_tr_timer.N_435_i ));
    InMux I__6484 (
            .O(N__33293),
            .I(N__33290));
    LocalMux I__6483 (
            .O(N__33290),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ));
    CascadeMux I__6482 (
            .O(N__33287),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0_cascade_ ));
    CascadeMux I__6481 (
            .O(N__33284),
            .I(\phase_controller_inst2.stoper_tr.running_1_sqmuxa_cascade_ ));
    InMux I__6480 (
            .O(N__33281),
            .I(N__33274));
    InMux I__6479 (
            .O(N__33280),
            .I(N__33274));
    InMux I__6478 (
            .O(N__33279),
            .I(N__33271));
    LocalMux I__6477 (
            .O(N__33274),
            .I(N__33268));
    LocalMux I__6476 (
            .O(N__33271),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    Odrv12 I__6475 (
            .O(N__33268),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__6474 (
            .O(N__33263),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__6473 (
            .O(N__33260),
            .I(N__33253));
    InMux I__6472 (
            .O(N__33259),
            .I(N__33253));
    InMux I__6471 (
            .O(N__33258),
            .I(N__33250));
    LocalMux I__6470 (
            .O(N__33253),
            .I(N__33247));
    LocalMux I__6469 (
            .O(N__33250),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    Odrv12 I__6468 (
            .O(N__33247),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__6467 (
            .O(N__33242),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__6466 (
            .O(N__33239),
            .I(N__33235));
    CascadeMux I__6465 (
            .O(N__33238),
            .I(N__33232));
    InMux I__6464 (
            .O(N__33235),
            .I(N__33226));
    InMux I__6463 (
            .O(N__33232),
            .I(N__33226));
    InMux I__6462 (
            .O(N__33231),
            .I(N__33223));
    LocalMux I__6461 (
            .O(N__33226),
            .I(N__33220));
    LocalMux I__6460 (
            .O(N__33223),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    Odrv12 I__6459 (
            .O(N__33220),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__6458 (
            .O(N__33215),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__6457 (
            .O(N__33212),
            .I(N__33208));
    CascadeMux I__6456 (
            .O(N__33211),
            .I(N__33205));
    InMux I__6455 (
            .O(N__33208),
            .I(N__33199));
    InMux I__6454 (
            .O(N__33205),
            .I(N__33199));
    InMux I__6453 (
            .O(N__33204),
            .I(N__33196));
    LocalMux I__6452 (
            .O(N__33199),
            .I(N__33193));
    LocalMux I__6451 (
            .O(N__33196),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    Odrv12 I__6450 (
            .O(N__33193),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__6449 (
            .O(N__33188),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__6448 (
            .O(N__33185),
            .I(N__33179));
    InMux I__6447 (
            .O(N__33184),
            .I(N__33179));
    LocalMux I__6446 (
            .O(N__33179),
            .I(N__33175));
    InMux I__6445 (
            .O(N__33178),
            .I(N__33172));
    Span4Mux_v I__6444 (
            .O(N__33175),
            .I(N__33169));
    LocalMux I__6443 (
            .O(N__33172),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    Odrv4 I__6442 (
            .O(N__33169),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__6441 (
            .O(N__33164),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__6440 (
            .O(N__33161),
            .I(N__33158));
    InMux I__6439 (
            .O(N__33158),
            .I(N__33154));
    InMux I__6438 (
            .O(N__33157),
            .I(N__33151));
    LocalMux I__6437 (
            .O(N__33154),
            .I(N__33145));
    LocalMux I__6436 (
            .O(N__33151),
            .I(N__33145));
    InMux I__6435 (
            .O(N__33150),
            .I(N__33142));
    Span4Mux_v I__6434 (
            .O(N__33145),
            .I(N__33139));
    LocalMux I__6433 (
            .O(N__33142),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    Odrv4 I__6432 (
            .O(N__33139),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__6431 (
            .O(N__33134),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__6430 (
            .O(N__33131),
            .I(N__33127));
    CascadeMux I__6429 (
            .O(N__33130),
            .I(N__33124));
    InMux I__6428 (
            .O(N__33127),
            .I(N__33121));
    InMux I__6427 (
            .O(N__33124),
            .I(N__33118));
    LocalMux I__6426 (
            .O(N__33121),
            .I(N__33112));
    LocalMux I__6425 (
            .O(N__33118),
            .I(N__33112));
    InMux I__6424 (
            .O(N__33117),
            .I(N__33109));
    Span4Mux_v I__6423 (
            .O(N__33112),
            .I(N__33106));
    LocalMux I__6422 (
            .O(N__33109),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    Odrv4 I__6421 (
            .O(N__33106),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__6420 (
            .O(N__33101),
            .I(bfn_13_12_0_));
    CascadeMux I__6419 (
            .O(N__33098),
            .I(N__33095));
    InMux I__6418 (
            .O(N__33095),
            .I(N__33090));
    InMux I__6417 (
            .O(N__33094),
            .I(N__33087));
    InMux I__6416 (
            .O(N__33093),
            .I(N__33084));
    LocalMux I__6415 (
            .O(N__33090),
            .I(N__33079));
    LocalMux I__6414 (
            .O(N__33087),
            .I(N__33079));
    LocalMux I__6413 (
            .O(N__33084),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    Odrv12 I__6412 (
            .O(N__33079),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    InMux I__6411 (
            .O(N__33074),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__6410 (
            .O(N__33071),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__6409 (
            .O(N__33068),
            .I(N__33062));
    InMux I__6408 (
            .O(N__33067),
            .I(N__33062));
    LocalMux I__6407 (
            .O(N__33062),
            .I(N__33058));
    InMux I__6406 (
            .O(N__33061),
            .I(N__33055));
    Span4Mux_v I__6405 (
            .O(N__33058),
            .I(N__33052));
    LocalMux I__6404 (
            .O(N__33055),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    Odrv4 I__6403 (
            .O(N__33052),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__6402 (
            .O(N__33047),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__6401 (
            .O(N__33044),
            .I(N__33038));
    InMux I__6400 (
            .O(N__33043),
            .I(N__33038));
    LocalMux I__6399 (
            .O(N__33038),
            .I(N__33034));
    InMux I__6398 (
            .O(N__33037),
            .I(N__33031));
    Span4Mux_v I__6397 (
            .O(N__33034),
            .I(N__33028));
    LocalMux I__6396 (
            .O(N__33031),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    Odrv4 I__6395 (
            .O(N__33028),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__6394 (
            .O(N__33023),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__6393 (
            .O(N__33020),
            .I(N__33016));
    CascadeMux I__6392 (
            .O(N__33019),
            .I(N__33013));
    InMux I__6391 (
            .O(N__33016),
            .I(N__33007));
    InMux I__6390 (
            .O(N__33013),
            .I(N__33007));
    InMux I__6389 (
            .O(N__33012),
            .I(N__33004));
    LocalMux I__6388 (
            .O(N__33007),
            .I(N__33001));
    LocalMux I__6387 (
            .O(N__33004),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    Odrv12 I__6386 (
            .O(N__33001),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__6385 (
            .O(N__32996),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__6384 (
            .O(N__32993),
            .I(N__32989));
    CascadeMux I__6383 (
            .O(N__32992),
            .I(N__32986));
    InMux I__6382 (
            .O(N__32989),
            .I(N__32980));
    InMux I__6381 (
            .O(N__32986),
            .I(N__32980));
    InMux I__6380 (
            .O(N__32985),
            .I(N__32977));
    LocalMux I__6379 (
            .O(N__32980),
            .I(N__32974));
    LocalMux I__6378 (
            .O(N__32977),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    Odrv12 I__6377 (
            .O(N__32974),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__6376 (
            .O(N__32969),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__6375 (
            .O(N__32966),
            .I(N__32960));
    InMux I__6374 (
            .O(N__32965),
            .I(N__32960));
    LocalMux I__6373 (
            .O(N__32960),
            .I(N__32956));
    InMux I__6372 (
            .O(N__32959),
            .I(N__32953));
    Span4Mux_v I__6371 (
            .O(N__32956),
            .I(N__32950));
    LocalMux I__6370 (
            .O(N__32953),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    Odrv4 I__6369 (
            .O(N__32950),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__6368 (
            .O(N__32945),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__6367 (
            .O(N__32942),
            .I(N__32939));
    InMux I__6366 (
            .O(N__32939),
            .I(N__32935));
    InMux I__6365 (
            .O(N__32938),
            .I(N__32932));
    LocalMux I__6364 (
            .O(N__32935),
            .I(N__32926));
    LocalMux I__6363 (
            .O(N__32932),
            .I(N__32926));
    InMux I__6362 (
            .O(N__32931),
            .I(N__32923));
    Span4Mux_v I__6361 (
            .O(N__32926),
            .I(N__32920));
    LocalMux I__6360 (
            .O(N__32923),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    Odrv4 I__6359 (
            .O(N__32920),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__6358 (
            .O(N__32915),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__6357 (
            .O(N__32912),
            .I(N__32909));
    InMux I__6356 (
            .O(N__32909),
            .I(N__32905));
    CascadeMux I__6355 (
            .O(N__32908),
            .I(N__32902));
    LocalMux I__6354 (
            .O(N__32905),
            .I(N__32898));
    InMux I__6353 (
            .O(N__32902),
            .I(N__32895));
    InMux I__6352 (
            .O(N__32901),
            .I(N__32892));
    Sp12to4 I__6351 (
            .O(N__32898),
            .I(N__32887));
    LocalMux I__6350 (
            .O(N__32895),
            .I(N__32887));
    LocalMux I__6349 (
            .O(N__32892),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    Odrv12 I__6348 (
            .O(N__32887),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__6347 (
            .O(N__32882),
            .I(bfn_13_11_0_));
    CascadeMux I__6346 (
            .O(N__32879),
            .I(N__32876));
    InMux I__6345 (
            .O(N__32876),
            .I(N__32873));
    LocalMux I__6344 (
            .O(N__32873),
            .I(N__32868));
    InMux I__6343 (
            .O(N__32872),
            .I(N__32865));
    InMux I__6342 (
            .O(N__32871),
            .I(N__32862));
    Sp12to4 I__6341 (
            .O(N__32868),
            .I(N__32857));
    LocalMux I__6340 (
            .O(N__32865),
            .I(N__32857));
    LocalMux I__6339 (
            .O(N__32862),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    Odrv12 I__6338 (
            .O(N__32857),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__6337 (
            .O(N__32852),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__6336 (
            .O(N__32849),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__6335 (
            .O(N__32846),
            .I(N__32842));
    InMux I__6334 (
            .O(N__32845),
            .I(N__32839));
    InMux I__6333 (
            .O(N__32842),
            .I(N__32836));
    LocalMux I__6332 (
            .O(N__32839),
            .I(N__32830));
    LocalMux I__6331 (
            .O(N__32836),
            .I(N__32830));
    InMux I__6330 (
            .O(N__32835),
            .I(N__32827));
    Span4Mux_v I__6329 (
            .O(N__32830),
            .I(N__32824));
    LocalMux I__6328 (
            .O(N__32827),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    Odrv4 I__6327 (
            .O(N__32824),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__6326 (
            .O(N__32819),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__6325 (
            .O(N__32816),
            .I(N__32810));
    InMux I__6324 (
            .O(N__32815),
            .I(N__32810));
    LocalMux I__6323 (
            .O(N__32810),
            .I(N__32806));
    InMux I__6322 (
            .O(N__32809),
            .I(N__32803));
    Span4Mux_v I__6321 (
            .O(N__32806),
            .I(N__32800));
    LocalMux I__6320 (
            .O(N__32803),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    Odrv4 I__6319 (
            .O(N__32800),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__6318 (
            .O(N__32795),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__6317 (
            .O(N__32792),
            .I(N__32788));
    CascadeMux I__6316 (
            .O(N__32791),
            .I(N__32785));
    InMux I__6315 (
            .O(N__32788),
            .I(N__32779));
    InMux I__6314 (
            .O(N__32785),
            .I(N__32779));
    InMux I__6313 (
            .O(N__32784),
            .I(N__32776));
    LocalMux I__6312 (
            .O(N__32779),
            .I(N__32773));
    LocalMux I__6311 (
            .O(N__32776),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    Odrv12 I__6310 (
            .O(N__32773),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__6309 (
            .O(N__32768),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__6308 (
            .O(N__32765),
            .I(N__32761));
    InMux I__6307 (
            .O(N__32764),
            .I(N__32757));
    InMux I__6306 (
            .O(N__32761),
            .I(N__32754));
    InMux I__6305 (
            .O(N__32760),
            .I(N__32751));
    LocalMux I__6304 (
            .O(N__32757),
            .I(N__32746));
    LocalMux I__6303 (
            .O(N__32754),
            .I(N__32746));
    LocalMux I__6302 (
            .O(N__32751),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    Odrv12 I__6301 (
            .O(N__32746),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__6300 (
            .O(N__32741),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__6299 (
            .O(N__32738),
            .I(N__32732));
    InMux I__6298 (
            .O(N__32737),
            .I(N__32732));
    LocalMux I__6297 (
            .O(N__32732),
            .I(N__32728));
    InMux I__6296 (
            .O(N__32731),
            .I(N__32725));
    Span4Mux_v I__6295 (
            .O(N__32728),
            .I(N__32722));
    LocalMux I__6294 (
            .O(N__32725),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    Odrv4 I__6293 (
            .O(N__32722),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__6292 (
            .O(N__32717),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__6291 (
            .O(N__32714),
            .I(N__32710));
    CascadeMux I__6290 (
            .O(N__32713),
            .I(N__32707));
    InMux I__6289 (
            .O(N__32710),
            .I(N__32702));
    InMux I__6288 (
            .O(N__32707),
            .I(N__32702));
    LocalMux I__6287 (
            .O(N__32702),
            .I(N__32698));
    InMux I__6286 (
            .O(N__32701),
            .I(N__32695));
    Span4Mux_v I__6285 (
            .O(N__32698),
            .I(N__32692));
    LocalMux I__6284 (
            .O(N__32695),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    Odrv4 I__6283 (
            .O(N__32692),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__6282 (
            .O(N__32687),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__6281 (
            .O(N__32684),
            .I(N__32681));
    InMux I__6280 (
            .O(N__32681),
            .I(N__32677));
    CascadeMux I__6279 (
            .O(N__32680),
            .I(N__32674));
    LocalMux I__6278 (
            .O(N__32677),
            .I(N__32670));
    InMux I__6277 (
            .O(N__32674),
            .I(N__32667));
    InMux I__6276 (
            .O(N__32673),
            .I(N__32664));
    Sp12to4 I__6275 (
            .O(N__32670),
            .I(N__32659));
    LocalMux I__6274 (
            .O(N__32667),
            .I(N__32659));
    LocalMux I__6273 (
            .O(N__32664),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    Odrv12 I__6272 (
            .O(N__32659),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__6271 (
            .O(N__32654),
            .I(bfn_13_10_0_));
    CascadeMux I__6270 (
            .O(N__32651),
            .I(N__32648));
    InMux I__6269 (
            .O(N__32648),
            .I(N__32645));
    LocalMux I__6268 (
            .O(N__32645),
            .I(N__32640));
    InMux I__6267 (
            .O(N__32644),
            .I(N__32637));
    InMux I__6266 (
            .O(N__32643),
            .I(N__32634));
    Sp12to4 I__6265 (
            .O(N__32640),
            .I(N__32629));
    LocalMux I__6264 (
            .O(N__32637),
            .I(N__32629));
    LocalMux I__6263 (
            .O(N__32634),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    Odrv12 I__6262 (
            .O(N__32629),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__6261 (
            .O(N__32624),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    InMux I__6260 (
            .O(N__32621),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    InMux I__6259 (
            .O(N__32618),
            .I(bfn_13_8_0_));
    InMux I__6258 (
            .O(N__32615),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    InMux I__6257 (
            .O(N__32612),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    InMux I__6256 (
            .O(N__32609),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__6255 (
            .O(N__32606),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__6254 (
            .O(N__32603),
            .I(N__32579));
    InMux I__6253 (
            .O(N__32602),
            .I(N__32579));
    InMux I__6252 (
            .O(N__32601),
            .I(N__32579));
    InMux I__6251 (
            .O(N__32600),
            .I(N__32579));
    InMux I__6250 (
            .O(N__32599),
            .I(N__32570));
    InMux I__6249 (
            .O(N__32598),
            .I(N__32570));
    InMux I__6248 (
            .O(N__32597),
            .I(N__32570));
    InMux I__6247 (
            .O(N__32596),
            .I(N__32570));
    InMux I__6246 (
            .O(N__32595),
            .I(N__32547));
    InMux I__6245 (
            .O(N__32594),
            .I(N__32547));
    InMux I__6244 (
            .O(N__32593),
            .I(N__32547));
    InMux I__6243 (
            .O(N__32592),
            .I(N__32547));
    InMux I__6242 (
            .O(N__32591),
            .I(N__32538));
    InMux I__6241 (
            .O(N__32590),
            .I(N__32538));
    InMux I__6240 (
            .O(N__32589),
            .I(N__32538));
    InMux I__6239 (
            .O(N__32588),
            .I(N__32538));
    LocalMux I__6238 (
            .O(N__32579),
            .I(N__32535));
    LocalMux I__6237 (
            .O(N__32570),
            .I(N__32532));
    InMux I__6236 (
            .O(N__32569),
            .I(N__32527));
    InMux I__6235 (
            .O(N__32568),
            .I(N__32527));
    InMux I__6234 (
            .O(N__32567),
            .I(N__32518));
    InMux I__6233 (
            .O(N__32566),
            .I(N__32518));
    InMux I__6232 (
            .O(N__32565),
            .I(N__32518));
    InMux I__6231 (
            .O(N__32564),
            .I(N__32518));
    InMux I__6230 (
            .O(N__32563),
            .I(N__32509));
    InMux I__6229 (
            .O(N__32562),
            .I(N__32509));
    InMux I__6228 (
            .O(N__32561),
            .I(N__32509));
    InMux I__6227 (
            .O(N__32560),
            .I(N__32509));
    InMux I__6226 (
            .O(N__32559),
            .I(N__32500));
    InMux I__6225 (
            .O(N__32558),
            .I(N__32500));
    InMux I__6224 (
            .O(N__32557),
            .I(N__32500));
    InMux I__6223 (
            .O(N__32556),
            .I(N__32500));
    LocalMux I__6222 (
            .O(N__32547),
            .I(N__32495));
    LocalMux I__6221 (
            .O(N__32538),
            .I(N__32495));
    Span4Mux_h I__6220 (
            .O(N__32535),
            .I(N__32490));
    Span4Mux_h I__6219 (
            .O(N__32532),
            .I(N__32490));
    LocalMux I__6218 (
            .O(N__32527),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    LocalMux I__6217 (
            .O(N__32518),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    LocalMux I__6216 (
            .O(N__32509),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    LocalMux I__6215 (
            .O(N__32500),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__6214 (
            .O(N__32495),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__6213 (
            .O(N__32490),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    InMux I__6212 (
            .O(N__32477),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    InMux I__6211 (
            .O(N__32474),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    InMux I__6210 (
            .O(N__32471),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    InMux I__6209 (
            .O(N__32468),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    InMux I__6208 (
            .O(N__32465),
            .I(bfn_13_7_0_));
    InMux I__6207 (
            .O(N__32462),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    InMux I__6206 (
            .O(N__32459),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    InMux I__6205 (
            .O(N__32456),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    InMux I__6204 (
            .O(N__32453),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    InMux I__6203 (
            .O(N__32450),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    InMux I__6202 (
            .O(N__32447),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    InMux I__6201 (
            .O(N__32444),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    InMux I__6200 (
            .O(N__32441),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    InMux I__6199 (
            .O(N__32438),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    InMux I__6198 (
            .O(N__32435),
            .I(bfn_13_6_0_));
    InMux I__6197 (
            .O(N__32432),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    InMux I__6196 (
            .O(N__32429),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    InMux I__6195 (
            .O(N__32426),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    InMux I__6194 (
            .O(N__32423),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    InMux I__6193 (
            .O(N__32420),
            .I(N__32415));
    InMux I__6192 (
            .O(N__32419),
            .I(N__32412));
    InMux I__6191 (
            .O(N__32418),
            .I(N__32409));
    LocalMux I__6190 (
            .O(N__32415),
            .I(N__32403));
    LocalMux I__6189 (
            .O(N__32412),
            .I(N__32403));
    LocalMux I__6188 (
            .O(N__32409),
            .I(N__32400));
    InMux I__6187 (
            .O(N__32408),
            .I(N__32395));
    Span4Mux_h I__6186 (
            .O(N__32403),
            .I(N__32392));
    Span12Mux_h I__6185 (
            .O(N__32400),
            .I(N__32389));
    InMux I__6184 (
            .O(N__32399),
            .I(N__32386));
    InMux I__6183 (
            .O(N__32398),
            .I(N__32383));
    LocalMux I__6182 (
            .O(N__32395),
            .I(N__32378));
    Span4Mux_h I__6181 (
            .O(N__32392),
            .I(N__32378));
    Odrv12 I__6180 (
            .O(N__32389),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    LocalMux I__6179 (
            .O(N__32386),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    LocalMux I__6178 (
            .O(N__32383),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv4 I__6177 (
            .O(N__32378),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    InMux I__6176 (
            .O(N__32369),
            .I(N__32363));
    InMux I__6175 (
            .O(N__32368),
            .I(N__32363));
    LocalMux I__6174 (
            .O(N__32363),
            .I(N__32358));
    InMux I__6173 (
            .O(N__32362),
            .I(N__32353));
    InMux I__6172 (
            .O(N__32361),
            .I(N__32353));
    Odrv4 I__6171 (
            .O(N__32358),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    LocalMux I__6170 (
            .O(N__32353),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    IoInMux I__6169 (
            .O(N__32348),
            .I(N__32345));
    LocalMux I__6168 (
            .O(N__32345),
            .I(N__32342));
    Span4Mux_s3_v I__6167 (
            .O(N__32342),
            .I(N__32339));
    Span4Mux_v I__6166 (
            .O(N__32339),
            .I(N__32336));
    Span4Mux_v I__6165 (
            .O(N__32336),
            .I(N__32332));
    InMux I__6164 (
            .O(N__32335),
            .I(N__32329));
    Odrv4 I__6163 (
            .O(N__32332),
            .I(T45_c));
    LocalMux I__6162 (
            .O(N__32329),
            .I(T45_c));
    InMux I__6161 (
            .O(N__32324),
            .I(N__32321));
    LocalMux I__6160 (
            .O(N__32321),
            .I(N__32318));
    Span12Mux_v I__6159 (
            .O(N__32318),
            .I(N__32315));
    Odrv12 I__6158 (
            .O(N__32315),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ));
    CEMux I__6157 (
            .O(N__32312),
            .I(N__32308));
    CEMux I__6156 (
            .O(N__32311),
            .I(N__32304));
    LocalMux I__6155 (
            .O(N__32308),
            .I(N__32301));
    CEMux I__6154 (
            .O(N__32307),
            .I(N__32298));
    LocalMux I__6153 (
            .O(N__32304),
            .I(N__32295));
    Span4Mux_h I__6152 (
            .O(N__32301),
            .I(N__32289));
    LocalMux I__6151 (
            .O(N__32298),
            .I(N__32289));
    Span4Mux_v I__6150 (
            .O(N__32295),
            .I(N__32286));
    CEMux I__6149 (
            .O(N__32294),
            .I(N__32283));
    Odrv4 I__6148 (
            .O(N__32289),
            .I(\delay_measurement_inst.delay_hc_timer.N_433_i ));
    Odrv4 I__6147 (
            .O(N__32286),
            .I(\delay_measurement_inst.delay_hc_timer.N_433_i ));
    LocalMux I__6146 (
            .O(N__32283),
            .I(\delay_measurement_inst.delay_hc_timer.N_433_i ));
    InMux I__6145 (
            .O(N__32276),
            .I(N__32272));
    InMux I__6144 (
            .O(N__32275),
            .I(N__32269));
    LocalMux I__6143 (
            .O(N__32272),
            .I(N__32262));
    LocalMux I__6142 (
            .O(N__32269),
            .I(N__32262));
    InMux I__6141 (
            .O(N__32268),
            .I(N__32259));
    InMux I__6140 (
            .O(N__32267),
            .I(N__32256));
    Span12Mux_v I__6139 (
            .O(N__32262),
            .I(N__32253));
    LocalMux I__6138 (
            .O(N__32259),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    LocalMux I__6137 (
            .O(N__32256),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    Odrv12 I__6136 (
            .O(N__32253),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    InMux I__6135 (
            .O(N__32246),
            .I(N__32241));
    InMux I__6134 (
            .O(N__32245),
            .I(N__32238));
    InMux I__6133 (
            .O(N__32244),
            .I(N__32235));
    LocalMux I__6132 (
            .O(N__32241),
            .I(N__32232));
    LocalMux I__6131 (
            .O(N__32238),
            .I(N__32225));
    LocalMux I__6130 (
            .O(N__32235),
            .I(N__32225));
    Sp12to4 I__6129 (
            .O(N__32232),
            .I(N__32225));
    Span12Mux_v I__6128 (
            .O(N__32225),
            .I(N__32222));
    Odrv12 I__6127 (
            .O(N__32222),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    InMux I__6126 (
            .O(N__32219),
            .I(N__32213));
    InMux I__6125 (
            .O(N__32218),
            .I(N__32210));
    InMux I__6124 (
            .O(N__32217),
            .I(N__32207));
    InMux I__6123 (
            .O(N__32216),
            .I(N__32204));
    LocalMux I__6122 (
            .O(N__32213),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__6121 (
            .O(N__32210),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__6120 (
            .O(N__32207),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__6119 (
            .O(N__32204),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    InMux I__6118 (
            .O(N__32195),
            .I(bfn_13_5_0_));
    InMux I__6117 (
            .O(N__32192),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    InMux I__6116 (
            .O(N__32189),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    InMux I__6115 (
            .O(N__32186),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    IoInMux I__6114 (
            .O(N__32183),
            .I(N__32180));
    LocalMux I__6113 (
            .O(N__32180),
            .I(N__32177));
    IoSpan4Mux I__6112 (
            .O(N__32177),
            .I(N__32174));
    Span4Mux_s1_v I__6111 (
            .O(N__32174),
            .I(N__32171));
    Sp12to4 I__6110 (
            .O(N__32171),
            .I(N__32168));
    Span12Mux_v I__6109 (
            .O(N__32168),
            .I(N__32164));
    InMux I__6108 (
            .O(N__32167),
            .I(N__32161));
    Odrv12 I__6107 (
            .O(N__32164),
            .I(T12_c));
    LocalMux I__6106 (
            .O(N__32161),
            .I(T12_c));
    InMux I__6105 (
            .O(N__32156),
            .I(N__32153));
    LocalMux I__6104 (
            .O(N__32153),
            .I(N__32150));
    Span4Mux_v I__6103 (
            .O(N__32150),
            .I(N__32145));
    InMux I__6102 (
            .O(N__32149),
            .I(N__32140));
    InMux I__6101 (
            .O(N__32148),
            .I(N__32140));
    Sp12to4 I__6100 (
            .O(N__32145),
            .I(N__32133));
    LocalMux I__6099 (
            .O(N__32140),
            .I(N__32133));
    InMux I__6098 (
            .O(N__32139),
            .I(N__32128));
    InMux I__6097 (
            .O(N__32138),
            .I(N__32128));
    Odrv12 I__6096 (
            .O(N__32133),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    LocalMux I__6095 (
            .O(N__32128),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    CascadeMux I__6094 (
            .O(N__32123),
            .I(N__32120));
    InMux I__6093 (
            .O(N__32120),
            .I(N__32117));
    LocalMux I__6092 (
            .O(N__32117),
            .I(N__32114));
    Span4Mux_h I__6091 (
            .O(N__32114),
            .I(N__32108));
    InMux I__6090 (
            .O(N__32113),
            .I(N__32105));
    InMux I__6089 (
            .O(N__32112),
            .I(N__32102));
    InMux I__6088 (
            .O(N__32111),
            .I(N__32099));
    Span4Mux_h I__6087 (
            .O(N__32108),
            .I(N__32096));
    LocalMux I__6086 (
            .O(N__32105),
            .I(N__32091));
    LocalMux I__6085 (
            .O(N__32102),
            .I(N__32091));
    LocalMux I__6084 (
            .O(N__32099),
            .I(\phase_controller_inst2.hc_time_passed ));
    Odrv4 I__6083 (
            .O(N__32096),
            .I(\phase_controller_inst2.hc_time_passed ));
    Odrv4 I__6082 (
            .O(N__32091),
            .I(\phase_controller_inst2.hc_time_passed ));
    InMux I__6081 (
            .O(N__32084),
            .I(N__32081));
    LocalMux I__6080 (
            .O(N__32081),
            .I(N__32078));
    Span4Mux_v I__6079 (
            .O(N__32078),
            .I(N__32075));
    Span4Mux_v I__6078 (
            .O(N__32075),
            .I(N__32071));
    CascadeMux I__6077 (
            .O(N__32074),
            .I(N__32068));
    Sp12to4 I__6076 (
            .O(N__32071),
            .I(N__32064));
    InMux I__6075 (
            .O(N__32068),
            .I(N__32059));
    InMux I__6074 (
            .O(N__32067),
            .I(N__32059));
    Span12Mux_h I__6073 (
            .O(N__32064),
            .I(N__32054));
    LocalMux I__6072 (
            .O(N__32059),
            .I(N__32054));
    Span12Mux_v I__6071 (
            .O(N__32054),
            .I(N__32051));
    Odrv12 I__6070 (
            .O(N__32051),
            .I(il_max_comp2_D2));
    CascadeMux I__6069 (
            .O(N__32048),
            .I(\phase_controller_inst2.time_passed_RNI9M3O_cascade_ ));
    InMux I__6068 (
            .O(N__32045),
            .I(N__32042));
    LocalMux I__6067 (
            .O(N__32042),
            .I(\phase_controller_inst2.time_passed_RNI9M3O ));
    IoInMux I__6066 (
            .O(N__32039),
            .I(N__32036));
    LocalMux I__6065 (
            .O(N__32036),
            .I(N__32033));
    Span4Mux_s3_v I__6064 (
            .O(N__32033),
            .I(N__32030));
    Span4Mux_h I__6063 (
            .O(N__32030),
            .I(N__32027));
    Span4Mux_v I__6062 (
            .O(N__32027),
            .I(N__32024));
    Span4Mux_v I__6061 (
            .O(N__32024),
            .I(N__32020));
    InMux I__6060 (
            .O(N__32023),
            .I(N__32017));
    Odrv4 I__6059 (
            .O(N__32020),
            .I(T23_c));
    LocalMux I__6058 (
            .O(N__32017),
            .I(T23_c));
    CascadeMux I__6057 (
            .O(N__32012),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_6_cascade_ ));
    InMux I__6056 (
            .O(N__32009),
            .I(N__32006));
    LocalMux I__6055 (
            .O(N__32006),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_5 ));
    InMux I__6054 (
            .O(N__32003),
            .I(N__31998));
    InMux I__6053 (
            .O(N__32002),
            .I(N__31993));
    InMux I__6052 (
            .O(N__32001),
            .I(N__31993));
    LocalMux I__6051 (
            .O(N__31998),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17 ));
    LocalMux I__6050 (
            .O(N__31993),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17 ));
    CascadeMux I__6049 (
            .O(N__31988),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17_cascade_ ));
    InMux I__6048 (
            .O(N__31985),
            .I(N__31982));
    LocalMux I__6047 (
            .O(N__31982),
            .I(N__31979));
    Span4Mux_h I__6046 (
            .O(N__31979),
            .I(N__31976));
    Odrv4 I__6045 (
            .O(N__31976),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58FZ0Z_31 ));
    InMux I__6044 (
            .O(N__31973),
            .I(N__31968));
    InMux I__6043 (
            .O(N__31972),
            .I(N__31963));
    InMux I__6042 (
            .O(N__31971),
            .I(N__31963));
    LocalMux I__6041 (
            .O(N__31968),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    LocalMux I__6040 (
            .O(N__31963),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    CascadeMux I__6039 (
            .O(N__31958),
            .I(N__31955));
    InMux I__6038 (
            .O(N__31955),
            .I(N__31952));
    LocalMux I__6037 (
            .O(N__31952),
            .I(N__31947));
    InMux I__6036 (
            .O(N__31951),
            .I(N__31944));
    InMux I__6035 (
            .O(N__31950),
            .I(N__31941));
    Odrv4 I__6034 (
            .O(N__31947),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    LocalMux I__6033 (
            .O(N__31944),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    LocalMux I__6032 (
            .O(N__31941),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    InMux I__6031 (
            .O(N__31934),
            .I(N__31930));
    CascadeMux I__6030 (
            .O(N__31933),
            .I(N__31927));
    LocalMux I__6029 (
            .O(N__31930),
            .I(N__31923));
    InMux I__6028 (
            .O(N__31927),
            .I(N__31920));
    InMux I__6027 (
            .O(N__31926),
            .I(N__31917));
    Span4Mux_v I__6026 (
            .O(N__31923),
            .I(N__31914));
    LocalMux I__6025 (
            .O(N__31920),
            .I(N__31911));
    LocalMux I__6024 (
            .O(N__31917),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    Odrv4 I__6023 (
            .O(N__31914),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    Odrv4 I__6022 (
            .O(N__31911),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    InMux I__6021 (
            .O(N__31904),
            .I(N__31901));
    LocalMux I__6020 (
            .O(N__31901),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16 ));
    InMux I__6019 (
            .O(N__31898),
            .I(N__31895));
    LocalMux I__6018 (
            .O(N__31895),
            .I(N__31891));
    InMux I__6017 (
            .O(N__31894),
            .I(N__31888));
    Span4Mux_h I__6016 (
            .O(N__31891),
            .I(N__31881));
    LocalMux I__6015 (
            .O(N__31888),
            .I(N__31881));
    InMux I__6014 (
            .O(N__31887),
            .I(N__31876));
    InMux I__6013 (
            .O(N__31886),
            .I(N__31876));
    Odrv4 I__6012 (
            .O(N__31881),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto14 ));
    LocalMux I__6011 (
            .O(N__31876),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto14 ));
    CascadeMux I__6010 (
            .O(N__31871),
            .I(N__31868));
    InMux I__6009 (
            .O(N__31868),
            .I(N__31865));
    LocalMux I__6008 (
            .O(N__31865),
            .I(N__31862));
    Span4Mux_v I__6007 (
            .O(N__31862),
            .I(N__31857));
    InMux I__6006 (
            .O(N__31861),
            .I(N__31852));
    InMux I__6005 (
            .O(N__31860),
            .I(N__31852));
    Odrv4 I__6004 (
            .O(N__31857),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto6 ));
    LocalMux I__6003 (
            .O(N__31852),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto6 ));
    CascadeMux I__6002 (
            .O(N__31847),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16_cascade_ ));
    CascadeMux I__6001 (
            .O(N__31844),
            .I(N__31841));
    InMux I__6000 (
            .O(N__31841),
            .I(N__31838));
    LocalMux I__5999 (
            .O(N__31838),
            .I(N__31834));
    InMux I__5998 (
            .O(N__31837),
            .I(N__31830));
    Span4Mux_h I__5997 (
            .O(N__31834),
            .I(N__31827));
    InMux I__5996 (
            .O(N__31833),
            .I(N__31824));
    LocalMux I__5995 (
            .O(N__31830),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6 ));
    Odrv4 I__5994 (
            .O(N__31827),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6 ));
    LocalMux I__5993 (
            .O(N__31824),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6 ));
    InMux I__5992 (
            .O(N__31817),
            .I(N__31814));
    LocalMux I__5991 (
            .O(N__31814),
            .I(N__31809));
    InMux I__5990 (
            .O(N__31813),
            .I(N__31806));
    InMux I__5989 (
            .O(N__31812),
            .I(N__31803));
    Odrv4 I__5988 (
            .O(N__31809),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15 ));
    LocalMux I__5987 (
            .O(N__31806),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15 ));
    LocalMux I__5986 (
            .O(N__31803),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15 ));
    CascadeMux I__5985 (
            .O(N__31796),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6_cascade_ ));
    InMux I__5984 (
            .O(N__31793),
            .I(N__31788));
    CascadeMux I__5983 (
            .O(N__31792),
            .I(N__31783));
    InMux I__5982 (
            .O(N__31791),
            .I(N__31780));
    LocalMux I__5981 (
            .O(N__31788),
            .I(N__31777));
    InMux I__5980 (
            .O(N__31787),
            .I(N__31772));
    InMux I__5979 (
            .O(N__31786),
            .I(N__31772));
    InMux I__5978 (
            .O(N__31783),
            .I(N__31768));
    LocalMux I__5977 (
            .O(N__31780),
            .I(N__31765));
    Span4Mux_h I__5976 (
            .O(N__31777),
            .I(N__31762));
    LocalMux I__5975 (
            .O(N__31772),
            .I(N__31759));
    InMux I__5974 (
            .O(N__31771),
            .I(N__31756));
    LocalMux I__5973 (
            .O(N__31768),
            .I(N__31753));
    Span4Mux_h I__5972 (
            .O(N__31765),
            .I(N__31750));
    Span4Mux_v I__5971 (
            .O(N__31762),
            .I(N__31747));
    Span4Mux_h I__5970 (
            .O(N__31759),
            .I(N__31740));
    LocalMux I__5969 (
            .O(N__31756),
            .I(N__31740));
    Span4Mux_h I__5968 (
            .O(N__31753),
            .I(N__31740));
    Odrv4 I__5967 (
            .O(N__31750),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    Odrv4 I__5966 (
            .O(N__31747),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    Odrv4 I__5965 (
            .O(N__31740),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    InMux I__5964 (
            .O(N__31733),
            .I(N__31729));
    InMux I__5963 (
            .O(N__31732),
            .I(N__31726));
    LocalMux I__5962 (
            .O(N__31729),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31 ));
    LocalMux I__5961 (
            .O(N__31726),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31 ));
    CascadeMux I__5960 (
            .O(N__31721),
            .I(N__31718));
    InMux I__5959 (
            .O(N__31718),
            .I(N__31715));
    LocalMux I__5958 (
            .O(N__31715),
            .I(N__31711));
    InMux I__5957 (
            .O(N__31714),
            .I(N__31708));
    Odrv4 I__5956 (
            .O(N__31711),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    LocalMux I__5955 (
            .O(N__31708),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    CascadeMux I__5954 (
            .O(N__31703),
            .I(N__31700));
    InMux I__5953 (
            .O(N__31700),
            .I(N__31697));
    LocalMux I__5952 (
            .O(N__31697),
            .I(N__31694));
    Span4Mux_v I__5951 (
            .O(N__31694),
            .I(N__31690));
    InMux I__5950 (
            .O(N__31693),
            .I(N__31687));
    Odrv4 I__5949 (
            .O(N__31690),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    LocalMux I__5948 (
            .O(N__31687),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    InMux I__5947 (
            .O(N__31682),
            .I(N__31676));
    InMux I__5946 (
            .O(N__31681),
            .I(N__31676));
    LocalMux I__5945 (
            .O(N__31676),
            .I(N__31672));
    CascadeMux I__5944 (
            .O(N__31675),
            .I(N__31669));
    Span4Mux_v I__5943 (
            .O(N__31672),
            .I(N__31666));
    InMux I__5942 (
            .O(N__31669),
            .I(N__31663));
    Odrv4 I__5941 (
            .O(N__31666),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2 ));
    LocalMux I__5940 (
            .O(N__31663),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2 ));
    IoInMux I__5939 (
            .O(N__31658),
            .I(N__31655));
    LocalMux I__5938 (
            .O(N__31655),
            .I(N__31652));
    Span4Mux_s2_v I__5937 (
            .O(N__31652),
            .I(N__31649));
    Sp12to4 I__5936 (
            .O(N__31649),
            .I(N__31646));
    Span12Mux_h I__5935 (
            .O(N__31646),
            .I(N__31643));
    Span12Mux_v I__5934 (
            .O(N__31643),
            .I(N__31639));
    InMux I__5933 (
            .O(N__31642),
            .I(N__31636));
    Odrv12 I__5932 (
            .O(N__31639),
            .I(T01_c));
    LocalMux I__5931 (
            .O(N__31636),
            .I(T01_c));
    CascadeMux I__5930 (
            .O(N__31631),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15_cascade_ ));
    InMux I__5929 (
            .O(N__31628),
            .I(N__31625));
    LocalMux I__5928 (
            .O(N__31625),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKRZ0Z_2 ));
    CascadeMux I__5927 (
            .O(N__31622),
            .I(N__31619));
    InMux I__5926 (
            .O(N__31619),
            .I(N__31616));
    LocalMux I__5925 (
            .O(N__31616),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847Z0Z_31 ));
    CascadeMux I__5924 (
            .O(N__31613),
            .I(N__31610));
    InMux I__5923 (
            .O(N__31610),
            .I(N__31607));
    LocalMux I__5922 (
            .O(N__31607),
            .I(N__31604));
    Span4Mux_h I__5921 (
            .O(N__31604),
            .I(N__31600));
    InMux I__5920 (
            .O(N__31603),
            .I(N__31597));
    Odrv4 I__5919 (
            .O(N__31600),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    LocalMux I__5918 (
            .O(N__31597),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    InMux I__5917 (
            .O(N__31592),
            .I(N__31588));
    InMux I__5916 (
            .O(N__31591),
            .I(N__31585));
    LocalMux I__5915 (
            .O(N__31588),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    LocalMux I__5914 (
            .O(N__31585),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    InMux I__5913 (
            .O(N__31580),
            .I(N__31577));
    LocalMux I__5912 (
            .O(N__31577),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4 ));
    CascadeMux I__5911 (
            .O(N__31574),
            .I(N__31570));
    InMux I__5910 (
            .O(N__31573),
            .I(N__31567));
    InMux I__5909 (
            .O(N__31570),
            .I(N__31564));
    LocalMux I__5908 (
            .O(N__31567),
            .I(N__31561));
    LocalMux I__5907 (
            .O(N__31564),
            .I(N__31558));
    Span4Mux_v I__5906 (
            .O(N__31561),
            .I(N__31555));
    Odrv4 I__5905 (
            .O(N__31558),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    Odrv4 I__5904 (
            .O(N__31555),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    CascadeMux I__5903 (
            .O(N__31550),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4_cascade_ ));
    InMux I__5902 (
            .O(N__31547),
            .I(N__31544));
    LocalMux I__5901 (
            .O(N__31544),
            .I(N__31541));
    Span4Mux_v I__5900 (
            .O(N__31541),
            .I(N__31536));
    InMux I__5899 (
            .O(N__31540),
            .I(N__31531));
    InMux I__5898 (
            .O(N__31539),
            .I(N__31531));
    Odrv4 I__5897 (
            .O(N__31536),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    LocalMux I__5896 (
            .O(N__31531),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    InMux I__5895 (
            .O(N__31526),
            .I(N__31523));
    LocalMux I__5894 (
            .O(N__31523),
            .I(N__31520));
    Span4Mux_h I__5893 (
            .O(N__31520),
            .I(N__31516));
    InMux I__5892 (
            .O(N__31519),
            .I(N__31513));
    Odrv4 I__5891 (
            .O(N__31516),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1 ));
    LocalMux I__5890 (
            .O(N__31513),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1 ));
    CascadeMux I__5889 (
            .O(N__31508),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1_cascade_ ));
    InMux I__5888 (
            .O(N__31505),
            .I(N__31502));
    LocalMux I__5887 (
            .O(N__31502),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4Z0Z_31 ));
    CascadeMux I__5886 (
            .O(N__31499),
            .I(N__31496));
    InMux I__5885 (
            .O(N__31496),
            .I(N__31492));
    InMux I__5884 (
            .O(N__31495),
            .I(N__31489));
    LocalMux I__5883 (
            .O(N__31492),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    LocalMux I__5882 (
            .O(N__31489),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    InMux I__5881 (
            .O(N__31484),
            .I(N__31481));
    LocalMux I__5880 (
            .O(N__31481),
            .I(N__31477));
    InMux I__5879 (
            .O(N__31480),
            .I(N__31474));
    Odrv4 I__5878 (
            .O(N__31477),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    LocalMux I__5877 (
            .O(N__31474),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    CascadeMux I__5876 (
            .O(N__31469),
            .I(N__31466));
    InMux I__5875 (
            .O(N__31466),
            .I(N__31463));
    LocalMux I__5874 (
            .O(N__31463),
            .I(N__31459));
    CascadeMux I__5873 (
            .O(N__31462),
            .I(N__31456));
    Span4Mux_h I__5872 (
            .O(N__31459),
            .I(N__31453));
    InMux I__5871 (
            .O(N__31456),
            .I(N__31450));
    Odrv4 I__5870 (
            .O(N__31453),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    LocalMux I__5869 (
            .O(N__31450),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    CascadeMux I__5868 (
            .O(N__31445),
            .I(N__31442));
    InMux I__5867 (
            .O(N__31442),
            .I(N__31439));
    LocalMux I__5866 (
            .O(N__31439),
            .I(N__31435));
    InMux I__5865 (
            .O(N__31438),
            .I(N__31432));
    Odrv4 I__5864 (
            .O(N__31435),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    LocalMux I__5863 (
            .O(N__31432),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    CascadeMux I__5862 (
            .O(N__31427),
            .I(N__31424));
    InMux I__5861 (
            .O(N__31424),
            .I(N__31420));
    InMux I__5860 (
            .O(N__31423),
            .I(N__31417));
    LocalMux I__5859 (
            .O(N__31420),
            .I(N__31414));
    LocalMux I__5858 (
            .O(N__31417),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10 ));
    Odrv4 I__5857 (
            .O(N__31414),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10 ));
    InMux I__5856 (
            .O(N__31409),
            .I(N__31406));
    LocalMux I__5855 (
            .O(N__31406),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15 ));
    InMux I__5854 (
            .O(N__31403),
            .I(N__31400));
    LocalMux I__5853 (
            .O(N__31400),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_a3_1_3 ));
    InMux I__5852 (
            .O(N__31397),
            .I(N__31394));
    LocalMux I__5851 (
            .O(N__31394),
            .I(N__31391));
    Odrv4 I__5850 (
            .O(N__31391),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ));
    InMux I__5849 (
            .O(N__31388),
            .I(N__31385));
    LocalMux I__5848 (
            .O(N__31385),
            .I(N__31380));
    CascadeMux I__5847 (
            .O(N__31384),
            .I(N__31377));
    InMux I__5846 (
            .O(N__31383),
            .I(N__31374));
    Span4Mux_h I__5845 (
            .O(N__31380),
            .I(N__31371));
    InMux I__5844 (
            .O(N__31377),
            .I(N__31368));
    LocalMux I__5843 (
            .O(N__31374),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ));
    Odrv4 I__5842 (
            .O(N__31371),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ));
    LocalMux I__5841 (
            .O(N__31368),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ));
    InMux I__5840 (
            .O(N__31361),
            .I(N__31358));
    LocalMux I__5839 (
            .O(N__31358),
            .I(N__31354));
    InMux I__5838 (
            .O(N__31357),
            .I(N__31350));
    Span4Mux_v I__5837 (
            .O(N__31354),
            .I(N__31347));
    InMux I__5836 (
            .O(N__31353),
            .I(N__31344));
    LocalMux I__5835 (
            .O(N__31350),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ));
    Odrv4 I__5834 (
            .O(N__31347),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ));
    LocalMux I__5833 (
            .O(N__31344),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ));
    CascadeMux I__5832 (
            .O(N__31337),
            .I(N__31334));
    InMux I__5831 (
            .O(N__31334),
            .I(N__31330));
    InMux I__5830 (
            .O(N__31333),
            .I(N__31326));
    LocalMux I__5829 (
            .O(N__31330),
            .I(N__31323));
    InMux I__5828 (
            .O(N__31329),
            .I(N__31320));
    LocalMux I__5827 (
            .O(N__31326),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ));
    Odrv4 I__5826 (
            .O(N__31323),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ));
    LocalMux I__5825 (
            .O(N__31320),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ));
    InMux I__5824 (
            .O(N__31313),
            .I(N__31310));
    LocalMux I__5823 (
            .O(N__31310),
            .I(N__31306));
    InMux I__5822 (
            .O(N__31309),
            .I(N__31302));
    Span4Mux_h I__5821 (
            .O(N__31306),
            .I(N__31299));
    InMux I__5820 (
            .O(N__31305),
            .I(N__31296));
    LocalMux I__5819 (
            .O(N__31302),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ));
    Odrv4 I__5818 (
            .O(N__31299),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ));
    LocalMux I__5817 (
            .O(N__31296),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ));
    InMux I__5816 (
            .O(N__31289),
            .I(N__31286));
    LocalMux I__5815 (
            .O(N__31286),
            .I(N__31282));
    InMux I__5814 (
            .O(N__31285),
            .I(N__31278));
    Span4Mux_h I__5813 (
            .O(N__31282),
            .I(N__31275));
    InMux I__5812 (
            .O(N__31281),
            .I(N__31272));
    LocalMux I__5811 (
            .O(N__31278),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ));
    Odrv4 I__5810 (
            .O(N__31275),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ));
    LocalMux I__5809 (
            .O(N__31272),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ));
    InMux I__5808 (
            .O(N__31265),
            .I(N__31262));
    LocalMux I__5807 (
            .O(N__31262),
            .I(N__31259));
    Odrv4 I__5806 (
            .O(N__31259),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ));
    CascadeMux I__5805 (
            .O(N__31256),
            .I(N__31253));
    InMux I__5804 (
            .O(N__31253),
            .I(N__31250));
    LocalMux I__5803 (
            .O(N__31250),
            .I(N__31247));
    Span4Mux_h I__5802 (
            .O(N__31247),
            .I(N__31242));
    InMux I__5801 (
            .O(N__31246),
            .I(N__31239));
    InMux I__5800 (
            .O(N__31245),
            .I(N__31236));
    Span4Mux_h I__5799 (
            .O(N__31242),
            .I(N__31232));
    LocalMux I__5798 (
            .O(N__31239),
            .I(N__31227));
    LocalMux I__5797 (
            .O(N__31236),
            .I(N__31227));
    InMux I__5796 (
            .O(N__31235),
            .I(N__31224));
    Span4Mux_h I__5795 (
            .O(N__31232),
            .I(N__31221));
    Span4Mux_v I__5794 (
            .O(N__31227),
            .I(N__31218));
    LocalMux I__5793 (
            .O(N__31224),
            .I(elapsed_time_ns_1_RNIO0MD11_0_11));
    Odrv4 I__5792 (
            .O(N__31221),
            .I(elapsed_time_ns_1_RNIO0MD11_0_11));
    Odrv4 I__5791 (
            .O(N__31218),
            .I(elapsed_time_ns_1_RNIO0MD11_0_11));
    InMux I__5790 (
            .O(N__31211),
            .I(N__31206));
    InMux I__5789 (
            .O(N__31210),
            .I(N__31203));
    InMux I__5788 (
            .O(N__31209),
            .I(N__31200));
    LocalMux I__5787 (
            .O(N__31206),
            .I(N__31197));
    LocalMux I__5786 (
            .O(N__31203),
            .I(N__31192));
    LocalMux I__5785 (
            .O(N__31200),
            .I(N__31192));
    Odrv4 I__5784 (
            .O(N__31197),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto15 ));
    Odrv4 I__5783 (
            .O(N__31192),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto15 ));
    InMux I__5782 (
            .O(N__31187),
            .I(N__31184));
    LocalMux I__5781 (
            .O(N__31184),
            .I(N__31179));
    InMux I__5780 (
            .O(N__31183),
            .I(N__31176));
    InMux I__5779 (
            .O(N__31182),
            .I(N__31173));
    Odrv4 I__5778 (
            .O(N__31179),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    LocalMux I__5777 (
            .O(N__31176),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    LocalMux I__5776 (
            .O(N__31173),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    InMux I__5775 (
            .O(N__31166),
            .I(N__31163));
    LocalMux I__5774 (
            .O(N__31163),
            .I(N__31158));
    InMux I__5773 (
            .O(N__31162),
            .I(N__31155));
    InMux I__5772 (
            .O(N__31161),
            .I(N__31152));
    Odrv4 I__5771 (
            .O(N__31158),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    LocalMux I__5770 (
            .O(N__31155),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    LocalMux I__5769 (
            .O(N__31152),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    InMux I__5768 (
            .O(N__31145),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ));
    InMux I__5767 (
            .O(N__31142),
            .I(bfn_12_12_0_));
    InMux I__5766 (
            .O(N__31139),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ));
    InMux I__5765 (
            .O(N__31136),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ));
    InMux I__5764 (
            .O(N__31133),
            .I(N__31129));
    CascadeMux I__5763 (
            .O(N__31132),
            .I(N__31126));
    LocalMux I__5762 (
            .O(N__31129),
            .I(N__31123));
    InMux I__5761 (
            .O(N__31126),
            .I(N__31120));
    Span4Mux_v I__5760 (
            .O(N__31123),
            .I(N__31114));
    LocalMux I__5759 (
            .O(N__31120),
            .I(N__31114));
    InMux I__5758 (
            .O(N__31119),
            .I(N__31111));
    Span4Mux_h I__5757 (
            .O(N__31114),
            .I(N__31108));
    LocalMux I__5756 (
            .O(N__31111),
            .I(N__31105));
    Odrv4 I__5755 (
            .O(N__31108),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    Odrv4 I__5754 (
            .O(N__31105),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    InMux I__5753 (
            .O(N__31100),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ));
    InMux I__5752 (
            .O(N__31097),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ));
    InMux I__5751 (
            .O(N__31094),
            .I(N__31091));
    LocalMux I__5750 (
            .O(N__31091),
            .I(N__31087));
    InMux I__5749 (
            .O(N__31090),
            .I(N__31084));
    Span4Mux_v I__5748 (
            .O(N__31087),
            .I(N__31079));
    LocalMux I__5747 (
            .O(N__31084),
            .I(N__31079));
    Span4Mux_h I__5746 (
            .O(N__31079),
            .I(N__31075));
    InMux I__5745 (
            .O(N__31078),
            .I(N__31072));
    Odrv4 I__5744 (
            .O(N__31075),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    LocalMux I__5743 (
            .O(N__31072),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    InMux I__5742 (
            .O(N__31067),
            .I(N__31064));
    LocalMux I__5741 (
            .O(N__31064),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ));
    InMux I__5740 (
            .O(N__31061),
            .I(N__31058));
    LocalMux I__5739 (
            .O(N__31058),
            .I(N__31054));
    InMux I__5738 (
            .O(N__31057),
            .I(N__31051));
    Span4Mux_v I__5737 (
            .O(N__31054),
            .I(N__31046));
    LocalMux I__5736 (
            .O(N__31051),
            .I(N__31046));
    Span4Mux_h I__5735 (
            .O(N__31046),
            .I(N__31042));
    InMux I__5734 (
            .O(N__31045),
            .I(N__31039));
    Odrv4 I__5733 (
            .O(N__31042),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    LocalMux I__5732 (
            .O(N__31039),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    InMux I__5731 (
            .O(N__31034),
            .I(N__31031));
    LocalMux I__5730 (
            .O(N__31031),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ));
    InMux I__5729 (
            .O(N__31028),
            .I(N__31025));
    LocalMux I__5728 (
            .O(N__31025),
            .I(N__31021));
    InMux I__5727 (
            .O(N__31024),
            .I(N__31018));
    Span4Mux_v I__5726 (
            .O(N__31021),
            .I(N__31013));
    LocalMux I__5725 (
            .O(N__31018),
            .I(N__31013));
    Span4Mux_h I__5724 (
            .O(N__31013),
            .I(N__31009));
    InMux I__5723 (
            .O(N__31012),
            .I(N__31006));
    Odrv4 I__5722 (
            .O(N__31009),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    LocalMux I__5721 (
            .O(N__31006),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    InMux I__5720 (
            .O(N__31001),
            .I(N__30998));
    LocalMux I__5719 (
            .O(N__30998),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ));
    InMux I__5718 (
            .O(N__30995),
            .I(N__30992));
    LocalMux I__5717 (
            .O(N__30992),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ));
    InMux I__5716 (
            .O(N__30989),
            .I(N__30986));
    LocalMux I__5715 (
            .O(N__30986),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ));
    InMux I__5714 (
            .O(N__30983),
            .I(N__30980));
    LocalMux I__5713 (
            .O(N__30980),
            .I(N__30976));
    InMux I__5712 (
            .O(N__30979),
            .I(N__30973));
    Odrv4 I__5711 (
            .O(N__30976),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    LocalMux I__5710 (
            .O(N__30973),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    InMux I__5709 (
            .O(N__30968),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ));
    InMux I__5708 (
            .O(N__30965),
            .I(N__30962));
    LocalMux I__5707 (
            .O(N__30962),
            .I(N__30958));
    InMux I__5706 (
            .O(N__30961),
            .I(N__30955));
    Odrv4 I__5705 (
            .O(N__30958),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    LocalMux I__5704 (
            .O(N__30955),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    InMux I__5703 (
            .O(N__30950),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ));
    InMux I__5702 (
            .O(N__30947),
            .I(N__30944));
    LocalMux I__5701 (
            .O(N__30944),
            .I(N__30941));
    Span4Mux_v I__5700 (
            .O(N__30941),
            .I(N__30938));
    Span4Mux_h I__5699 (
            .O(N__30938),
            .I(N__30934));
    InMux I__5698 (
            .O(N__30937),
            .I(N__30931));
    Odrv4 I__5697 (
            .O(N__30934),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    LocalMux I__5696 (
            .O(N__30931),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    InMux I__5695 (
            .O(N__30926),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ));
    CascadeMux I__5694 (
            .O(N__30923),
            .I(N__30919));
    InMux I__5693 (
            .O(N__30922),
            .I(N__30916));
    InMux I__5692 (
            .O(N__30919),
            .I(N__30913));
    LocalMux I__5691 (
            .O(N__30916),
            .I(N__30908));
    LocalMux I__5690 (
            .O(N__30913),
            .I(N__30908));
    Span4Mux_h I__5689 (
            .O(N__30908),
            .I(N__30904));
    InMux I__5688 (
            .O(N__30907),
            .I(N__30901));
    Odrv4 I__5687 (
            .O(N__30904),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    LocalMux I__5686 (
            .O(N__30901),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    InMux I__5685 (
            .O(N__30896),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ));
    InMux I__5684 (
            .O(N__30893),
            .I(N__30889));
    InMux I__5683 (
            .O(N__30892),
            .I(N__30886));
    LocalMux I__5682 (
            .O(N__30889),
            .I(N__30880));
    LocalMux I__5681 (
            .O(N__30886),
            .I(N__30880));
    InMux I__5680 (
            .O(N__30885),
            .I(N__30877));
    Odrv4 I__5679 (
            .O(N__30880),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    LocalMux I__5678 (
            .O(N__30877),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    InMux I__5677 (
            .O(N__30872),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ));
    InMux I__5676 (
            .O(N__30869),
            .I(N__30865));
    CascadeMux I__5675 (
            .O(N__30868),
            .I(N__30862));
    LocalMux I__5674 (
            .O(N__30865),
            .I(N__30859));
    InMux I__5673 (
            .O(N__30862),
            .I(N__30856));
    Span4Mux_h I__5672 (
            .O(N__30859),
            .I(N__30853));
    LocalMux I__5671 (
            .O(N__30856),
            .I(N__30850));
    Span4Mux_h I__5670 (
            .O(N__30853),
            .I(N__30846));
    Span4Mux_h I__5669 (
            .O(N__30850),
            .I(N__30843));
    InMux I__5668 (
            .O(N__30849),
            .I(N__30840));
    Odrv4 I__5667 (
            .O(N__30846),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    Odrv4 I__5666 (
            .O(N__30843),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    LocalMux I__5665 (
            .O(N__30840),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    InMux I__5664 (
            .O(N__30833),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ));
    CascadeMux I__5663 (
            .O(N__30830),
            .I(N__30826));
    InMux I__5662 (
            .O(N__30829),
            .I(N__30823));
    InMux I__5661 (
            .O(N__30826),
            .I(N__30820));
    LocalMux I__5660 (
            .O(N__30823),
            .I(N__30815));
    LocalMux I__5659 (
            .O(N__30820),
            .I(N__30815));
    Span4Mux_h I__5658 (
            .O(N__30815),
            .I(N__30811));
    InMux I__5657 (
            .O(N__30814),
            .I(N__30808));
    Odrv4 I__5656 (
            .O(N__30811),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    LocalMux I__5655 (
            .O(N__30808),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    CascadeMux I__5654 (
            .O(N__30803),
            .I(N__30800));
    InMux I__5653 (
            .O(N__30800),
            .I(N__30797));
    LocalMux I__5652 (
            .O(N__30797),
            .I(N__30794));
    Span12Mux_s8_h I__5651 (
            .O(N__30794),
            .I(N__30791));
    Odrv12 I__5650 (
            .O(N__30791),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ));
    InMux I__5649 (
            .O(N__30788),
            .I(N__30785));
    LocalMux I__5648 (
            .O(N__30785),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ));
    CascadeMux I__5647 (
            .O(N__30782),
            .I(N__30778));
    CascadeMux I__5646 (
            .O(N__30781),
            .I(N__30775));
    InMux I__5645 (
            .O(N__30778),
            .I(N__30772));
    InMux I__5644 (
            .O(N__30775),
            .I(N__30769));
    LocalMux I__5643 (
            .O(N__30772),
            .I(N__30764));
    LocalMux I__5642 (
            .O(N__30769),
            .I(N__30761));
    InMux I__5641 (
            .O(N__30768),
            .I(N__30758));
    InMux I__5640 (
            .O(N__30767),
            .I(N__30755));
    Span4Mux_v I__5639 (
            .O(N__30764),
            .I(N__30752));
    Span4Mux_v I__5638 (
            .O(N__30761),
            .I(N__30747));
    LocalMux I__5637 (
            .O(N__30758),
            .I(N__30747));
    LocalMux I__5636 (
            .O(N__30755),
            .I(N__30741));
    Span4Mux_h I__5635 (
            .O(N__30752),
            .I(N__30741));
    Span4Mux_h I__5634 (
            .O(N__30747),
            .I(N__30738));
    InMux I__5633 (
            .O(N__30746),
            .I(N__30735));
    Odrv4 I__5632 (
            .O(N__30741),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv4 I__5631 (
            .O(N__30738),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    LocalMux I__5630 (
            .O(N__30735),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    InMux I__5629 (
            .O(N__30728),
            .I(N__30725));
    LocalMux I__5628 (
            .O(N__30725),
            .I(N__30722));
    Span4Mux_v I__5627 (
            .O(N__30722),
            .I(N__30719));
    Odrv4 I__5626 (
            .O(N__30719),
            .I(\current_shift_inst.PI_CTRL.integrator_i_8 ));
    InMux I__5625 (
            .O(N__30716),
            .I(N__30713));
    LocalMux I__5624 (
            .O(N__30713),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ));
    InMux I__5623 (
            .O(N__30710),
            .I(N__30707));
    LocalMux I__5622 (
            .O(N__30707),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ));
    InMux I__5621 (
            .O(N__30704),
            .I(N__30701));
    LocalMux I__5620 (
            .O(N__30701),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ));
    InMux I__5619 (
            .O(N__30698),
            .I(N__30693));
    InMux I__5618 (
            .O(N__30697),
            .I(N__30690));
    InMux I__5617 (
            .O(N__30696),
            .I(N__30687));
    LocalMux I__5616 (
            .O(N__30693),
            .I(N__30684));
    LocalMux I__5615 (
            .O(N__30690),
            .I(N__30681));
    LocalMux I__5614 (
            .O(N__30687),
            .I(N__30676));
    Span4Mux_h I__5613 (
            .O(N__30684),
            .I(N__30671));
    Span4Mux_h I__5612 (
            .O(N__30681),
            .I(N__30671));
    InMux I__5611 (
            .O(N__30680),
            .I(N__30668));
    InMux I__5610 (
            .O(N__30679),
            .I(N__30665));
    Span4Mux_v I__5609 (
            .O(N__30676),
            .I(N__30662));
    Odrv4 I__5608 (
            .O(N__30671),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    LocalMux I__5607 (
            .O(N__30668),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    LocalMux I__5606 (
            .O(N__30665),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv4 I__5605 (
            .O(N__30662),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    InMux I__5604 (
            .O(N__30653),
            .I(N__30650));
    LocalMux I__5603 (
            .O(N__30650),
            .I(N__30647));
    Odrv4 I__5602 (
            .O(N__30647),
            .I(\current_shift_inst.PI_CTRL.integrator_i_21 ));
    InMux I__5601 (
            .O(N__30644),
            .I(N__30641));
    LocalMux I__5600 (
            .O(N__30641),
            .I(N__30636));
    InMux I__5599 (
            .O(N__30640),
            .I(N__30633));
    InMux I__5598 (
            .O(N__30639),
            .I(N__30630));
    Span4Mux_h I__5597 (
            .O(N__30636),
            .I(N__30627));
    LocalMux I__5596 (
            .O(N__30633),
            .I(N__30624));
    LocalMux I__5595 (
            .O(N__30630),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ));
    Odrv4 I__5594 (
            .O(N__30627),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ));
    Odrv4 I__5593 (
            .O(N__30624),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ));
    IoInMux I__5592 (
            .O(N__30617),
            .I(N__30614));
    LocalMux I__5591 (
            .O(N__30614),
            .I(N__30611));
    Span4Mux_s2_v I__5590 (
            .O(N__30611),
            .I(N__30608));
    Span4Mux_h I__5589 (
            .O(N__30608),
            .I(N__30605));
    Span4Mux_v I__5588 (
            .O(N__30605),
            .I(N__30602));
    Odrv4 I__5587 (
            .O(N__30602),
            .I(\delay_measurement_inst.delay_hc_timer.N_432_i ));
    InMux I__5586 (
            .O(N__30599),
            .I(N__30596));
    LocalMux I__5585 (
            .O(N__30596),
            .I(N__30593));
    Span4Mux_h I__5584 (
            .O(N__30593),
            .I(N__30590));
    Odrv4 I__5583 (
            .O(N__30590),
            .I(il_min_comp1_c));
    InMux I__5582 (
            .O(N__30587),
            .I(N__30584));
    LocalMux I__5581 (
            .O(N__30584),
            .I(il_min_comp1_D1));
    ClkMux I__5580 (
            .O(N__30581),
            .I(N__30575));
    ClkMux I__5579 (
            .O(N__30580),
            .I(N__30575));
    GlobalMux I__5578 (
            .O(N__30575),
            .I(N__30572));
    gio2CtrlBuf I__5577 (
            .O(N__30572),
            .I(delay_hc_input_c_g));
    CascadeMux I__5576 (
            .O(N__30569),
            .I(N__30565));
    InMux I__5575 (
            .O(N__30568),
            .I(N__30562));
    InMux I__5574 (
            .O(N__30565),
            .I(N__30559));
    LocalMux I__5573 (
            .O(N__30562),
            .I(N__30554));
    LocalMux I__5572 (
            .O(N__30559),
            .I(N__30551));
    InMux I__5571 (
            .O(N__30558),
            .I(N__30548));
    InMux I__5570 (
            .O(N__30557),
            .I(N__30545));
    Span4Mux_h I__5569 (
            .O(N__30554),
            .I(N__30542));
    Span4Mux_v I__5568 (
            .O(N__30551),
            .I(N__30539));
    LocalMux I__5567 (
            .O(N__30548),
            .I(N__30534));
    LocalMux I__5566 (
            .O(N__30545),
            .I(N__30534));
    Odrv4 I__5565 (
            .O(N__30542),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__5564 (
            .O(N__30539),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv12 I__5563 (
            .O(N__30534),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    InMux I__5562 (
            .O(N__30527),
            .I(N__30524));
    LocalMux I__5561 (
            .O(N__30524),
            .I(N__30521));
    Odrv12 I__5560 (
            .O(N__30521),
            .I(\current_shift_inst.PI_CTRL.integrator_i_1 ));
    CascadeMux I__5559 (
            .O(N__30518),
            .I(N__30515));
    InMux I__5558 (
            .O(N__30515),
            .I(N__30511));
    InMux I__5557 (
            .O(N__30514),
            .I(N__30508));
    LocalMux I__5556 (
            .O(N__30511),
            .I(N__30503));
    LocalMux I__5555 (
            .O(N__30508),
            .I(N__30503));
    Odrv12 I__5554 (
            .O(N__30503),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_i_12 ));
    CascadeMux I__5553 (
            .O(N__30500),
            .I(N__30496));
    InMux I__5552 (
            .O(N__30499),
            .I(N__30492));
    InMux I__5551 (
            .O(N__30496),
            .I(N__30489));
    InMux I__5550 (
            .O(N__30495),
            .I(N__30486));
    LocalMux I__5549 (
            .O(N__30492),
            .I(N__30483));
    LocalMux I__5548 (
            .O(N__30489),
            .I(N__30480));
    LocalMux I__5547 (
            .O(N__30486),
            .I(N__30477));
    Span4Mux_h I__5546 (
            .O(N__30483),
            .I(N__30472));
    Span4Mux_v I__5545 (
            .O(N__30480),
            .I(N__30469));
    Span4Mux_v I__5544 (
            .O(N__30477),
            .I(N__30466));
    InMux I__5543 (
            .O(N__30476),
            .I(N__30463));
    InMux I__5542 (
            .O(N__30475),
            .I(N__30460));
    Odrv4 I__5541 (
            .O(N__30472),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__5540 (
            .O(N__30469),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__5539 (
            .O(N__30466),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    LocalMux I__5538 (
            .O(N__30463),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    LocalMux I__5537 (
            .O(N__30460),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    InMux I__5536 (
            .O(N__30449),
            .I(N__30446));
    LocalMux I__5535 (
            .O(N__30446),
            .I(N__30443));
    Span4Mux_h I__5534 (
            .O(N__30443),
            .I(N__30440));
    Odrv4 I__5533 (
            .O(N__30440),
            .I(\current_shift_inst.PI_CTRL.integrator_i_24 ));
    CascadeMux I__5532 (
            .O(N__30437),
            .I(N__30433));
    CascadeMux I__5531 (
            .O(N__30436),
            .I(N__30430));
    InMux I__5530 (
            .O(N__30433),
            .I(N__30424));
    InMux I__5529 (
            .O(N__30430),
            .I(N__30424));
    InMux I__5528 (
            .O(N__30429),
            .I(N__30421));
    LocalMux I__5527 (
            .O(N__30424),
            .I(N__30418));
    LocalMux I__5526 (
            .O(N__30421),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    Odrv12 I__5525 (
            .O(N__30418),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__5524 (
            .O(N__30413),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    CascadeMux I__5523 (
            .O(N__30410),
            .I(N__30406));
    CascadeMux I__5522 (
            .O(N__30409),
            .I(N__30403));
    InMux I__5521 (
            .O(N__30406),
            .I(N__30397));
    InMux I__5520 (
            .O(N__30403),
            .I(N__30397));
    InMux I__5519 (
            .O(N__30402),
            .I(N__30394));
    LocalMux I__5518 (
            .O(N__30397),
            .I(N__30391));
    LocalMux I__5517 (
            .O(N__30394),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    Odrv12 I__5516 (
            .O(N__30391),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__5515 (
            .O(N__30386),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    CascadeMux I__5514 (
            .O(N__30383),
            .I(N__30380));
    InMux I__5513 (
            .O(N__30380),
            .I(N__30375));
    InMux I__5512 (
            .O(N__30379),
            .I(N__30372));
    InMux I__5511 (
            .O(N__30378),
            .I(N__30369));
    LocalMux I__5510 (
            .O(N__30375),
            .I(N__30364));
    LocalMux I__5509 (
            .O(N__30372),
            .I(N__30364));
    LocalMux I__5508 (
            .O(N__30369),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv12 I__5507 (
            .O(N__30364),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__5506 (
            .O(N__30359),
            .I(bfn_11_22_0_));
    InMux I__5505 (
            .O(N__30356),
            .I(N__30352));
    InMux I__5504 (
            .O(N__30355),
            .I(N__30349));
    LocalMux I__5503 (
            .O(N__30352),
            .I(N__30343));
    LocalMux I__5502 (
            .O(N__30349),
            .I(N__30343));
    InMux I__5501 (
            .O(N__30348),
            .I(N__30340));
    Span4Mux_v I__5500 (
            .O(N__30343),
            .I(N__30337));
    LocalMux I__5499 (
            .O(N__30340),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__5498 (
            .O(N__30337),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__5497 (
            .O(N__30332),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    CascadeMux I__5496 (
            .O(N__30329),
            .I(N__30326));
    InMux I__5495 (
            .O(N__30326),
            .I(N__30322));
    InMux I__5494 (
            .O(N__30325),
            .I(N__30319));
    LocalMux I__5493 (
            .O(N__30322),
            .I(N__30313));
    LocalMux I__5492 (
            .O(N__30319),
            .I(N__30313));
    InMux I__5491 (
            .O(N__30318),
            .I(N__30310));
    Span4Mux_h I__5490 (
            .O(N__30313),
            .I(N__30307));
    LocalMux I__5489 (
            .O(N__30310),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    Odrv4 I__5488 (
            .O(N__30307),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    InMux I__5487 (
            .O(N__30302),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    CascadeMux I__5486 (
            .O(N__30299),
            .I(N__30295));
    CascadeMux I__5485 (
            .O(N__30298),
            .I(N__30292));
    InMux I__5484 (
            .O(N__30295),
            .I(N__30286));
    InMux I__5483 (
            .O(N__30292),
            .I(N__30286));
    InMux I__5482 (
            .O(N__30291),
            .I(N__30283));
    LocalMux I__5481 (
            .O(N__30286),
            .I(N__30280));
    LocalMux I__5480 (
            .O(N__30283),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    Odrv12 I__5479 (
            .O(N__30280),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__5478 (
            .O(N__30275),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    InMux I__5477 (
            .O(N__30272),
            .I(N__30268));
    InMux I__5476 (
            .O(N__30271),
            .I(N__30265));
    LocalMux I__5475 (
            .O(N__30268),
            .I(N__30262));
    LocalMux I__5474 (
            .O(N__30265),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    Odrv12 I__5473 (
            .O(N__30262),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    InMux I__5472 (
            .O(N__30257),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__5471 (
            .O(N__30254),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    InMux I__5470 (
            .O(N__30251),
            .I(N__30247));
    InMux I__5469 (
            .O(N__30250),
            .I(N__30244));
    LocalMux I__5468 (
            .O(N__30247),
            .I(N__30241));
    LocalMux I__5467 (
            .O(N__30244),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    Odrv12 I__5466 (
            .O(N__30241),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    InMux I__5465 (
            .O(N__30236),
            .I(N__30204));
    InMux I__5464 (
            .O(N__30235),
            .I(N__30204));
    InMux I__5463 (
            .O(N__30234),
            .I(N__30204));
    InMux I__5462 (
            .O(N__30233),
            .I(N__30204));
    InMux I__5461 (
            .O(N__30232),
            .I(N__30195));
    InMux I__5460 (
            .O(N__30231),
            .I(N__30195));
    InMux I__5459 (
            .O(N__30230),
            .I(N__30195));
    InMux I__5458 (
            .O(N__30229),
            .I(N__30195));
    InMux I__5457 (
            .O(N__30228),
            .I(N__30180));
    InMux I__5456 (
            .O(N__30227),
            .I(N__30180));
    InMux I__5455 (
            .O(N__30226),
            .I(N__30180));
    InMux I__5454 (
            .O(N__30225),
            .I(N__30180));
    InMux I__5453 (
            .O(N__30224),
            .I(N__30171));
    InMux I__5452 (
            .O(N__30223),
            .I(N__30171));
    InMux I__5451 (
            .O(N__30222),
            .I(N__30171));
    InMux I__5450 (
            .O(N__30221),
            .I(N__30171));
    InMux I__5449 (
            .O(N__30220),
            .I(N__30162));
    InMux I__5448 (
            .O(N__30219),
            .I(N__30162));
    InMux I__5447 (
            .O(N__30218),
            .I(N__30162));
    InMux I__5446 (
            .O(N__30217),
            .I(N__30162));
    InMux I__5445 (
            .O(N__30216),
            .I(N__30153));
    InMux I__5444 (
            .O(N__30215),
            .I(N__30153));
    InMux I__5443 (
            .O(N__30214),
            .I(N__30153));
    InMux I__5442 (
            .O(N__30213),
            .I(N__30153));
    LocalMux I__5441 (
            .O(N__30204),
            .I(N__30150));
    LocalMux I__5440 (
            .O(N__30195),
            .I(N__30147));
    InMux I__5439 (
            .O(N__30194),
            .I(N__30142));
    InMux I__5438 (
            .O(N__30193),
            .I(N__30142));
    InMux I__5437 (
            .O(N__30192),
            .I(N__30133));
    InMux I__5436 (
            .O(N__30191),
            .I(N__30133));
    InMux I__5435 (
            .O(N__30190),
            .I(N__30133));
    InMux I__5434 (
            .O(N__30189),
            .I(N__30133));
    LocalMux I__5433 (
            .O(N__30180),
            .I(N__30130));
    LocalMux I__5432 (
            .O(N__30171),
            .I(N__30119));
    LocalMux I__5431 (
            .O(N__30162),
            .I(N__30119));
    LocalMux I__5430 (
            .O(N__30153),
            .I(N__30119));
    Span4Mux_h I__5429 (
            .O(N__30150),
            .I(N__30119));
    Span4Mux_h I__5428 (
            .O(N__30147),
            .I(N__30119));
    LocalMux I__5427 (
            .O(N__30142),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    LocalMux I__5426 (
            .O(N__30133),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__5425 (
            .O(N__30130),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__5424 (
            .O(N__30119),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    CascadeMux I__5423 (
            .O(N__30110),
            .I(N__30107));
    InMux I__5422 (
            .O(N__30107),
            .I(N__30103));
    InMux I__5421 (
            .O(N__30106),
            .I(N__30100));
    LocalMux I__5420 (
            .O(N__30103),
            .I(N__30094));
    LocalMux I__5419 (
            .O(N__30100),
            .I(N__30094));
    InMux I__5418 (
            .O(N__30099),
            .I(N__30091));
    Span4Mux_v I__5417 (
            .O(N__30094),
            .I(N__30088));
    LocalMux I__5416 (
            .O(N__30091),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    Odrv4 I__5415 (
            .O(N__30088),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__5414 (
            .O(N__30083),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    InMux I__5413 (
            .O(N__30080),
            .I(N__30074));
    InMux I__5412 (
            .O(N__30079),
            .I(N__30074));
    LocalMux I__5411 (
            .O(N__30074),
            .I(N__30070));
    InMux I__5410 (
            .O(N__30073),
            .I(N__30067));
    Span4Mux_v I__5409 (
            .O(N__30070),
            .I(N__30064));
    LocalMux I__5408 (
            .O(N__30067),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    Odrv4 I__5407 (
            .O(N__30064),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__5406 (
            .O(N__30059),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    CascadeMux I__5405 (
            .O(N__30056),
            .I(N__30053));
    InMux I__5404 (
            .O(N__30053),
            .I(N__30049));
    InMux I__5403 (
            .O(N__30052),
            .I(N__30046));
    LocalMux I__5402 (
            .O(N__30049),
            .I(N__30042));
    LocalMux I__5401 (
            .O(N__30046),
            .I(N__30039));
    InMux I__5400 (
            .O(N__30045),
            .I(N__30036));
    Span4Mux_v I__5399 (
            .O(N__30042),
            .I(N__30031));
    Span4Mux_v I__5398 (
            .O(N__30039),
            .I(N__30031));
    LocalMux I__5397 (
            .O(N__30036),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__5396 (
            .O(N__30031),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__5395 (
            .O(N__30026),
            .I(bfn_11_21_0_));
    CascadeMux I__5394 (
            .O(N__30023),
            .I(N__30019));
    CascadeMux I__5393 (
            .O(N__30022),
            .I(N__30016));
    InMux I__5392 (
            .O(N__30019),
            .I(N__30013));
    InMux I__5391 (
            .O(N__30016),
            .I(N__30010));
    LocalMux I__5390 (
            .O(N__30013),
            .I(N__30004));
    LocalMux I__5389 (
            .O(N__30010),
            .I(N__30004));
    InMux I__5388 (
            .O(N__30009),
            .I(N__30001));
    Span4Mux_v I__5387 (
            .O(N__30004),
            .I(N__29998));
    LocalMux I__5386 (
            .O(N__30001),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__5385 (
            .O(N__29998),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__5384 (
            .O(N__29993),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    CascadeMux I__5383 (
            .O(N__29990),
            .I(N__29987));
    InMux I__5382 (
            .O(N__29987),
            .I(N__29983));
    InMux I__5381 (
            .O(N__29986),
            .I(N__29980));
    LocalMux I__5380 (
            .O(N__29983),
            .I(N__29974));
    LocalMux I__5379 (
            .O(N__29980),
            .I(N__29974));
    InMux I__5378 (
            .O(N__29979),
            .I(N__29971));
    Span4Mux_h I__5377 (
            .O(N__29974),
            .I(N__29968));
    LocalMux I__5376 (
            .O(N__29971),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    Odrv4 I__5375 (
            .O(N__29968),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__5374 (
            .O(N__29963),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    InMux I__5373 (
            .O(N__29960),
            .I(N__29953));
    InMux I__5372 (
            .O(N__29959),
            .I(N__29953));
    InMux I__5371 (
            .O(N__29958),
            .I(N__29950));
    LocalMux I__5370 (
            .O(N__29953),
            .I(N__29947));
    LocalMux I__5369 (
            .O(N__29950),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    Odrv12 I__5368 (
            .O(N__29947),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__5367 (
            .O(N__29942),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    InMux I__5366 (
            .O(N__29939),
            .I(N__29932));
    InMux I__5365 (
            .O(N__29938),
            .I(N__29932));
    InMux I__5364 (
            .O(N__29937),
            .I(N__29929));
    LocalMux I__5363 (
            .O(N__29932),
            .I(N__29926));
    LocalMux I__5362 (
            .O(N__29929),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    Odrv12 I__5361 (
            .O(N__29926),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__5360 (
            .O(N__29921),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    CascadeMux I__5359 (
            .O(N__29918),
            .I(N__29914));
    InMux I__5358 (
            .O(N__29917),
            .I(N__29910));
    InMux I__5357 (
            .O(N__29914),
            .I(N__29907));
    InMux I__5356 (
            .O(N__29913),
            .I(N__29904));
    LocalMux I__5355 (
            .O(N__29910),
            .I(N__29899));
    LocalMux I__5354 (
            .O(N__29907),
            .I(N__29899));
    LocalMux I__5353 (
            .O(N__29904),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    Odrv12 I__5352 (
            .O(N__29899),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__5351 (
            .O(N__29894),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    InMux I__5350 (
            .O(N__29891),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    CascadeMux I__5349 (
            .O(N__29888),
            .I(N__29885));
    InMux I__5348 (
            .O(N__29885),
            .I(N__29881));
    InMux I__5347 (
            .O(N__29884),
            .I(N__29878));
    LocalMux I__5346 (
            .O(N__29881),
            .I(N__29872));
    LocalMux I__5345 (
            .O(N__29878),
            .I(N__29872));
    InMux I__5344 (
            .O(N__29877),
            .I(N__29869));
    Span4Mux_v I__5343 (
            .O(N__29872),
            .I(N__29866));
    LocalMux I__5342 (
            .O(N__29869),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    Odrv4 I__5341 (
            .O(N__29866),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__5340 (
            .O(N__29861),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    InMux I__5339 (
            .O(N__29858),
            .I(N__29852));
    InMux I__5338 (
            .O(N__29857),
            .I(N__29852));
    LocalMux I__5337 (
            .O(N__29852),
            .I(N__29848));
    InMux I__5336 (
            .O(N__29851),
            .I(N__29845));
    Span4Mux_v I__5335 (
            .O(N__29848),
            .I(N__29842));
    LocalMux I__5334 (
            .O(N__29845),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    Odrv4 I__5333 (
            .O(N__29842),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__5332 (
            .O(N__29837),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    CascadeMux I__5331 (
            .O(N__29834),
            .I(N__29831));
    InMux I__5330 (
            .O(N__29831),
            .I(N__29828));
    LocalMux I__5329 (
            .O(N__29828),
            .I(N__29823));
    InMux I__5328 (
            .O(N__29827),
            .I(N__29820));
    InMux I__5327 (
            .O(N__29826),
            .I(N__29817));
    Span4Mux_v I__5326 (
            .O(N__29823),
            .I(N__29814));
    LocalMux I__5325 (
            .O(N__29820),
            .I(N__29811));
    LocalMux I__5324 (
            .O(N__29817),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv4 I__5323 (
            .O(N__29814),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv12 I__5322 (
            .O(N__29811),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__5321 (
            .O(N__29804),
            .I(bfn_11_20_0_));
    InMux I__5320 (
            .O(N__29801),
            .I(N__29797));
    CascadeMux I__5319 (
            .O(N__29800),
            .I(N__29794));
    LocalMux I__5318 (
            .O(N__29797),
            .I(N__29790));
    InMux I__5317 (
            .O(N__29794),
            .I(N__29787));
    InMux I__5316 (
            .O(N__29793),
            .I(N__29784));
    Span4Mux_h I__5315 (
            .O(N__29790),
            .I(N__29781));
    LocalMux I__5314 (
            .O(N__29787),
            .I(N__29778));
    LocalMux I__5313 (
            .O(N__29784),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv4 I__5312 (
            .O(N__29781),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv12 I__5311 (
            .O(N__29778),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__5310 (
            .O(N__29771),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    InMux I__5309 (
            .O(N__29768),
            .I(N__29762));
    InMux I__5308 (
            .O(N__29767),
            .I(N__29762));
    LocalMux I__5307 (
            .O(N__29762),
            .I(N__29758));
    InMux I__5306 (
            .O(N__29761),
            .I(N__29755));
    Span4Mux_v I__5305 (
            .O(N__29758),
            .I(N__29752));
    LocalMux I__5304 (
            .O(N__29755),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    Odrv4 I__5303 (
            .O(N__29752),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__5302 (
            .O(N__29747),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    CascadeMux I__5301 (
            .O(N__29744),
            .I(N__29740));
    CascadeMux I__5300 (
            .O(N__29743),
            .I(N__29737));
    InMux I__5299 (
            .O(N__29740),
            .I(N__29731));
    InMux I__5298 (
            .O(N__29737),
            .I(N__29731));
    InMux I__5297 (
            .O(N__29736),
            .I(N__29728));
    LocalMux I__5296 (
            .O(N__29731),
            .I(N__29725));
    LocalMux I__5295 (
            .O(N__29728),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    Odrv12 I__5294 (
            .O(N__29725),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__5293 (
            .O(N__29720),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    CascadeMux I__5292 (
            .O(N__29717),
            .I(N__29713));
    CascadeMux I__5291 (
            .O(N__29716),
            .I(N__29710));
    InMux I__5290 (
            .O(N__29713),
            .I(N__29704));
    InMux I__5289 (
            .O(N__29710),
            .I(N__29704));
    InMux I__5288 (
            .O(N__29709),
            .I(N__29701));
    LocalMux I__5287 (
            .O(N__29704),
            .I(N__29698));
    LocalMux I__5286 (
            .O(N__29701),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    Odrv12 I__5285 (
            .O(N__29698),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__5284 (
            .O(N__29693),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    CascadeMux I__5283 (
            .O(N__29690),
            .I(N__29687));
    InMux I__5282 (
            .O(N__29687),
            .I(N__29683));
    InMux I__5281 (
            .O(N__29686),
            .I(N__29680));
    LocalMux I__5280 (
            .O(N__29683),
            .I(N__29674));
    LocalMux I__5279 (
            .O(N__29680),
            .I(N__29674));
    InMux I__5278 (
            .O(N__29679),
            .I(N__29671));
    Span4Mux_v I__5277 (
            .O(N__29674),
            .I(N__29668));
    LocalMux I__5276 (
            .O(N__29671),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    Odrv4 I__5275 (
            .O(N__29668),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__5274 (
            .O(N__29663),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    InMux I__5273 (
            .O(N__29660),
            .I(N__29657));
    LocalMux I__5272 (
            .O(N__29657),
            .I(N__29654));
    Span4Mux_h I__5271 (
            .O(N__29654),
            .I(N__29650));
    InMux I__5270 (
            .O(N__29653),
            .I(N__29647));
    Odrv4 I__5269 (
            .O(N__29650),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    LocalMux I__5268 (
            .O(N__29647),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    InMux I__5267 (
            .O(N__29642),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__5266 (
            .O(N__29639),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__5265 (
            .O(N__29636),
            .I(N__29632));
    InMux I__5264 (
            .O(N__29635),
            .I(N__29628));
    LocalMux I__5263 (
            .O(N__29632),
            .I(N__29625));
    InMux I__5262 (
            .O(N__29631),
            .I(N__29622));
    LocalMux I__5261 (
            .O(N__29628),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    Odrv12 I__5260 (
            .O(N__29625),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__5259 (
            .O(N__29622),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    InMux I__5258 (
            .O(N__29615),
            .I(bfn_11_19_0_));
    InMux I__5257 (
            .O(N__29612),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    InMux I__5256 (
            .O(N__29609),
            .I(N__29605));
    CascadeMux I__5255 (
            .O(N__29608),
            .I(N__29602));
    LocalMux I__5254 (
            .O(N__29605),
            .I(N__29598));
    InMux I__5253 (
            .O(N__29602),
            .I(N__29595));
    InMux I__5252 (
            .O(N__29601),
            .I(N__29592));
    Span4Mux_h I__5251 (
            .O(N__29598),
            .I(N__29589));
    LocalMux I__5250 (
            .O(N__29595),
            .I(N__29586));
    LocalMux I__5249 (
            .O(N__29592),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    Odrv4 I__5248 (
            .O(N__29589),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    Odrv12 I__5247 (
            .O(N__29586),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__5246 (
            .O(N__29579),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    CascadeMux I__5245 (
            .O(N__29576),
            .I(N__29572));
    InMux I__5244 (
            .O(N__29575),
            .I(N__29569));
    InMux I__5243 (
            .O(N__29572),
            .I(N__29566));
    LocalMux I__5242 (
            .O(N__29569),
            .I(N__29560));
    LocalMux I__5241 (
            .O(N__29566),
            .I(N__29560));
    InMux I__5240 (
            .O(N__29565),
            .I(N__29557));
    Span4Mux_h I__5239 (
            .O(N__29560),
            .I(N__29554));
    LocalMux I__5238 (
            .O(N__29557),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    Odrv4 I__5237 (
            .O(N__29554),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__5236 (
            .O(N__29549),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    CascadeMux I__5235 (
            .O(N__29546),
            .I(N__29542));
    CascadeMux I__5234 (
            .O(N__29545),
            .I(N__29539));
    InMux I__5233 (
            .O(N__29542),
            .I(N__29533));
    InMux I__5232 (
            .O(N__29539),
            .I(N__29533));
    InMux I__5231 (
            .O(N__29538),
            .I(N__29530));
    LocalMux I__5230 (
            .O(N__29533),
            .I(N__29527));
    LocalMux I__5229 (
            .O(N__29530),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    Odrv12 I__5228 (
            .O(N__29527),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__5227 (
            .O(N__29522),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    CascadeMux I__5226 (
            .O(N__29519),
            .I(N__29515));
    CascadeMux I__5225 (
            .O(N__29518),
            .I(N__29512));
    InMux I__5224 (
            .O(N__29515),
            .I(N__29507));
    InMux I__5223 (
            .O(N__29512),
            .I(N__29507));
    LocalMux I__5222 (
            .O(N__29507),
            .I(N__29503));
    InMux I__5221 (
            .O(N__29506),
            .I(N__29500));
    Span4Mux_h I__5220 (
            .O(N__29503),
            .I(N__29497));
    LocalMux I__5219 (
            .O(N__29500),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    Odrv4 I__5218 (
            .O(N__29497),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__5217 (
            .O(N__29492),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__5216 (
            .O(N__29489),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__5215 (
            .O(N__29486),
            .I(N__29483));
    LocalMux I__5214 (
            .O(N__29483),
            .I(N__29479));
    InMux I__5213 (
            .O(N__29482),
            .I(N__29476));
    Odrv4 I__5212 (
            .O(N__29479),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    LocalMux I__5211 (
            .O(N__29476),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__5210 (
            .O(N__29471),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__5209 (
            .O(N__29468),
            .I(N__29465));
    LocalMux I__5208 (
            .O(N__29465),
            .I(N__29461));
    InMux I__5207 (
            .O(N__29464),
            .I(N__29458));
    Odrv4 I__5206 (
            .O(N__29461),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    LocalMux I__5205 (
            .O(N__29458),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    InMux I__5204 (
            .O(N__29453),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__5203 (
            .O(N__29450),
            .I(N__29447));
    LocalMux I__5202 (
            .O(N__29447),
            .I(N__29443));
    CascadeMux I__5201 (
            .O(N__29446),
            .I(N__29440));
    Span4Mux_h I__5200 (
            .O(N__29443),
            .I(N__29437));
    InMux I__5199 (
            .O(N__29440),
            .I(N__29434));
    Odrv4 I__5198 (
            .O(N__29437),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    LocalMux I__5197 (
            .O(N__29434),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    InMux I__5196 (
            .O(N__29429),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__5195 (
            .O(N__29426),
            .I(N__29423));
    InMux I__5194 (
            .O(N__29423),
            .I(N__29420));
    LocalMux I__5193 (
            .O(N__29420),
            .I(N__29417));
    Span4Mux_v I__5192 (
            .O(N__29417),
            .I(N__29413));
    InMux I__5191 (
            .O(N__29416),
            .I(N__29410));
    Odrv4 I__5190 (
            .O(N__29413),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    LocalMux I__5189 (
            .O(N__29410),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    InMux I__5188 (
            .O(N__29405),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__5187 (
            .O(N__29402),
            .I(N__29399));
    InMux I__5186 (
            .O(N__29399),
            .I(N__29396));
    LocalMux I__5185 (
            .O(N__29396),
            .I(N__29393));
    Span4Mux_v I__5184 (
            .O(N__29393),
            .I(N__29390));
    Span4Mux_v I__5183 (
            .O(N__29390),
            .I(N__29386));
    InMux I__5182 (
            .O(N__29389),
            .I(N__29383));
    Odrv4 I__5181 (
            .O(N__29386),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    LocalMux I__5180 (
            .O(N__29383),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    InMux I__5179 (
            .O(N__29378),
            .I(bfn_11_18_0_));
    CascadeMux I__5178 (
            .O(N__29375),
            .I(N__29372));
    InMux I__5177 (
            .O(N__29372),
            .I(N__29369));
    LocalMux I__5176 (
            .O(N__29369),
            .I(N__29365));
    CascadeMux I__5175 (
            .O(N__29368),
            .I(N__29362));
    Span4Mux_v I__5174 (
            .O(N__29365),
            .I(N__29359));
    InMux I__5173 (
            .O(N__29362),
            .I(N__29356));
    Odrv4 I__5172 (
            .O(N__29359),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    LocalMux I__5171 (
            .O(N__29356),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    InMux I__5170 (
            .O(N__29351),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    CascadeMux I__5169 (
            .O(N__29348),
            .I(N__29345));
    InMux I__5168 (
            .O(N__29345),
            .I(N__29342));
    LocalMux I__5167 (
            .O(N__29342),
            .I(N__29339));
    Span4Mux_v I__5166 (
            .O(N__29339),
            .I(N__29335));
    InMux I__5165 (
            .O(N__29338),
            .I(N__29332));
    Odrv4 I__5164 (
            .O(N__29335),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    LocalMux I__5163 (
            .O(N__29332),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    InMux I__5162 (
            .O(N__29327),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__5161 (
            .O(N__29324),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__5160 (
            .O(N__29321),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__5159 (
            .O(N__29318),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__5158 (
            .O(N__29315),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__5157 (
            .O(N__29312),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__5156 (
            .O(N__29309),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__5155 (
            .O(N__29306),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__5154 (
            .O(N__29303),
            .I(bfn_11_17_0_));
    InMux I__5153 (
            .O(N__29300),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__5152 (
            .O(N__29297),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__5151 (
            .O(N__29294),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__5150 (
            .O(N__29291),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__5149 (
            .O(N__29288),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__5148 (
            .O(N__29285),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__5147 (
            .O(N__29282),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__5146 (
            .O(N__29279),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__5145 (
            .O(N__29276),
            .I(bfn_11_16_0_));
    InMux I__5144 (
            .O(N__29273),
            .I(N__29268));
    InMux I__5143 (
            .O(N__29272),
            .I(N__29265));
    CascadeMux I__5142 (
            .O(N__29271),
            .I(N__29260));
    LocalMux I__5141 (
            .O(N__29268),
            .I(N__29257));
    LocalMux I__5140 (
            .O(N__29265),
            .I(N__29254));
    InMux I__5139 (
            .O(N__29264),
            .I(N__29247));
    InMux I__5138 (
            .O(N__29263),
            .I(N__29247));
    InMux I__5137 (
            .O(N__29260),
            .I(N__29247));
    Span4Mux_h I__5136 (
            .O(N__29257),
            .I(N__29244));
    Span4Mux_h I__5135 (
            .O(N__29254),
            .I(N__29239));
    LocalMux I__5134 (
            .O(N__29247),
            .I(N__29239));
    Odrv4 I__5133 (
            .O(N__29244),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__5132 (
            .O(N__29239),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    InMux I__5131 (
            .O(N__29234),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_31 ));
    CascadeMux I__5130 (
            .O(N__29231),
            .I(N__29228));
    InMux I__5129 (
            .O(N__29228),
            .I(N__29225));
    LocalMux I__5128 (
            .O(N__29225),
            .I(N__29222));
    Span4Mux_h I__5127 (
            .O(N__29222),
            .I(N__29219));
    Odrv4 I__5126 (
            .O(N__29219),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0 ));
    CascadeMux I__5125 (
            .O(N__29216),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i_cascade_ ));
    InMux I__5124 (
            .O(N__29213),
            .I(N__29209));
    InMux I__5123 (
            .O(N__29212),
            .I(N__29206));
    LocalMux I__5122 (
            .O(N__29209),
            .I(elapsed_time_ns_1_RNIP3OD11_0_30));
    LocalMux I__5121 (
            .O(N__29206),
            .I(elapsed_time_ns_1_RNIP3OD11_0_30));
    CascadeMux I__5120 (
            .O(N__29201),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91Z0Z_7_cascade_ ));
    CascadeMux I__5119 (
            .O(N__29198),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2Z0Z_15_cascade_ ));
    InMux I__5118 (
            .O(N__29195),
            .I(N__29192));
    LocalMux I__5117 (
            .O(N__29192),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719Z0Z_21 ));
    CascadeMux I__5116 (
            .O(N__29189),
            .I(N__29185));
    InMux I__5115 (
            .O(N__29188),
            .I(N__29177));
    InMux I__5114 (
            .O(N__29185),
            .I(N__29177));
    InMux I__5113 (
            .O(N__29184),
            .I(N__29177));
    LocalMux I__5112 (
            .O(N__29177),
            .I(N__29174));
    Odrv4 I__5111 (
            .O(N__29174),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992Z0Z_24 ));
    InMux I__5110 (
            .O(N__29171),
            .I(N__29168));
    LocalMux I__5109 (
            .O(N__29168),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9Z0Z_24 ));
    InMux I__5108 (
            .O(N__29165),
            .I(N__29161));
    InMux I__5107 (
            .O(N__29164),
            .I(N__29158));
    LocalMux I__5106 (
            .O(N__29161),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ));
    LocalMux I__5105 (
            .O(N__29158),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ));
    InMux I__5104 (
            .O(N__29153),
            .I(N__29150));
    LocalMux I__5103 (
            .O(N__29150),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO ));
    InMux I__5102 (
            .O(N__29147),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ));
    InMux I__5101 (
            .O(N__29144),
            .I(N__29141));
    LocalMux I__5100 (
            .O(N__29141),
            .I(N__29138));
    Odrv4 I__5099 (
            .O(N__29138),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO ));
    InMux I__5098 (
            .O(N__29135),
            .I(bfn_11_13_0_));
    InMux I__5097 (
            .O(N__29132),
            .I(N__29129));
    LocalMux I__5096 (
            .O(N__29129),
            .I(N__29126));
    Odrv4 I__5095 (
            .O(N__29126),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO ));
    InMux I__5094 (
            .O(N__29123),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ));
    CascadeMux I__5093 (
            .O(N__29120),
            .I(N__29117));
    InMux I__5092 (
            .O(N__29117),
            .I(N__29114));
    LocalMux I__5091 (
            .O(N__29114),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ));
    InMux I__5090 (
            .O(N__29111),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ));
    InMux I__5089 (
            .O(N__29108),
            .I(N__29103));
    InMux I__5088 (
            .O(N__29107),
            .I(N__29100));
    InMux I__5087 (
            .O(N__29106),
            .I(N__29097));
    LocalMux I__5086 (
            .O(N__29103),
            .I(N__29092));
    LocalMux I__5085 (
            .O(N__29100),
            .I(N__29092));
    LocalMux I__5084 (
            .O(N__29097),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ));
    Odrv4 I__5083 (
            .O(N__29092),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ));
    CascadeMux I__5082 (
            .O(N__29087),
            .I(N__29084));
    InMux I__5081 (
            .O(N__29084),
            .I(N__29081));
    LocalMux I__5080 (
            .O(N__29081),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ));
    InMux I__5079 (
            .O(N__29078),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ));
    InMux I__5078 (
            .O(N__29075),
            .I(N__29072));
    LocalMux I__5077 (
            .O(N__29072),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ));
    InMux I__5076 (
            .O(N__29069),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ));
    InMux I__5075 (
            .O(N__29066),
            .I(N__29063));
    LocalMux I__5074 (
            .O(N__29063),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ));
    InMux I__5073 (
            .O(N__29060),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ));
    InMux I__5072 (
            .O(N__29057),
            .I(N__29053));
    InMux I__5071 (
            .O(N__29056),
            .I(N__29050));
    LocalMux I__5070 (
            .O(N__29053),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ));
    LocalMux I__5069 (
            .O(N__29050),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ));
    InMux I__5068 (
            .O(N__29045),
            .I(N__29042));
    LocalMux I__5067 (
            .O(N__29042),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ));
    InMux I__5066 (
            .O(N__29039),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ));
    InMux I__5065 (
            .O(N__29036),
            .I(N__29032));
    InMux I__5064 (
            .O(N__29035),
            .I(N__29029));
    LocalMux I__5063 (
            .O(N__29032),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ));
    LocalMux I__5062 (
            .O(N__29029),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ));
    InMux I__5061 (
            .O(N__29024),
            .I(N__29021));
    LocalMux I__5060 (
            .O(N__29021),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO ));
    InMux I__5059 (
            .O(N__29018),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ));
    InMux I__5058 (
            .O(N__29015),
            .I(N__29010));
    InMux I__5057 (
            .O(N__29014),
            .I(N__29007));
    InMux I__5056 (
            .O(N__29013),
            .I(N__29004));
    LocalMux I__5055 (
            .O(N__29010),
            .I(N__29001));
    LocalMux I__5054 (
            .O(N__29007),
            .I(N__28998));
    LocalMux I__5053 (
            .O(N__29004),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ));
    Odrv4 I__5052 (
            .O(N__29001),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ));
    Odrv12 I__5051 (
            .O(N__28998),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ));
    InMux I__5050 (
            .O(N__28991),
            .I(N__28988));
    LocalMux I__5049 (
            .O(N__28988),
            .I(N__28985));
    Odrv4 I__5048 (
            .O(N__28985),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO ));
    InMux I__5047 (
            .O(N__28982),
            .I(bfn_11_12_0_));
    InMux I__5046 (
            .O(N__28979),
            .I(N__28976));
    LocalMux I__5045 (
            .O(N__28976),
            .I(N__28971));
    InMux I__5044 (
            .O(N__28975),
            .I(N__28968));
    InMux I__5043 (
            .O(N__28974),
            .I(N__28965));
    Span4Mux_h I__5042 (
            .O(N__28971),
            .I(N__28962));
    LocalMux I__5041 (
            .O(N__28968),
            .I(N__28959));
    LocalMux I__5040 (
            .O(N__28965),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ));
    Odrv4 I__5039 (
            .O(N__28962),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ));
    Odrv12 I__5038 (
            .O(N__28959),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ));
    CascadeMux I__5037 (
            .O(N__28952),
            .I(N__28949));
    InMux I__5036 (
            .O(N__28949),
            .I(N__28946));
    LocalMux I__5035 (
            .O(N__28946),
            .I(N__28943));
    Odrv4 I__5034 (
            .O(N__28943),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO ));
    InMux I__5033 (
            .O(N__28940),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ));
    InMux I__5032 (
            .O(N__28937),
            .I(N__28934));
    LocalMux I__5031 (
            .O(N__28934),
            .I(N__28930));
    InMux I__5030 (
            .O(N__28933),
            .I(N__28926));
    Sp12to4 I__5029 (
            .O(N__28930),
            .I(N__28923));
    InMux I__5028 (
            .O(N__28929),
            .I(N__28920));
    LocalMux I__5027 (
            .O(N__28926),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ));
    Odrv12 I__5026 (
            .O(N__28923),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ));
    LocalMux I__5025 (
            .O(N__28920),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ));
    CascadeMux I__5024 (
            .O(N__28913),
            .I(N__28910));
    InMux I__5023 (
            .O(N__28910),
            .I(N__28907));
    LocalMux I__5022 (
            .O(N__28907),
            .I(N__28904));
    Odrv4 I__5021 (
            .O(N__28904),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO ));
    InMux I__5020 (
            .O(N__28901),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ));
    InMux I__5019 (
            .O(N__28898),
            .I(N__28893));
    CascadeMux I__5018 (
            .O(N__28897),
            .I(N__28890));
    InMux I__5017 (
            .O(N__28896),
            .I(N__28887));
    LocalMux I__5016 (
            .O(N__28893),
            .I(N__28884));
    InMux I__5015 (
            .O(N__28890),
            .I(N__28881));
    LocalMux I__5014 (
            .O(N__28887),
            .I(N__28876));
    Span4Mux_v I__5013 (
            .O(N__28884),
            .I(N__28876));
    LocalMux I__5012 (
            .O(N__28881),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ));
    Odrv4 I__5011 (
            .O(N__28876),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ));
    InMux I__5010 (
            .O(N__28871),
            .I(N__28868));
    LocalMux I__5009 (
            .O(N__28868),
            .I(N__28865));
    Odrv4 I__5008 (
            .O(N__28865),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO ));
    InMux I__5007 (
            .O(N__28862),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ));
    InMux I__5006 (
            .O(N__28859),
            .I(N__28856));
    LocalMux I__5005 (
            .O(N__28856),
            .I(N__28853));
    Odrv4 I__5004 (
            .O(N__28853),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO ));
    InMux I__5003 (
            .O(N__28850),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ));
    CascadeMux I__5002 (
            .O(N__28847),
            .I(N__28844));
    InMux I__5001 (
            .O(N__28844),
            .I(N__28841));
    LocalMux I__5000 (
            .O(N__28841),
            .I(N__28836));
    InMux I__4999 (
            .O(N__28840),
            .I(N__28833));
    InMux I__4998 (
            .O(N__28839),
            .I(N__28830));
    Span4Mux_h I__4997 (
            .O(N__28836),
            .I(N__28827));
    LocalMux I__4996 (
            .O(N__28833),
            .I(N__28824));
    LocalMux I__4995 (
            .O(N__28830),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ));
    Odrv4 I__4994 (
            .O(N__28827),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ));
    Odrv12 I__4993 (
            .O(N__28824),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ));
    InMux I__4992 (
            .O(N__28817),
            .I(N__28814));
    LocalMux I__4991 (
            .O(N__28814),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO ));
    InMux I__4990 (
            .O(N__28811),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ));
    CascadeMux I__4989 (
            .O(N__28808),
            .I(N__28805));
    InMux I__4988 (
            .O(N__28805),
            .I(N__28802));
    LocalMux I__4987 (
            .O(N__28802),
            .I(N__28797));
    InMux I__4986 (
            .O(N__28801),
            .I(N__28794));
    InMux I__4985 (
            .O(N__28800),
            .I(N__28791));
    Span4Mux_v I__4984 (
            .O(N__28797),
            .I(N__28788));
    LocalMux I__4983 (
            .O(N__28794),
            .I(N__28785));
    LocalMux I__4982 (
            .O(N__28791),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ));
    Odrv4 I__4981 (
            .O(N__28788),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ));
    Odrv12 I__4980 (
            .O(N__28785),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ));
    InMux I__4979 (
            .O(N__28778),
            .I(N__28775));
    LocalMux I__4978 (
            .O(N__28775),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO ));
    InMux I__4977 (
            .O(N__28772),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ));
    InMux I__4976 (
            .O(N__28769),
            .I(N__28766));
    LocalMux I__4975 (
            .O(N__28766),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_7 ));
    InMux I__4974 (
            .O(N__28763),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ));
    InMux I__4973 (
            .O(N__28760),
            .I(N__28757));
    LocalMux I__4972 (
            .O(N__28757),
            .I(N__28754));
    Span4Mux_v I__4971 (
            .O(N__28754),
            .I(N__28751));
    Span4Mux_v I__4970 (
            .O(N__28751),
            .I(N__28748));
    Odrv4 I__4969 (
            .O(N__28748),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_8 ));
    InMux I__4968 (
            .O(N__28745),
            .I(bfn_11_11_0_));
    InMux I__4967 (
            .O(N__28742),
            .I(N__28739));
    LocalMux I__4966 (
            .O(N__28739),
            .I(N__28736));
    Span4Mux_h I__4965 (
            .O(N__28736),
            .I(N__28733));
    Odrv4 I__4964 (
            .O(N__28733),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_9 ));
    InMux I__4963 (
            .O(N__28730),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ));
    CascadeMux I__4962 (
            .O(N__28727),
            .I(N__28724));
    InMux I__4961 (
            .O(N__28724),
            .I(N__28721));
    LocalMux I__4960 (
            .O(N__28721),
            .I(N__28718));
    Odrv12 I__4959 (
            .O(N__28718),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_10 ));
    InMux I__4958 (
            .O(N__28715),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ));
    InMux I__4957 (
            .O(N__28712),
            .I(N__28709));
    LocalMux I__4956 (
            .O(N__28709),
            .I(N__28706));
    Span4Mux_h I__4955 (
            .O(N__28706),
            .I(N__28703));
    Odrv4 I__4954 (
            .O(N__28703),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_11 ));
    InMux I__4953 (
            .O(N__28700),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ));
    InMux I__4952 (
            .O(N__28697),
            .I(N__28692));
    InMux I__4951 (
            .O(N__28696),
            .I(N__28689));
    InMux I__4950 (
            .O(N__28695),
            .I(N__28686));
    LocalMux I__4949 (
            .O(N__28692),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ));
    LocalMux I__4948 (
            .O(N__28689),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ));
    LocalMux I__4947 (
            .O(N__28686),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ));
    InMux I__4946 (
            .O(N__28679),
            .I(N__28676));
    LocalMux I__4945 (
            .O(N__28676),
            .I(N__28673));
    Odrv4 I__4944 (
            .O(N__28673),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO ));
    InMux I__4943 (
            .O(N__28670),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ));
    InMux I__4942 (
            .O(N__28667),
            .I(N__28664));
    LocalMux I__4941 (
            .O(N__28664),
            .I(N__28659));
    InMux I__4940 (
            .O(N__28663),
            .I(N__28656));
    InMux I__4939 (
            .O(N__28662),
            .I(N__28653));
    Odrv4 I__4938 (
            .O(N__28659),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ));
    LocalMux I__4937 (
            .O(N__28656),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ));
    LocalMux I__4936 (
            .O(N__28653),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ));
    InMux I__4935 (
            .O(N__28646),
            .I(N__28643));
    LocalMux I__4934 (
            .O(N__28643),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO ));
    InMux I__4933 (
            .O(N__28640),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ));
    InMux I__4932 (
            .O(N__28637),
            .I(N__28632));
    InMux I__4931 (
            .O(N__28636),
            .I(N__28629));
    InMux I__4930 (
            .O(N__28635),
            .I(N__28626));
    LocalMux I__4929 (
            .O(N__28632),
            .I(N__28623));
    LocalMux I__4928 (
            .O(N__28629),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ));
    LocalMux I__4927 (
            .O(N__28626),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ));
    Odrv4 I__4926 (
            .O(N__28623),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ));
    CascadeMux I__4925 (
            .O(N__28616),
            .I(N__28613));
    InMux I__4924 (
            .O(N__28613),
            .I(N__28610));
    LocalMux I__4923 (
            .O(N__28610),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO ));
    InMux I__4922 (
            .O(N__28607),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ));
    CascadeMux I__4921 (
            .O(N__28604),
            .I(N__28601));
    InMux I__4920 (
            .O(N__28601),
            .I(N__28598));
    LocalMux I__4919 (
            .O(N__28598),
            .I(N__28595));
    Span4Mux_h I__4918 (
            .O(N__28595),
            .I(N__28592));
    Odrv4 I__4917 (
            .O(N__28592),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    CascadeMux I__4916 (
            .O(N__28589),
            .I(N__28586));
    InMux I__4915 (
            .O(N__28586),
            .I(N__28583));
    LocalMux I__4914 (
            .O(N__28583),
            .I(N__28580));
    Span4Mux_h I__4913 (
            .O(N__28580),
            .I(N__28577));
    Odrv4 I__4912 (
            .O(N__28577),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    InMux I__4911 (
            .O(N__28574),
            .I(N__28570));
    InMux I__4910 (
            .O(N__28573),
            .I(N__28567));
    LocalMux I__4909 (
            .O(N__28570),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    LocalMux I__4908 (
            .O(N__28567),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    InMux I__4907 (
            .O(N__28562),
            .I(N__28559));
    LocalMux I__4906 (
            .O(N__28559),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ));
    InMux I__4905 (
            .O(N__28556),
            .I(N__28553));
    LocalMux I__4904 (
            .O(N__28553),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ));
    InMux I__4903 (
            .O(N__28550),
            .I(N__28547));
    LocalMux I__4902 (
            .O(N__28547),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ));
    InMux I__4901 (
            .O(N__28544),
            .I(N__28541));
    LocalMux I__4900 (
            .O(N__28541),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ));
    InMux I__4899 (
            .O(N__28538),
            .I(N__28535));
    LocalMux I__4898 (
            .O(N__28535),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_4 ));
    InMux I__4897 (
            .O(N__28532),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ));
    CascadeMux I__4896 (
            .O(N__28529),
            .I(N__28526));
    InMux I__4895 (
            .O(N__28526),
            .I(N__28523));
    LocalMux I__4894 (
            .O(N__28523),
            .I(N__28520));
    Odrv4 I__4893 (
            .O(N__28520),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_5 ));
    InMux I__4892 (
            .O(N__28517),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ));
    InMux I__4891 (
            .O(N__28514),
            .I(N__28511));
    LocalMux I__4890 (
            .O(N__28511),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_6 ));
    InMux I__4889 (
            .O(N__28508),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ));
    InMux I__4888 (
            .O(N__28505),
            .I(N__28502));
    LocalMux I__4887 (
            .O(N__28502),
            .I(N__28499));
    Span4Mux_h I__4886 (
            .O(N__28499),
            .I(N__28496));
    Span4Mux_h I__4885 (
            .O(N__28496),
            .I(N__28493));
    Odrv4 I__4884 (
            .O(N__28493),
            .I(\current_shift_inst.PI_CTRL.integrator_i_19 ));
    CascadeMux I__4883 (
            .O(N__28490),
            .I(N__28487));
    InMux I__4882 (
            .O(N__28487),
            .I(N__28484));
    LocalMux I__4881 (
            .O(N__28484),
            .I(N__28480));
    InMux I__4880 (
            .O(N__28483),
            .I(N__28475));
    Span4Mux_v I__4879 (
            .O(N__28480),
            .I(N__28472));
    CascadeMux I__4878 (
            .O(N__28479),
            .I(N__28469));
    CascadeMux I__4877 (
            .O(N__28478),
            .I(N__28466));
    LocalMux I__4876 (
            .O(N__28475),
            .I(N__28462));
    Span4Mux_h I__4875 (
            .O(N__28472),
            .I(N__28459));
    InMux I__4874 (
            .O(N__28469),
            .I(N__28454));
    InMux I__4873 (
            .O(N__28466),
            .I(N__28454));
    InMux I__4872 (
            .O(N__28465),
            .I(N__28451));
    Odrv4 I__4871 (
            .O(N__28462),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__4870 (
            .O(N__28459),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    LocalMux I__4869 (
            .O(N__28454),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    LocalMux I__4868 (
            .O(N__28451),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    CascadeMux I__4867 (
            .O(N__28442),
            .I(N__28439));
    InMux I__4866 (
            .O(N__28439),
            .I(N__28436));
    LocalMux I__4865 (
            .O(N__28436),
            .I(N__28433));
    Span4Mux_v I__4864 (
            .O(N__28433),
            .I(N__28430));
    Odrv4 I__4863 (
            .O(N__28430),
            .I(\current_shift_inst.PI_CTRL.integrator_i_12 ));
    InMux I__4862 (
            .O(N__28427),
            .I(N__28423));
    InMux I__4861 (
            .O(N__28426),
            .I(N__28420));
    LocalMux I__4860 (
            .O(N__28423),
            .I(N__28416));
    LocalMux I__4859 (
            .O(N__28420),
            .I(N__28412));
    CascadeMux I__4858 (
            .O(N__28419),
            .I(N__28409));
    Span4Mux_v I__4857 (
            .O(N__28416),
            .I(N__28405));
    InMux I__4856 (
            .O(N__28415),
            .I(N__28402));
    Span4Mux_h I__4855 (
            .O(N__28412),
            .I(N__28399));
    InMux I__4854 (
            .O(N__28409),
            .I(N__28396));
    InMux I__4853 (
            .O(N__28408),
            .I(N__28393));
    Odrv4 I__4852 (
            .O(N__28405),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    LocalMux I__4851 (
            .O(N__28402),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__4850 (
            .O(N__28399),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    LocalMux I__4849 (
            .O(N__28396),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    LocalMux I__4848 (
            .O(N__28393),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    CascadeMux I__4847 (
            .O(N__28382),
            .I(N__28379));
    InMux I__4846 (
            .O(N__28379),
            .I(N__28376));
    LocalMux I__4845 (
            .O(N__28376),
            .I(N__28373));
    Odrv4 I__4844 (
            .O(N__28373),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10 ));
    CascadeMux I__4843 (
            .O(N__28370),
            .I(N__28367));
    InMux I__4842 (
            .O(N__28367),
            .I(N__28364));
    LocalMux I__4841 (
            .O(N__28364),
            .I(N__28361));
    Odrv4 I__4840 (
            .O(N__28361),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5 ));
    InMux I__4839 (
            .O(N__28358),
            .I(N__28355));
    LocalMux I__4838 (
            .O(N__28355),
            .I(N__28352));
    Span4Mux_h I__4837 (
            .O(N__28352),
            .I(N__28349));
    Odrv4 I__4836 (
            .O(N__28349),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ));
    InMux I__4835 (
            .O(N__28346),
            .I(N__28343));
    LocalMux I__4834 (
            .O(N__28343),
            .I(N__28340));
    Odrv12 I__4833 (
            .O(N__28340),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    InMux I__4832 (
            .O(N__28337),
            .I(N__28334));
    LocalMux I__4831 (
            .O(N__28334),
            .I(N__28331));
    Odrv12 I__4830 (
            .O(N__28331),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    InMux I__4829 (
            .O(N__28328),
            .I(N__28325));
    LocalMux I__4828 (
            .O(N__28325),
            .I(N__28322));
    Odrv4 I__4827 (
            .O(N__28322),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    CascadeMux I__4826 (
            .O(N__28319),
            .I(N__28310));
    InMux I__4825 (
            .O(N__28318),
            .I(N__28293));
    InMux I__4824 (
            .O(N__28317),
            .I(N__28290));
    InMux I__4823 (
            .O(N__28316),
            .I(N__28281));
    InMux I__4822 (
            .O(N__28315),
            .I(N__28281));
    InMux I__4821 (
            .O(N__28314),
            .I(N__28281));
    InMux I__4820 (
            .O(N__28313),
            .I(N__28281));
    InMux I__4819 (
            .O(N__28310),
            .I(N__28270));
    InMux I__4818 (
            .O(N__28309),
            .I(N__28270));
    InMux I__4817 (
            .O(N__28308),
            .I(N__28270));
    InMux I__4816 (
            .O(N__28307),
            .I(N__28270));
    InMux I__4815 (
            .O(N__28306),
            .I(N__28270));
    InMux I__4814 (
            .O(N__28305),
            .I(N__28257));
    InMux I__4813 (
            .O(N__28304),
            .I(N__28246));
    InMux I__4812 (
            .O(N__28303),
            .I(N__28246));
    InMux I__4811 (
            .O(N__28302),
            .I(N__28246));
    InMux I__4810 (
            .O(N__28301),
            .I(N__28246));
    InMux I__4809 (
            .O(N__28300),
            .I(N__28246));
    InMux I__4808 (
            .O(N__28299),
            .I(N__28237));
    InMux I__4807 (
            .O(N__28298),
            .I(N__28237));
    InMux I__4806 (
            .O(N__28297),
            .I(N__28237));
    InMux I__4805 (
            .O(N__28296),
            .I(N__28237));
    LocalMux I__4804 (
            .O(N__28293),
            .I(N__28234));
    LocalMux I__4803 (
            .O(N__28290),
            .I(N__28230));
    LocalMux I__4802 (
            .O(N__28281),
            .I(N__28225));
    LocalMux I__4801 (
            .O(N__28270),
            .I(N__28225));
    InMux I__4800 (
            .O(N__28269),
            .I(N__28222));
    InMux I__4799 (
            .O(N__28268),
            .I(N__28211));
    InMux I__4798 (
            .O(N__28267),
            .I(N__28211));
    InMux I__4797 (
            .O(N__28266),
            .I(N__28211));
    InMux I__4796 (
            .O(N__28265),
            .I(N__28211));
    InMux I__4795 (
            .O(N__28264),
            .I(N__28211));
    InMux I__4794 (
            .O(N__28263),
            .I(N__28202));
    InMux I__4793 (
            .O(N__28262),
            .I(N__28202));
    InMux I__4792 (
            .O(N__28261),
            .I(N__28202));
    InMux I__4791 (
            .O(N__28260),
            .I(N__28202));
    LocalMux I__4790 (
            .O(N__28257),
            .I(N__28199));
    LocalMux I__4789 (
            .O(N__28246),
            .I(N__28194));
    LocalMux I__4788 (
            .O(N__28237),
            .I(N__28194));
    Span4Mux_v I__4787 (
            .O(N__28234),
            .I(N__28191));
    InMux I__4786 (
            .O(N__28233),
            .I(N__28188));
    Span4Mux_h I__4785 (
            .O(N__28230),
            .I(N__28183));
    Span4Mux_h I__4784 (
            .O(N__28225),
            .I(N__28183));
    LocalMux I__4783 (
            .O(N__28222),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__4782 (
            .O(N__28211),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__4781 (
            .O(N__28202),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__4780 (
            .O(N__28199),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__4779 (
            .O(N__28194),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__4778 (
            .O(N__28191),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__4777 (
            .O(N__28188),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__4776 (
            .O(N__28183),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    CascadeMux I__4775 (
            .O(N__28166),
            .I(N__28153));
    CascadeMux I__4774 (
            .O(N__28165),
            .I(N__28140));
    CascadeMux I__4773 (
            .O(N__28164),
            .I(N__28136));
    CascadeMux I__4772 (
            .O(N__28163),
            .I(N__28133));
    CascadeMux I__4771 (
            .O(N__28162),
            .I(N__28130));
    CascadeMux I__4770 (
            .O(N__28161),
            .I(N__28126));
    CascadeMux I__4769 (
            .O(N__28160),
            .I(N__28123));
    InMux I__4768 (
            .O(N__28159),
            .I(N__28114));
    InMux I__4767 (
            .O(N__28158),
            .I(N__28114));
    InMux I__4766 (
            .O(N__28157),
            .I(N__28114));
    InMux I__4765 (
            .O(N__28156),
            .I(N__28114));
    InMux I__4764 (
            .O(N__28153),
            .I(N__28111));
    CascadeMux I__4763 (
            .O(N__28152),
            .I(N__28108));
    CascadeMux I__4762 (
            .O(N__28151),
            .I(N__28105));
    CascadeMux I__4761 (
            .O(N__28150),
            .I(N__28102));
    CascadeMux I__4760 (
            .O(N__28149),
            .I(N__28095));
    CascadeMux I__4759 (
            .O(N__28148),
            .I(N__28092));
    CascadeMux I__4758 (
            .O(N__28147),
            .I(N__28089));
    CascadeMux I__4757 (
            .O(N__28146),
            .I(N__28086));
    InMux I__4756 (
            .O(N__28145),
            .I(N__28077));
    InMux I__4755 (
            .O(N__28144),
            .I(N__28077));
    InMux I__4754 (
            .O(N__28143),
            .I(N__28077));
    InMux I__4753 (
            .O(N__28140),
            .I(N__28077));
    InMux I__4752 (
            .O(N__28139),
            .I(N__28068));
    InMux I__4751 (
            .O(N__28136),
            .I(N__28068));
    InMux I__4750 (
            .O(N__28133),
            .I(N__28068));
    InMux I__4749 (
            .O(N__28130),
            .I(N__28068));
    InMux I__4748 (
            .O(N__28129),
            .I(N__28061));
    InMux I__4747 (
            .O(N__28126),
            .I(N__28061));
    InMux I__4746 (
            .O(N__28123),
            .I(N__28061));
    LocalMux I__4745 (
            .O(N__28114),
            .I(N__28056));
    LocalMux I__4744 (
            .O(N__28111),
            .I(N__28056));
    InMux I__4743 (
            .O(N__28108),
            .I(N__28053));
    InMux I__4742 (
            .O(N__28105),
            .I(N__28046));
    InMux I__4741 (
            .O(N__28102),
            .I(N__28046));
    InMux I__4740 (
            .O(N__28101),
            .I(N__28046));
    InMux I__4739 (
            .O(N__28100),
            .I(N__28035));
    InMux I__4738 (
            .O(N__28099),
            .I(N__28035));
    InMux I__4737 (
            .O(N__28098),
            .I(N__28035));
    InMux I__4736 (
            .O(N__28095),
            .I(N__28035));
    InMux I__4735 (
            .O(N__28092),
            .I(N__28035));
    InMux I__4734 (
            .O(N__28089),
            .I(N__28030));
    InMux I__4733 (
            .O(N__28086),
            .I(N__28030));
    LocalMux I__4732 (
            .O(N__28077),
            .I(N__28027));
    LocalMux I__4731 (
            .O(N__28068),
            .I(N__28024));
    LocalMux I__4730 (
            .O(N__28061),
            .I(N__28019));
    Span4Mux_v I__4729 (
            .O(N__28056),
            .I(N__28019));
    LocalMux I__4728 (
            .O(N__28053),
            .I(\current_shift_inst.PI_CTRL.N_103 ));
    LocalMux I__4727 (
            .O(N__28046),
            .I(\current_shift_inst.PI_CTRL.N_103 ));
    LocalMux I__4726 (
            .O(N__28035),
            .I(\current_shift_inst.PI_CTRL.N_103 ));
    LocalMux I__4725 (
            .O(N__28030),
            .I(\current_shift_inst.PI_CTRL.N_103 ));
    Odrv4 I__4724 (
            .O(N__28027),
            .I(\current_shift_inst.PI_CTRL.N_103 ));
    Odrv4 I__4723 (
            .O(N__28024),
            .I(\current_shift_inst.PI_CTRL.N_103 ));
    Odrv4 I__4722 (
            .O(N__28019),
            .I(\current_shift_inst.PI_CTRL.N_103 ));
    InMux I__4721 (
            .O(N__28004),
            .I(N__27985));
    InMux I__4720 (
            .O(N__28003),
            .I(N__27985));
    InMux I__4719 (
            .O(N__28002),
            .I(N__27985));
    InMux I__4718 (
            .O(N__28001),
            .I(N__27985));
    InMux I__4717 (
            .O(N__28000),
            .I(N__27985));
    CascadeMux I__4716 (
            .O(N__27999),
            .I(N__27971));
    CascadeMux I__4715 (
            .O(N__27998),
            .I(N__27968));
    InMux I__4714 (
            .O(N__27997),
            .I(N__27962));
    CascadeMux I__4713 (
            .O(N__27996),
            .I(N__27957));
    LocalMux I__4712 (
            .O(N__27985),
            .I(N__27948));
    InMux I__4711 (
            .O(N__27984),
            .I(N__27939));
    InMux I__4710 (
            .O(N__27983),
            .I(N__27939));
    InMux I__4709 (
            .O(N__27982),
            .I(N__27939));
    InMux I__4708 (
            .O(N__27981),
            .I(N__27939));
    CascadeMux I__4707 (
            .O(N__27980),
            .I(N__27936));
    CascadeMux I__4706 (
            .O(N__27979),
            .I(N__27932));
    CascadeMux I__4705 (
            .O(N__27978),
            .I(N__27929));
    InMux I__4704 (
            .O(N__27977),
            .I(N__27926));
    InMux I__4703 (
            .O(N__27976),
            .I(N__27921));
    InMux I__4702 (
            .O(N__27975),
            .I(N__27921));
    InMux I__4701 (
            .O(N__27974),
            .I(N__27912));
    InMux I__4700 (
            .O(N__27971),
            .I(N__27912));
    InMux I__4699 (
            .O(N__27968),
            .I(N__27912));
    InMux I__4698 (
            .O(N__27967),
            .I(N__27912));
    InMux I__4697 (
            .O(N__27966),
            .I(N__27907));
    InMux I__4696 (
            .O(N__27965),
            .I(N__27907));
    LocalMux I__4695 (
            .O(N__27962),
            .I(N__27904));
    InMux I__4694 (
            .O(N__27961),
            .I(N__27901));
    InMux I__4693 (
            .O(N__27960),
            .I(N__27892));
    InMux I__4692 (
            .O(N__27957),
            .I(N__27892));
    InMux I__4691 (
            .O(N__27956),
            .I(N__27892));
    InMux I__4690 (
            .O(N__27955),
            .I(N__27892));
    InMux I__4689 (
            .O(N__27954),
            .I(N__27883));
    InMux I__4688 (
            .O(N__27953),
            .I(N__27883));
    InMux I__4687 (
            .O(N__27952),
            .I(N__27883));
    InMux I__4686 (
            .O(N__27951),
            .I(N__27883));
    Span4Mux_v I__4685 (
            .O(N__27948),
            .I(N__27878));
    LocalMux I__4684 (
            .O(N__27939),
            .I(N__27878));
    InMux I__4683 (
            .O(N__27936),
            .I(N__27875));
    InMux I__4682 (
            .O(N__27935),
            .I(N__27868));
    InMux I__4681 (
            .O(N__27932),
            .I(N__27868));
    InMux I__4680 (
            .O(N__27929),
            .I(N__27868));
    LocalMux I__4679 (
            .O(N__27926),
            .I(N__27865));
    LocalMux I__4678 (
            .O(N__27921),
            .I(N__27856));
    LocalMux I__4677 (
            .O(N__27912),
            .I(N__27856));
    LocalMux I__4676 (
            .O(N__27907),
            .I(N__27856));
    Span4Mux_v I__4675 (
            .O(N__27904),
            .I(N__27856));
    LocalMux I__4674 (
            .O(N__27901),
            .I(N__27847));
    LocalMux I__4673 (
            .O(N__27892),
            .I(N__27847));
    LocalMux I__4672 (
            .O(N__27883),
            .I(N__27847));
    Span4Mux_v I__4671 (
            .O(N__27878),
            .I(N__27847));
    LocalMux I__4670 (
            .O(N__27875),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    LocalMux I__4669 (
            .O(N__27868),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    Odrv4 I__4668 (
            .O(N__27865),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    Odrv4 I__4667 (
            .O(N__27856),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    Odrv4 I__4666 (
            .O(N__27847),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    CascadeMux I__4665 (
            .O(N__27836),
            .I(N__27833));
    InMux I__4664 (
            .O(N__27833),
            .I(N__27828));
    InMux I__4663 (
            .O(N__27832),
            .I(N__27825));
    InMux I__4662 (
            .O(N__27831),
            .I(N__27822));
    LocalMux I__4661 (
            .O(N__27828),
            .I(N__27810));
    LocalMux I__4660 (
            .O(N__27825),
            .I(N__27810));
    LocalMux I__4659 (
            .O(N__27822),
            .I(N__27810));
    InMux I__4658 (
            .O(N__27821),
            .I(N__27805));
    InMux I__4657 (
            .O(N__27820),
            .I(N__27805));
    InMux I__4656 (
            .O(N__27819),
            .I(N__27802));
    InMux I__4655 (
            .O(N__27818),
            .I(N__27799));
    InMux I__4654 (
            .O(N__27817),
            .I(N__27796));
    Span4Mux_v I__4653 (
            .O(N__27810),
            .I(N__27793));
    LocalMux I__4652 (
            .O(N__27805),
            .I(elapsed_time_ns_1_RNIS4MD11_0_15));
    LocalMux I__4651 (
            .O(N__27802),
            .I(elapsed_time_ns_1_RNIS4MD11_0_15));
    LocalMux I__4650 (
            .O(N__27799),
            .I(elapsed_time_ns_1_RNIS4MD11_0_15));
    LocalMux I__4649 (
            .O(N__27796),
            .I(elapsed_time_ns_1_RNIS4MD11_0_15));
    Odrv4 I__4648 (
            .O(N__27793),
            .I(elapsed_time_ns_1_RNIS4MD11_0_15));
    InMux I__4647 (
            .O(N__27782),
            .I(N__27778));
    InMux I__4646 (
            .O(N__27781),
            .I(N__27775));
    LocalMux I__4645 (
            .O(N__27778),
            .I(N__27772));
    LocalMux I__4644 (
            .O(N__27775),
            .I(N__27769));
    Span4Mux_v I__4643 (
            .O(N__27772),
            .I(N__27766));
    Odrv4 I__4642 (
            .O(N__27769),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_CO ));
    Odrv4 I__4641 (
            .O(N__27766),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_CO ));
    InMux I__4640 (
            .O(N__27761),
            .I(N__27758));
    LocalMux I__4639 (
            .O(N__27758),
            .I(N__27755));
    Odrv12 I__4638 (
            .O(N__27755),
            .I(\phase_controller_inst2.stoper_hc.running_1_sqmuxa ));
    InMux I__4637 (
            .O(N__27752),
            .I(N__27744));
    InMux I__4636 (
            .O(N__27751),
            .I(N__27744));
    CascadeMux I__4635 (
            .O(N__27750),
            .I(N__27740));
    InMux I__4634 (
            .O(N__27749),
            .I(N__27735));
    LocalMux I__4633 (
            .O(N__27744),
            .I(N__27732));
    InMux I__4632 (
            .O(N__27743),
            .I(N__27725));
    InMux I__4631 (
            .O(N__27740),
            .I(N__27725));
    InMux I__4630 (
            .O(N__27739),
            .I(N__27725));
    InMux I__4629 (
            .O(N__27738),
            .I(N__27722));
    LocalMux I__4628 (
            .O(N__27735),
            .I(N__27719));
    Span4Mux_h I__4627 (
            .O(N__27732),
            .I(N__27714));
    LocalMux I__4626 (
            .O(N__27725),
            .I(N__27714));
    LocalMux I__4625 (
            .O(N__27722),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv12 I__4624 (
            .O(N__27719),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv4 I__4623 (
            .O(N__27714),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    InMux I__4622 (
            .O(N__27707),
            .I(N__27700));
    InMux I__4621 (
            .O(N__27706),
            .I(N__27700));
    InMux I__4620 (
            .O(N__27705),
            .I(N__27693));
    LocalMux I__4619 (
            .O(N__27700),
            .I(N__27690));
    InMux I__4618 (
            .O(N__27699),
            .I(N__27681));
    InMux I__4617 (
            .O(N__27698),
            .I(N__27681));
    InMux I__4616 (
            .O(N__27697),
            .I(N__27681));
    InMux I__4615 (
            .O(N__27696),
            .I(N__27681));
    LocalMux I__4614 (
            .O(N__27693),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    Odrv4 I__4613 (
            .O(N__27690),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    LocalMux I__4612 (
            .O(N__27681),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    CascadeMux I__4611 (
            .O(N__27674),
            .I(\phase_controller_inst2.stoper_hc.running_1_sqmuxa_cascade_ ));
    InMux I__4610 (
            .O(N__27671),
            .I(N__27668));
    LocalMux I__4609 (
            .O(N__27668),
            .I(N__27663));
    InMux I__4608 (
            .O(N__27667),
            .I(N__27658));
    InMux I__4607 (
            .O(N__27666),
            .I(N__27658));
    Odrv4 I__4606 (
            .O(N__27663),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    LocalMux I__4605 (
            .O(N__27658),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    InMux I__4604 (
            .O(N__27653),
            .I(N__27650));
    LocalMux I__4603 (
            .O(N__27650),
            .I(N__27647));
    Odrv12 I__4602 (
            .O(N__27647),
            .I(\phase_controller_inst2.stoper_hc.un1_start_latched2_0 ));
    IoInMux I__4601 (
            .O(N__27644),
            .I(N__27641));
    LocalMux I__4600 (
            .O(N__27641),
            .I(N__27638));
    Span4Mux_s2_v I__4599 (
            .O(N__27638),
            .I(N__27635));
    Span4Mux_v I__4598 (
            .O(N__27635),
            .I(N__27632));
    Odrv4 I__4597 (
            .O(N__27632),
            .I(s4_phy_c));
    InMux I__4596 (
            .O(N__27629),
            .I(N__27626));
    LocalMux I__4595 (
            .O(N__27626),
            .I(N__27623));
    Odrv4 I__4594 (
            .O(N__27623),
            .I(il_max_comp1_D1));
    InMux I__4593 (
            .O(N__27620),
            .I(N__27617));
    LocalMux I__4592 (
            .O(N__27617),
            .I(N__27614));
    Span4Mux_v I__4591 (
            .O(N__27614),
            .I(N__27611));
    Span4Mux_h I__4590 (
            .O(N__27611),
            .I(N__27608));
    Odrv4 I__4589 (
            .O(N__27608),
            .I(il_min_comp2_c));
    InMux I__4588 (
            .O(N__27605),
            .I(N__27602));
    LocalMux I__4587 (
            .O(N__27602),
            .I(il_min_comp2_D1));
    InMux I__4586 (
            .O(N__27599),
            .I(N__27592));
    InMux I__4585 (
            .O(N__27598),
            .I(N__27589));
    CascadeMux I__4584 (
            .O(N__27597),
            .I(N__27586));
    CascadeMux I__4583 (
            .O(N__27596),
            .I(N__27583));
    InMux I__4582 (
            .O(N__27595),
            .I(N__27580));
    LocalMux I__4581 (
            .O(N__27592),
            .I(N__27577));
    LocalMux I__4580 (
            .O(N__27589),
            .I(N__27574));
    InMux I__4579 (
            .O(N__27586),
            .I(N__27571));
    InMux I__4578 (
            .O(N__27583),
            .I(N__27568));
    LocalMux I__4577 (
            .O(N__27580),
            .I(N__27565));
    Span4Mux_v I__4576 (
            .O(N__27577),
            .I(N__27562));
    Span4Mux_v I__4575 (
            .O(N__27574),
            .I(N__27555));
    LocalMux I__4574 (
            .O(N__27571),
            .I(N__27555));
    LocalMux I__4573 (
            .O(N__27568),
            .I(N__27555));
    Span4Mux_h I__4572 (
            .O(N__27565),
            .I(N__27552));
    Odrv4 I__4571 (
            .O(N__27562),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__4570 (
            .O(N__27555),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__4569 (
            .O(N__27552),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    InMux I__4568 (
            .O(N__27545),
            .I(N__27542));
    LocalMux I__4567 (
            .O(N__27542),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_5 ));
    CascadeMux I__4566 (
            .O(N__27539),
            .I(N__27536));
    InMux I__4565 (
            .O(N__27536),
            .I(N__27533));
    LocalMux I__4564 (
            .O(N__27533),
            .I(N__27530));
    Span4Mux_h I__4563 (
            .O(N__27530),
            .I(N__27526));
    InMux I__4562 (
            .O(N__27529),
            .I(N__27522));
    Span4Mux_h I__4561 (
            .O(N__27526),
            .I(N__27519));
    InMux I__4560 (
            .O(N__27525),
            .I(N__27516));
    LocalMux I__4559 (
            .O(N__27522),
            .I(elapsed_time_ns_1_RNINVLD11_0_10));
    Odrv4 I__4558 (
            .O(N__27519),
            .I(elapsed_time_ns_1_RNINVLD11_0_10));
    LocalMux I__4557 (
            .O(N__27516),
            .I(elapsed_time_ns_1_RNINVLD11_0_10));
    InMux I__4556 (
            .O(N__27509),
            .I(N__27506));
    LocalMux I__4555 (
            .O(N__27506),
            .I(N__27500));
    CascadeMux I__4554 (
            .O(N__27505),
            .I(N__27497));
    InMux I__4553 (
            .O(N__27504),
            .I(N__27494));
    InMux I__4552 (
            .O(N__27503),
            .I(N__27491));
    Span4Mux_h I__4551 (
            .O(N__27500),
            .I(N__27488));
    InMux I__4550 (
            .O(N__27497),
            .I(N__27485));
    LocalMux I__4549 (
            .O(N__27494),
            .I(N__27482));
    LocalMux I__4548 (
            .O(N__27491),
            .I(elapsed_time_ns_1_RNIQ2MD11_0_13));
    Odrv4 I__4547 (
            .O(N__27488),
            .I(elapsed_time_ns_1_RNIQ2MD11_0_13));
    LocalMux I__4546 (
            .O(N__27485),
            .I(elapsed_time_ns_1_RNIQ2MD11_0_13));
    Odrv4 I__4545 (
            .O(N__27482),
            .I(elapsed_time_ns_1_RNIQ2MD11_0_13));
    CascadeMux I__4544 (
            .O(N__27473),
            .I(elapsed_time_ns_1_RNINVLD11_0_10_cascade_));
    CascadeMux I__4543 (
            .O(N__27470),
            .I(N__27466));
    CascadeMux I__4542 (
            .O(N__27469),
            .I(N__27463));
    InMux I__4541 (
            .O(N__27466),
            .I(N__27460));
    InMux I__4540 (
            .O(N__27463),
            .I(N__27457));
    LocalMux I__4539 (
            .O(N__27460),
            .I(N__27454));
    LocalMux I__4538 (
            .O(N__27457),
            .I(N__27449));
    Span4Mux_h I__4537 (
            .O(N__27454),
            .I(N__27449));
    Span4Mux_h I__4536 (
            .O(N__27449),
            .I(N__27444));
    InMux I__4535 (
            .O(N__27448),
            .I(N__27439));
    InMux I__4534 (
            .O(N__27447),
            .I(N__27439));
    Odrv4 I__4533 (
            .O(N__27444),
            .I(elapsed_time_ns_1_RNIP1MD11_0_12));
    LocalMux I__4532 (
            .O(N__27439),
            .I(elapsed_time_ns_1_RNIP1MD11_0_12));
    CascadeMux I__4531 (
            .O(N__27434),
            .I(\phase_controller_inst1.stoper_hc.N_319_cascade_ ));
    CascadeMux I__4530 (
            .O(N__27431),
            .I(N__27428));
    InMux I__4529 (
            .O(N__27428),
            .I(N__27423));
    InMux I__4528 (
            .O(N__27427),
            .I(N__27420));
    InMux I__4527 (
            .O(N__27426),
            .I(N__27417));
    LocalMux I__4526 (
            .O(N__27423),
            .I(N__27413));
    LocalMux I__4525 (
            .O(N__27420),
            .I(N__27408));
    LocalMux I__4524 (
            .O(N__27417),
            .I(N__27408));
    InMux I__4523 (
            .O(N__27416),
            .I(N__27405));
    Span12Mux_s10_h I__4522 (
            .O(N__27413),
            .I(N__27400));
    Sp12to4 I__4521 (
            .O(N__27408),
            .I(N__27395));
    LocalMux I__4520 (
            .O(N__27405),
            .I(N__27395));
    InMux I__4519 (
            .O(N__27404),
            .I(N__27390));
    InMux I__4518 (
            .O(N__27403),
            .I(N__27390));
    Odrv12 I__4517 (
            .O(N__27400),
            .I(elapsed_time_ns_1_RNI1TBED1_0_14));
    Odrv12 I__4516 (
            .O(N__27395),
            .I(elapsed_time_ns_1_RNI1TBED1_0_14));
    LocalMux I__4515 (
            .O(N__27390),
            .I(elapsed_time_ns_1_RNI1TBED1_0_14));
    InMux I__4514 (
            .O(N__27383),
            .I(N__27380));
    LocalMux I__4513 (
            .O(N__27380),
            .I(\phase_controller_inst1.stoper_hc.N_275 ));
    InMux I__4512 (
            .O(N__27377),
            .I(N__27373));
    InMux I__4511 (
            .O(N__27376),
            .I(N__27370));
    LocalMux I__4510 (
            .O(N__27373),
            .I(\phase_controller_inst1.stoper_hc.N_319 ));
    LocalMux I__4509 (
            .O(N__27370),
            .I(\phase_controller_inst1.stoper_hc.N_319 ));
    InMux I__4508 (
            .O(N__27365),
            .I(N__27362));
    LocalMux I__4507 (
            .O(N__27362),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_a5_1_0Z0Z_9 ));
    CascadeMux I__4506 (
            .O(N__27359),
            .I(N__27351));
    InMux I__4505 (
            .O(N__27358),
            .I(N__27333));
    InMux I__4504 (
            .O(N__27357),
            .I(N__27326));
    InMux I__4503 (
            .O(N__27356),
            .I(N__27326));
    InMux I__4502 (
            .O(N__27355),
            .I(N__27326));
    InMux I__4501 (
            .O(N__27354),
            .I(N__27315));
    InMux I__4500 (
            .O(N__27351),
            .I(N__27315));
    InMux I__4499 (
            .O(N__27350),
            .I(N__27315));
    InMux I__4498 (
            .O(N__27349),
            .I(N__27315));
    InMux I__4497 (
            .O(N__27348),
            .I(N__27315));
    InMux I__4496 (
            .O(N__27347),
            .I(N__27306));
    InMux I__4495 (
            .O(N__27346),
            .I(N__27306));
    InMux I__4494 (
            .O(N__27345),
            .I(N__27306));
    InMux I__4493 (
            .O(N__27344),
            .I(N__27306));
    CascadeMux I__4492 (
            .O(N__27343),
            .I(N__27301));
    InMux I__4491 (
            .O(N__27342),
            .I(N__27277));
    InMux I__4490 (
            .O(N__27341),
            .I(N__27277));
    InMux I__4489 (
            .O(N__27340),
            .I(N__27277));
    InMux I__4488 (
            .O(N__27339),
            .I(N__27277));
    InMux I__4487 (
            .O(N__27338),
            .I(N__27277));
    InMux I__4486 (
            .O(N__27337),
            .I(N__27277));
    InMux I__4485 (
            .O(N__27336),
            .I(N__27277));
    LocalMux I__4484 (
            .O(N__27333),
            .I(N__27270));
    LocalMux I__4483 (
            .O(N__27326),
            .I(N__27270));
    LocalMux I__4482 (
            .O(N__27315),
            .I(N__27270));
    LocalMux I__4481 (
            .O(N__27306),
            .I(N__27267));
    InMux I__4480 (
            .O(N__27305),
            .I(N__27263));
    InMux I__4479 (
            .O(N__27304),
            .I(N__27256));
    InMux I__4478 (
            .O(N__27301),
            .I(N__27256));
    InMux I__4477 (
            .O(N__27300),
            .I(N__27256));
    CascadeMux I__4476 (
            .O(N__27299),
            .I(N__27252));
    InMux I__4475 (
            .O(N__27298),
            .I(N__27248));
    InMux I__4474 (
            .O(N__27297),
            .I(N__27235));
    InMux I__4473 (
            .O(N__27296),
            .I(N__27235));
    InMux I__4472 (
            .O(N__27295),
            .I(N__27235));
    InMux I__4471 (
            .O(N__27294),
            .I(N__27235));
    InMux I__4470 (
            .O(N__27293),
            .I(N__27235));
    InMux I__4469 (
            .O(N__27292),
            .I(N__27235));
    LocalMux I__4468 (
            .O(N__27277),
            .I(N__27232));
    Sp12to4 I__4467 (
            .O(N__27270),
            .I(N__27227));
    Span12Mux_s9_h I__4466 (
            .O(N__27267),
            .I(N__27227));
    InMux I__4465 (
            .O(N__27266),
            .I(N__27224));
    LocalMux I__4464 (
            .O(N__27263),
            .I(N__27219));
    LocalMux I__4463 (
            .O(N__27256),
            .I(N__27219));
    InMux I__4462 (
            .O(N__27255),
            .I(N__27212));
    InMux I__4461 (
            .O(N__27252),
            .I(N__27212));
    InMux I__4460 (
            .O(N__27251),
            .I(N__27212));
    LocalMux I__4459 (
            .O(N__27248),
            .I(elapsed_time_ns_1_RNIQ4OD11_0_31));
    LocalMux I__4458 (
            .O(N__27235),
            .I(elapsed_time_ns_1_RNIQ4OD11_0_31));
    Odrv4 I__4457 (
            .O(N__27232),
            .I(elapsed_time_ns_1_RNIQ4OD11_0_31));
    Odrv12 I__4456 (
            .O(N__27227),
            .I(elapsed_time_ns_1_RNIQ4OD11_0_31));
    LocalMux I__4455 (
            .O(N__27224),
            .I(elapsed_time_ns_1_RNIQ4OD11_0_31));
    Odrv4 I__4454 (
            .O(N__27219),
            .I(elapsed_time_ns_1_RNIQ4OD11_0_31));
    LocalMux I__4453 (
            .O(N__27212),
            .I(elapsed_time_ns_1_RNIQ4OD11_0_31));
    CascadeMux I__4452 (
            .O(N__27197),
            .I(N__27193));
    InMux I__4451 (
            .O(N__27196),
            .I(N__27189));
    InMux I__4450 (
            .O(N__27193),
            .I(N__27185));
    InMux I__4449 (
            .O(N__27192),
            .I(N__27182));
    LocalMux I__4448 (
            .O(N__27189),
            .I(N__27179));
    InMux I__4447 (
            .O(N__27188),
            .I(N__27176));
    LocalMux I__4446 (
            .O(N__27185),
            .I(N__27171));
    LocalMux I__4445 (
            .O(N__27182),
            .I(N__27171));
    Odrv4 I__4444 (
            .O(N__27179),
            .I(\phase_controller_inst1.stoper_hc.N_278 ));
    LocalMux I__4443 (
            .O(N__27176),
            .I(\phase_controller_inst1.stoper_hc.N_278 ));
    Odrv4 I__4442 (
            .O(N__27171),
            .I(\phase_controller_inst1.stoper_hc.N_278 ));
    InMux I__4441 (
            .O(N__27164),
            .I(N__27151));
    InMux I__4440 (
            .O(N__27163),
            .I(N__27151));
    InMux I__4439 (
            .O(N__27162),
            .I(N__27151));
    InMux I__4438 (
            .O(N__27161),
            .I(N__27151));
    CascadeMux I__4437 (
            .O(N__27160),
            .I(N__27143));
    LocalMux I__4436 (
            .O(N__27151),
            .I(N__27139));
    InMux I__4435 (
            .O(N__27150),
            .I(N__27136));
    InMux I__4434 (
            .O(N__27149),
            .I(N__27133));
    InMux I__4433 (
            .O(N__27148),
            .I(N__27126));
    InMux I__4432 (
            .O(N__27147),
            .I(N__27126));
    InMux I__4431 (
            .O(N__27146),
            .I(N__27126));
    InMux I__4430 (
            .O(N__27143),
            .I(N__27123));
    InMux I__4429 (
            .O(N__27142),
            .I(N__27107));
    Span4Mux_h I__4428 (
            .O(N__27139),
            .I(N__27102));
    LocalMux I__4427 (
            .O(N__27136),
            .I(N__27093));
    LocalMux I__4426 (
            .O(N__27133),
            .I(N__27093));
    LocalMux I__4425 (
            .O(N__27126),
            .I(N__27093));
    LocalMux I__4424 (
            .O(N__27123),
            .I(N__27093));
    InMux I__4423 (
            .O(N__27122),
            .I(N__27090));
    InMux I__4422 (
            .O(N__27121),
            .I(N__27085));
    InMux I__4421 (
            .O(N__27120),
            .I(N__27085));
    InMux I__4420 (
            .O(N__27119),
            .I(N__27076));
    InMux I__4419 (
            .O(N__27118),
            .I(N__27076));
    InMux I__4418 (
            .O(N__27117),
            .I(N__27076));
    InMux I__4417 (
            .O(N__27116),
            .I(N__27076));
    InMux I__4416 (
            .O(N__27115),
            .I(N__27063));
    InMux I__4415 (
            .O(N__27114),
            .I(N__27063));
    InMux I__4414 (
            .O(N__27113),
            .I(N__27063));
    InMux I__4413 (
            .O(N__27112),
            .I(N__27063));
    InMux I__4412 (
            .O(N__27111),
            .I(N__27063));
    InMux I__4411 (
            .O(N__27110),
            .I(N__27063));
    LocalMux I__4410 (
            .O(N__27107),
            .I(N__27060));
    InMux I__4409 (
            .O(N__27106),
            .I(N__27055));
    InMux I__4408 (
            .O(N__27105),
            .I(N__27055));
    Span4Mux_h I__4407 (
            .O(N__27102),
            .I(N__27050));
    Span4Mux_v I__4406 (
            .O(N__27093),
            .I(N__27050));
    LocalMux I__4405 (
            .O(N__27090),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ));
    LocalMux I__4404 (
            .O(N__27085),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ));
    LocalMux I__4403 (
            .O(N__27076),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ));
    LocalMux I__4402 (
            .O(N__27063),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ));
    Odrv12 I__4401 (
            .O(N__27060),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ));
    LocalMux I__4400 (
            .O(N__27055),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ));
    Odrv4 I__4399 (
            .O(N__27050),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ));
    CascadeMux I__4398 (
            .O(N__27035),
            .I(N__27032));
    InMux I__4397 (
            .O(N__27032),
            .I(N__27029));
    LocalMux I__4396 (
            .O(N__27029),
            .I(N__27026));
    Odrv4 I__4395 (
            .O(N__27026),
            .I(\phase_controller_inst2.stoper_hc.un6_running_15 ));
    CEMux I__4394 (
            .O(N__27023),
            .I(N__27017));
    CEMux I__4393 (
            .O(N__27022),
            .I(N__27010));
    CEMux I__4392 (
            .O(N__27021),
            .I(N__27003));
    CEMux I__4391 (
            .O(N__27020),
            .I(N__27000));
    LocalMux I__4390 (
            .O(N__27017),
            .I(N__26997));
    CEMux I__4389 (
            .O(N__27016),
            .I(N__26994));
    InMux I__4388 (
            .O(N__27015),
            .I(N__26991));
    CEMux I__4387 (
            .O(N__27014),
            .I(N__26988));
    CEMux I__4386 (
            .O(N__27013),
            .I(N__26985));
    LocalMux I__4385 (
            .O(N__27010),
            .I(N__26982));
    InMux I__4384 (
            .O(N__27009),
            .I(N__26973));
    InMux I__4383 (
            .O(N__27008),
            .I(N__26973));
    InMux I__4382 (
            .O(N__27007),
            .I(N__26973));
    InMux I__4381 (
            .O(N__27006),
            .I(N__26973));
    LocalMux I__4380 (
            .O(N__27003),
            .I(N__26970));
    LocalMux I__4379 (
            .O(N__27000),
            .I(N__26967));
    Span4Mux_h I__4378 (
            .O(N__26997),
            .I(N__26950));
    LocalMux I__4377 (
            .O(N__26994),
            .I(N__26947));
    LocalMux I__4376 (
            .O(N__26991),
            .I(N__26942));
    LocalMux I__4375 (
            .O(N__26988),
            .I(N__26942));
    LocalMux I__4374 (
            .O(N__26985),
            .I(N__26939));
    Span4Mux_h I__4373 (
            .O(N__26982),
            .I(N__26936));
    LocalMux I__4372 (
            .O(N__26973),
            .I(N__26929));
    Span4Mux_v I__4371 (
            .O(N__26970),
            .I(N__26929));
    Span4Mux_v I__4370 (
            .O(N__26967),
            .I(N__26929));
    InMux I__4369 (
            .O(N__26966),
            .I(N__26922));
    InMux I__4368 (
            .O(N__26965),
            .I(N__26922));
    InMux I__4367 (
            .O(N__26964),
            .I(N__26922));
    InMux I__4366 (
            .O(N__26963),
            .I(N__26913));
    InMux I__4365 (
            .O(N__26962),
            .I(N__26913));
    InMux I__4364 (
            .O(N__26961),
            .I(N__26913));
    InMux I__4363 (
            .O(N__26960),
            .I(N__26913));
    InMux I__4362 (
            .O(N__26959),
            .I(N__26910));
    InMux I__4361 (
            .O(N__26958),
            .I(N__26905));
    InMux I__4360 (
            .O(N__26957),
            .I(N__26905));
    InMux I__4359 (
            .O(N__26956),
            .I(N__26896));
    InMux I__4358 (
            .O(N__26955),
            .I(N__26896));
    InMux I__4357 (
            .O(N__26954),
            .I(N__26896));
    InMux I__4356 (
            .O(N__26953),
            .I(N__26896));
    Span4Mux_v I__4355 (
            .O(N__26950),
            .I(N__26893));
    Span4Mux_h I__4354 (
            .O(N__26947),
            .I(N__26888));
    Span4Mux_h I__4353 (
            .O(N__26942),
            .I(N__26888));
    Span12Mux_v I__4352 (
            .O(N__26939),
            .I(N__26885));
    Odrv4 I__4351 (
            .O(N__26936),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv4 I__4350 (
            .O(N__26929),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    LocalMux I__4349 (
            .O(N__26922),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    LocalMux I__4348 (
            .O(N__26913),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    LocalMux I__4347 (
            .O(N__26910),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    LocalMux I__4346 (
            .O(N__26905),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    LocalMux I__4345 (
            .O(N__26896),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv4 I__4344 (
            .O(N__26893),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv4 I__4343 (
            .O(N__26888),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv12 I__4342 (
            .O(N__26885),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    InMux I__4341 (
            .O(N__26864),
            .I(N__26861));
    LocalMux I__4340 (
            .O(N__26861),
            .I(N__26857));
    InMux I__4339 (
            .O(N__26860),
            .I(N__26854));
    Span4Mux_h I__4338 (
            .O(N__26857),
            .I(N__26848));
    LocalMux I__4337 (
            .O(N__26854),
            .I(N__26848));
    InMux I__4336 (
            .O(N__26853),
            .I(N__26844));
    Span4Mux_v I__4335 (
            .O(N__26848),
            .I(N__26841));
    InMux I__4334 (
            .O(N__26847),
            .I(N__26838));
    LocalMux I__4333 (
            .O(N__26844),
            .I(elapsed_time_ns_1_RNID6DJ11_0_7));
    Odrv4 I__4332 (
            .O(N__26841),
            .I(elapsed_time_ns_1_RNID6DJ11_0_7));
    LocalMux I__4331 (
            .O(N__26838),
            .I(elapsed_time_ns_1_RNID6DJ11_0_7));
    InMux I__4330 (
            .O(N__26831),
            .I(N__26828));
    LocalMux I__4329 (
            .O(N__26828),
            .I(N__26823));
    InMux I__4328 (
            .O(N__26827),
            .I(N__26820));
    InMux I__4327 (
            .O(N__26826),
            .I(N__26816));
    Span4Mux_h I__4326 (
            .O(N__26823),
            .I(N__26813));
    LocalMux I__4325 (
            .O(N__26820),
            .I(N__26810));
    InMux I__4324 (
            .O(N__26819),
            .I(N__26807));
    LocalMux I__4323 (
            .O(N__26816),
            .I(elapsed_time_ns_1_RNIE7DJ11_0_8));
    Odrv4 I__4322 (
            .O(N__26813),
            .I(elapsed_time_ns_1_RNIE7DJ11_0_8));
    Odrv4 I__4321 (
            .O(N__26810),
            .I(elapsed_time_ns_1_RNIE7DJ11_0_8));
    LocalMux I__4320 (
            .O(N__26807),
            .I(elapsed_time_ns_1_RNIE7DJ11_0_8));
    CascadeMux I__4319 (
            .O(N__26798),
            .I(N__26794));
    CascadeMux I__4318 (
            .O(N__26797),
            .I(N__26791));
    InMux I__4317 (
            .O(N__26794),
            .I(N__26788));
    InMux I__4316 (
            .O(N__26791),
            .I(N__26783));
    LocalMux I__4315 (
            .O(N__26788),
            .I(N__26780));
    InMux I__4314 (
            .O(N__26787),
            .I(N__26777));
    InMux I__4313 (
            .O(N__26786),
            .I(N__26774));
    LocalMux I__4312 (
            .O(N__26783),
            .I(N__26771));
    Span4Mux_h I__4311 (
            .O(N__26780),
            .I(N__26768));
    LocalMux I__4310 (
            .O(N__26777),
            .I(N__26765));
    LocalMux I__4309 (
            .O(N__26774),
            .I(elapsed_time_ns_1_RNIB4DJ11_0_5));
    Odrv4 I__4308 (
            .O(N__26771),
            .I(elapsed_time_ns_1_RNIB4DJ11_0_5));
    Odrv4 I__4307 (
            .O(N__26768),
            .I(elapsed_time_ns_1_RNIB4DJ11_0_5));
    Odrv4 I__4306 (
            .O(N__26765),
            .I(elapsed_time_ns_1_RNIB4DJ11_0_5));
    InMux I__4305 (
            .O(N__26756),
            .I(N__26753));
    LocalMux I__4304 (
            .O(N__26753),
            .I(N__26745));
    InMux I__4303 (
            .O(N__26752),
            .I(N__26742));
    InMux I__4302 (
            .O(N__26751),
            .I(N__26739));
    InMux I__4301 (
            .O(N__26750),
            .I(N__26736));
    InMux I__4300 (
            .O(N__26749),
            .I(N__26731));
    InMux I__4299 (
            .O(N__26748),
            .I(N__26728));
    Span4Mux_v I__4298 (
            .O(N__26745),
            .I(N__26719));
    LocalMux I__4297 (
            .O(N__26742),
            .I(N__26719));
    LocalMux I__4296 (
            .O(N__26739),
            .I(N__26719));
    LocalMux I__4295 (
            .O(N__26736),
            .I(N__26719));
    InMux I__4294 (
            .O(N__26735),
            .I(N__26714));
    InMux I__4293 (
            .O(N__26734),
            .I(N__26714));
    LocalMux I__4292 (
            .O(N__26731),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa ));
    LocalMux I__4291 (
            .O(N__26728),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa ));
    Odrv4 I__4290 (
            .O(N__26719),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa ));
    LocalMux I__4289 (
            .O(N__26714),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa ));
    CascadeMux I__4288 (
            .O(N__26705),
            .I(elapsed_time_ns_1_RNI3VBED1_0_16_cascade_));
    InMux I__4287 (
            .O(N__26702),
            .I(N__26699));
    LocalMux I__4286 (
            .O(N__26699),
            .I(N__26695));
    InMux I__4285 (
            .O(N__26698),
            .I(N__26692));
    Span4Mux_h I__4284 (
            .O(N__26695),
            .I(N__26688));
    LocalMux I__4283 (
            .O(N__26692),
            .I(N__26685));
    InMux I__4282 (
            .O(N__26691),
            .I(N__26682));
    Odrv4 I__4281 (
            .O(N__26688),
            .I(elapsed_time_ns_1_RNIA3DJ11_0_4));
    Odrv4 I__4280 (
            .O(N__26685),
            .I(elapsed_time_ns_1_RNIA3DJ11_0_4));
    LocalMux I__4279 (
            .O(N__26682),
            .I(elapsed_time_ns_1_RNIA3DJ11_0_4));
    InMux I__4278 (
            .O(N__26675),
            .I(N__26668));
    InMux I__4277 (
            .O(N__26674),
            .I(N__26663));
    InMux I__4276 (
            .O(N__26673),
            .I(N__26663));
    InMux I__4275 (
            .O(N__26672),
            .I(N__26658));
    InMux I__4274 (
            .O(N__26671),
            .I(N__26658));
    LocalMux I__4273 (
            .O(N__26668),
            .I(elapsed_time_ns_1_RNI40CED1_0_17));
    LocalMux I__4272 (
            .O(N__26663),
            .I(elapsed_time_ns_1_RNI40CED1_0_17));
    LocalMux I__4271 (
            .O(N__26658),
            .I(elapsed_time_ns_1_RNI40CED1_0_17));
    CascadeMux I__4270 (
            .O(N__26651),
            .I(elapsed_time_ns_1_RNIA3DJ11_0_4_cascade_));
    InMux I__4269 (
            .O(N__26648),
            .I(N__26643));
    InMux I__4268 (
            .O(N__26647),
            .I(N__26640));
    InMux I__4267 (
            .O(N__26646),
            .I(N__26635));
    LocalMux I__4266 (
            .O(N__26643),
            .I(N__26630));
    LocalMux I__4265 (
            .O(N__26640),
            .I(N__26630));
    InMux I__4264 (
            .O(N__26639),
            .I(N__26625));
    InMux I__4263 (
            .O(N__26638),
            .I(N__26625));
    LocalMux I__4262 (
            .O(N__26635),
            .I(elapsed_time_ns_1_RNI51CED1_0_18));
    Odrv12 I__4261 (
            .O(N__26630),
            .I(elapsed_time_ns_1_RNI51CED1_0_18));
    LocalMux I__4260 (
            .O(N__26625),
            .I(elapsed_time_ns_1_RNI51CED1_0_18));
    CascadeMux I__4259 (
            .O(N__26618),
            .I(N__26614));
    InMux I__4258 (
            .O(N__26617),
            .I(N__26609));
    InMux I__4257 (
            .O(N__26614),
            .I(N__26604));
    InMux I__4256 (
            .O(N__26613),
            .I(N__26604));
    InMux I__4255 (
            .O(N__26612),
            .I(N__26601));
    LocalMux I__4254 (
            .O(N__26609),
            .I(elapsed_time_ns_1_RNI62CED1_0_19));
    LocalMux I__4253 (
            .O(N__26604),
            .I(elapsed_time_ns_1_RNI62CED1_0_19));
    LocalMux I__4252 (
            .O(N__26601),
            .I(elapsed_time_ns_1_RNI62CED1_0_19));
    CascadeMux I__4251 (
            .O(N__26594),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2_cascade_ ));
    InMux I__4250 (
            .O(N__26591),
            .I(N__26587));
    InMux I__4249 (
            .O(N__26590),
            .I(N__26584));
    LocalMux I__4248 (
            .O(N__26587),
            .I(N__26579));
    LocalMux I__4247 (
            .O(N__26584),
            .I(N__26579));
    Odrv4 I__4246 (
            .O(N__26579),
            .I(\phase_controller_inst1.stoper_hc.N_328 ));
    CascadeMux I__4245 (
            .O(N__26576),
            .I(N__26571));
    InMux I__4244 (
            .O(N__26575),
            .I(N__26564));
    InMux I__4243 (
            .O(N__26574),
            .I(N__26564));
    InMux I__4242 (
            .O(N__26571),
            .I(N__26564));
    LocalMux I__4241 (
            .O(N__26564),
            .I(\phase_controller_inst1.stoper_hc.N_337 ));
    InMux I__4240 (
            .O(N__26561),
            .I(N__26558));
    LocalMux I__4239 (
            .O(N__26558),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_4 ));
    CascadeMux I__4238 (
            .O(N__26555),
            .I(N__26551));
    InMux I__4237 (
            .O(N__26554),
            .I(N__26547));
    InMux I__4236 (
            .O(N__26551),
            .I(N__26544));
    InMux I__4235 (
            .O(N__26550),
            .I(N__26541));
    LocalMux I__4234 (
            .O(N__26547),
            .I(N__26538));
    LocalMux I__4233 (
            .O(N__26544),
            .I(N__26533));
    LocalMux I__4232 (
            .O(N__26541),
            .I(N__26528));
    Span4Mux_v I__4231 (
            .O(N__26538),
            .I(N__26528));
    InMux I__4230 (
            .O(N__26537),
            .I(N__26523));
    InMux I__4229 (
            .O(N__26536),
            .I(N__26523));
    Odrv4 I__4228 (
            .O(N__26533),
            .I(elapsed_time_ns_1_RNIQURR91_0_3));
    Odrv4 I__4227 (
            .O(N__26528),
            .I(elapsed_time_ns_1_RNIQURR91_0_3));
    LocalMux I__4226 (
            .O(N__26523),
            .I(elapsed_time_ns_1_RNIQURR91_0_3));
    InMux I__4225 (
            .O(N__26516),
            .I(N__26513));
    LocalMux I__4224 (
            .O(N__26513),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3 ));
    CascadeMux I__4223 (
            .O(N__26510),
            .I(N__26507));
    InMux I__4222 (
            .O(N__26507),
            .I(N__26503));
    InMux I__4221 (
            .O(N__26506),
            .I(N__26500));
    LocalMux I__4220 (
            .O(N__26503),
            .I(N__26497));
    LocalMux I__4219 (
            .O(N__26500),
            .I(elapsed_time_ns_1_RNIP2ND11_0_21));
    Odrv12 I__4218 (
            .O(N__26497),
            .I(elapsed_time_ns_1_RNIP2ND11_0_21));
    InMux I__4217 (
            .O(N__26492),
            .I(N__26488));
    InMux I__4216 (
            .O(N__26491),
            .I(N__26485));
    LocalMux I__4215 (
            .O(N__26488),
            .I(elapsed_time_ns_1_RNIS5ND11_0_24));
    LocalMux I__4214 (
            .O(N__26485),
            .I(elapsed_time_ns_1_RNIS5ND11_0_24));
    InMux I__4213 (
            .O(N__26480),
            .I(N__26477));
    LocalMux I__4212 (
            .O(N__26477),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15 ));
    CascadeMux I__4211 (
            .O(N__26474),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15_cascade_ ));
    InMux I__4210 (
            .O(N__26471),
            .I(N__26468));
    LocalMux I__4209 (
            .O(N__26468),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15 ));
    CascadeMux I__4208 (
            .O(N__26465),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15_cascade_ ));
    InMux I__4207 (
            .O(N__26462),
            .I(N__26459));
    LocalMux I__4206 (
            .O(N__26459),
            .I(N__26456));
    Span4Mux_v I__4205 (
            .O(N__26456),
            .I(N__26453));
    Odrv4 I__4204 (
            .O(N__26453),
            .I(\phase_controller_inst2.stoper_hc.un6_running_17 ));
    InMux I__4203 (
            .O(N__26450),
            .I(N__26444));
    InMux I__4202 (
            .O(N__26449),
            .I(N__26444));
    LocalMux I__4201 (
            .O(N__26444),
            .I(elapsed_time_ns_1_RNIQ3ND11_0_22));
    CascadeMux I__4200 (
            .O(N__26441),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17_cascade_ ));
    InMux I__4199 (
            .O(N__26438),
            .I(N__26432));
    InMux I__4198 (
            .O(N__26437),
            .I(N__26432));
    LocalMux I__4197 (
            .O(N__26432),
            .I(elapsed_time_ns_1_RNIR4ND11_0_23));
    InMux I__4196 (
            .O(N__26429),
            .I(N__26426));
    LocalMux I__4195 (
            .O(N__26426),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19 ));
    CascadeMux I__4194 (
            .O(N__26423),
            .I(elapsed_time_ns_1_RNIL13KD1_0_9_cascade_));
    InMux I__4193 (
            .O(N__26420),
            .I(N__26417));
    LocalMux I__4192 (
            .O(N__26417),
            .I(elapsed_time_ns_1_RNI1BND11_0_29));
    CascadeMux I__4191 (
            .O(N__26414),
            .I(elapsed_time_ns_1_RNI1BND11_0_29_cascade_));
    CascadeMux I__4190 (
            .O(N__26411),
            .I(N__26408));
    InMux I__4189 (
            .O(N__26408),
            .I(N__26405));
    LocalMux I__4188 (
            .O(N__26405),
            .I(elapsed_time_ns_1_RNIT6ND11_0_25));
    InMux I__4187 (
            .O(N__26402),
            .I(N__26396));
    InMux I__4186 (
            .O(N__26401),
            .I(N__26396));
    LocalMux I__4185 (
            .O(N__26396),
            .I(elapsed_time_ns_1_RNI0AND11_0_28));
    InMux I__4184 (
            .O(N__26393),
            .I(N__26389));
    InMux I__4183 (
            .O(N__26392),
            .I(N__26386));
    LocalMux I__4182 (
            .O(N__26389),
            .I(elapsed_time_ns_1_RNIV8ND11_0_27));
    LocalMux I__4181 (
            .O(N__26386),
            .I(elapsed_time_ns_1_RNIV8ND11_0_27));
    CascadeMux I__4180 (
            .O(N__26381),
            .I(elapsed_time_ns_1_RNIT6ND11_0_25_cascade_));
    InMux I__4179 (
            .O(N__26378),
            .I(N__26374));
    InMux I__4178 (
            .O(N__26377),
            .I(N__26371));
    LocalMux I__4177 (
            .O(N__26374),
            .I(elapsed_time_ns_1_RNIU7ND11_0_26));
    LocalMux I__4176 (
            .O(N__26371),
            .I(elapsed_time_ns_1_RNIU7ND11_0_26));
    InMux I__4175 (
            .O(N__26366),
            .I(N__26360));
    InMux I__4174 (
            .O(N__26365),
            .I(N__26352));
    InMux I__4173 (
            .O(N__26364),
            .I(N__26352));
    InMux I__4172 (
            .O(N__26363),
            .I(N__26352));
    LocalMux I__4171 (
            .O(N__26360),
            .I(N__26349));
    InMux I__4170 (
            .O(N__26359),
            .I(N__26346));
    LocalMux I__4169 (
            .O(N__26352),
            .I(N__26343));
    Span4Mux_v I__4168 (
            .O(N__26349),
            .I(N__26340));
    LocalMux I__4167 (
            .O(N__26346),
            .I(N__26337));
    Span4Mux_h I__4166 (
            .O(N__26343),
            .I(N__26334));
    Odrv4 I__4165 (
            .O(N__26340),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv12 I__4164 (
            .O(N__26337),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__4163 (
            .O(N__26334),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    CascadeMux I__4162 (
            .O(N__26327),
            .I(N__26324));
    InMux I__4161 (
            .O(N__26324),
            .I(N__26321));
    LocalMux I__4160 (
            .O(N__26321),
            .I(N__26318));
    Odrv4 I__4159 (
            .O(N__26318),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0 ));
    CascadeMux I__4158 (
            .O(N__26315),
            .I(N__26312));
    InMux I__4157 (
            .O(N__26312),
            .I(N__26309));
    LocalMux I__4156 (
            .O(N__26309),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0 ));
    CascadeMux I__4155 (
            .O(N__26306),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5_cascade_ ));
    CascadeMux I__4154 (
            .O(N__26303),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14_cascade_ ));
    InMux I__4153 (
            .O(N__26300),
            .I(N__26295));
    InMux I__4152 (
            .O(N__26299),
            .I(N__26292));
    InMux I__4151 (
            .O(N__26298),
            .I(N__26289));
    LocalMux I__4150 (
            .O(N__26295),
            .I(N__26286));
    LocalMux I__4149 (
            .O(N__26292),
            .I(N__26283));
    LocalMux I__4148 (
            .O(N__26289),
            .I(N__26280));
    Span4Mux_h I__4147 (
            .O(N__26286),
            .I(N__26275));
    Span4Mux_h I__4146 (
            .O(N__26283),
            .I(N__26270));
    Span4Mux_h I__4145 (
            .O(N__26280),
            .I(N__26270));
    InMux I__4144 (
            .O(N__26279),
            .I(N__26265));
    InMux I__4143 (
            .O(N__26278),
            .I(N__26265));
    Odrv4 I__4142 (
            .O(N__26275),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__4141 (
            .O(N__26270),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    LocalMux I__4140 (
            .O(N__26265),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    InMux I__4139 (
            .O(N__26258),
            .I(N__26255));
    LocalMux I__4138 (
            .O(N__26255),
            .I(N__26252));
    Odrv4 I__4137 (
            .O(N__26252),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0 ));
    CascadeMux I__4136 (
            .O(N__26249),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23_cascade_ ));
    CascadeMux I__4135 (
            .O(N__26246),
            .I(N__26243));
    InMux I__4134 (
            .O(N__26243),
            .I(N__26240));
    LocalMux I__4133 (
            .O(N__26240),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0 ));
    CascadeMux I__4132 (
            .O(N__26237),
            .I(N__26233));
    InMux I__4131 (
            .O(N__26236),
            .I(N__26230));
    InMux I__4130 (
            .O(N__26233),
            .I(N__26227));
    LocalMux I__4129 (
            .O(N__26230),
            .I(N__26222));
    LocalMux I__4128 (
            .O(N__26227),
            .I(N__26219));
    InMux I__4127 (
            .O(N__26226),
            .I(N__26216));
    InMux I__4126 (
            .O(N__26225),
            .I(N__26212));
    Span4Mux_h I__4125 (
            .O(N__26222),
            .I(N__26207));
    Span4Mux_h I__4124 (
            .O(N__26219),
            .I(N__26207));
    LocalMux I__4123 (
            .O(N__26216),
            .I(N__26204));
    InMux I__4122 (
            .O(N__26215),
            .I(N__26201));
    LocalMux I__4121 (
            .O(N__26212),
            .I(N__26198));
    Odrv4 I__4120 (
            .O(N__26207),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__4119 (
            .O(N__26204),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    LocalMux I__4118 (
            .O(N__26201),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__4117 (
            .O(N__26198),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    CascadeMux I__4116 (
            .O(N__26189),
            .I(N__26186));
    InMux I__4115 (
            .O(N__26186),
            .I(N__26183));
    LocalMux I__4114 (
            .O(N__26183),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0 ));
    CascadeMux I__4113 (
            .O(N__26180),
            .I(N__26177));
    InMux I__4112 (
            .O(N__26177),
            .I(N__26172));
    InMux I__4111 (
            .O(N__26176),
            .I(N__26169));
    InMux I__4110 (
            .O(N__26175),
            .I(N__26166));
    LocalMux I__4109 (
            .O(N__26172),
            .I(N__26162));
    LocalMux I__4108 (
            .O(N__26169),
            .I(N__26159));
    LocalMux I__4107 (
            .O(N__26166),
            .I(N__26156));
    InMux I__4106 (
            .O(N__26165),
            .I(N__26153));
    Span4Mux_h I__4105 (
            .O(N__26162),
            .I(N__26150));
    Span4Mux_v I__4104 (
            .O(N__26159),
            .I(N__26145));
    Span4Mux_v I__4103 (
            .O(N__26156),
            .I(N__26145));
    LocalMux I__4102 (
            .O(N__26153),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    Odrv4 I__4101 (
            .O(N__26150),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    Odrv4 I__4100 (
            .O(N__26145),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    InMux I__4099 (
            .O(N__26138),
            .I(N__26135));
    LocalMux I__4098 (
            .O(N__26135),
            .I(N__26132));
    Span4Mux_h I__4097 (
            .O(N__26132),
            .I(N__26129));
    Odrv4 I__4096 (
            .O(N__26129),
            .I(\current_shift_inst.PI_CTRL.integrator_i_2 ));
    CascadeMux I__4095 (
            .O(N__26126),
            .I(N__26122));
    InMux I__4094 (
            .O(N__26125),
            .I(N__26118));
    InMux I__4093 (
            .O(N__26122),
            .I(N__26115));
    InMux I__4092 (
            .O(N__26121),
            .I(N__26112));
    LocalMux I__4091 (
            .O(N__26118),
            .I(N__26109));
    LocalMux I__4090 (
            .O(N__26115),
            .I(N__26106));
    LocalMux I__4089 (
            .O(N__26112),
            .I(N__26103));
    Span4Mux_h I__4088 (
            .O(N__26109),
            .I(N__26096));
    Span4Mux_h I__4087 (
            .O(N__26106),
            .I(N__26096));
    Span4Mux_h I__4086 (
            .O(N__26103),
            .I(N__26093));
    InMux I__4085 (
            .O(N__26102),
            .I(N__26088));
    InMux I__4084 (
            .O(N__26101),
            .I(N__26088));
    Odrv4 I__4083 (
            .O(N__26096),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__4082 (
            .O(N__26093),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    LocalMux I__4081 (
            .O(N__26088),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    CascadeMux I__4080 (
            .O(N__26081),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30_cascade_ ));
    InMux I__4079 (
            .O(N__26078),
            .I(N__26075));
    LocalMux I__4078 (
            .O(N__26075),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0 ));
    CascadeMux I__4077 (
            .O(N__26072),
            .I(N__26068));
    InMux I__4076 (
            .O(N__26071),
            .I(N__26065));
    InMux I__4075 (
            .O(N__26068),
            .I(N__26062));
    LocalMux I__4074 (
            .O(N__26065),
            .I(N__26058));
    LocalMux I__4073 (
            .O(N__26062),
            .I(N__26055));
    InMux I__4072 (
            .O(N__26061),
            .I(N__26050));
    Span4Mux_v I__4071 (
            .O(N__26058),
            .I(N__26045));
    Span4Mux_v I__4070 (
            .O(N__26055),
            .I(N__26045));
    InMux I__4069 (
            .O(N__26054),
            .I(N__26042));
    InMux I__4068 (
            .O(N__26053),
            .I(N__26039));
    LocalMux I__4067 (
            .O(N__26050),
            .I(N__26036));
    Odrv4 I__4066 (
            .O(N__26045),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    LocalMux I__4065 (
            .O(N__26042),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    LocalMux I__4064 (
            .O(N__26039),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__4063 (
            .O(N__26036),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    CascadeMux I__4062 (
            .O(N__26027),
            .I(N__26024));
    InMux I__4061 (
            .O(N__26024),
            .I(N__26021));
    LocalMux I__4060 (
            .O(N__26021),
            .I(N__26018));
    Odrv4 I__4059 (
            .O(N__26018),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0 ));
    CascadeMux I__4058 (
            .O(N__26015),
            .I(N__26010));
    CascadeMux I__4057 (
            .O(N__26014),
            .I(N__26007));
    InMux I__4056 (
            .O(N__26013),
            .I(N__26002));
    InMux I__4055 (
            .O(N__26010),
            .I(N__25999));
    InMux I__4054 (
            .O(N__26007),
            .I(N__25994));
    InMux I__4053 (
            .O(N__26006),
            .I(N__25994));
    InMux I__4052 (
            .O(N__26005),
            .I(N__25991));
    LocalMux I__4051 (
            .O(N__26002),
            .I(N__25988));
    LocalMux I__4050 (
            .O(N__25999),
            .I(N__25985));
    LocalMux I__4049 (
            .O(N__25994),
            .I(N__25980));
    LocalMux I__4048 (
            .O(N__25991),
            .I(N__25980));
    Span4Mux_h I__4047 (
            .O(N__25988),
            .I(N__25973));
    Span4Mux_h I__4046 (
            .O(N__25985),
            .I(N__25973));
    Span4Mux_v I__4045 (
            .O(N__25980),
            .I(N__25973));
    Odrv4 I__4044 (
            .O(N__25973),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    CascadeMux I__4043 (
            .O(N__25970),
            .I(N__25967));
    InMux I__4042 (
            .O(N__25967),
            .I(N__25964));
    LocalMux I__4041 (
            .O(N__25964),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0 ));
    CascadeMux I__4040 (
            .O(N__25961),
            .I(N__25958));
    InMux I__4039 (
            .O(N__25958),
            .I(N__25955));
    LocalMux I__4038 (
            .O(N__25955),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0 ));
    InMux I__4037 (
            .O(N__25952),
            .I(N__25949));
    LocalMux I__4036 (
            .O(N__25949),
            .I(N__25945));
    InMux I__4035 (
            .O(N__25948),
            .I(N__25942));
    Span4Mux_h I__4034 (
            .O(N__25945),
            .I(N__25937));
    LocalMux I__4033 (
            .O(N__25942),
            .I(N__25937));
    Span4Mux_h I__4032 (
            .O(N__25937),
            .I(N__25931));
    InMux I__4031 (
            .O(N__25936),
            .I(N__25928));
    InMux I__4030 (
            .O(N__25935),
            .I(N__25923));
    InMux I__4029 (
            .O(N__25934),
            .I(N__25923));
    Odrv4 I__4028 (
            .O(N__25931),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    LocalMux I__4027 (
            .O(N__25928),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    LocalMux I__4026 (
            .O(N__25923),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    CascadeMux I__4025 (
            .O(N__25916),
            .I(N__25913));
    InMux I__4024 (
            .O(N__25913),
            .I(N__25910));
    LocalMux I__4023 (
            .O(N__25910),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0 ));
    CascadeMux I__4022 (
            .O(N__25907),
            .I(N__25903));
    InMux I__4021 (
            .O(N__25906),
            .I(N__25900));
    InMux I__4020 (
            .O(N__25903),
            .I(N__25897));
    LocalMux I__4019 (
            .O(N__25900),
            .I(N__25894));
    LocalMux I__4018 (
            .O(N__25897),
            .I(N__25891));
    Span4Mux_h I__4017 (
            .O(N__25894),
            .I(N__25883));
    Span4Mux_h I__4016 (
            .O(N__25891),
            .I(N__25883));
    InMux I__4015 (
            .O(N__25890),
            .I(N__25880));
    InMux I__4014 (
            .O(N__25889),
            .I(N__25877));
    InMux I__4013 (
            .O(N__25888),
            .I(N__25874));
    Odrv4 I__4012 (
            .O(N__25883),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__4011 (
            .O(N__25880),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__4010 (
            .O(N__25877),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__4009 (
            .O(N__25874),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    CascadeMux I__4008 (
            .O(N__25865),
            .I(N__25862));
    InMux I__4007 (
            .O(N__25862),
            .I(N__25859));
    LocalMux I__4006 (
            .O(N__25859),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0 ));
    InMux I__4005 (
            .O(N__25856),
            .I(N__25852));
    InMux I__4004 (
            .O(N__25855),
            .I(N__25849));
    LocalMux I__4003 (
            .O(N__25852),
            .I(N__25846));
    LocalMux I__4002 (
            .O(N__25849),
            .I(N__25843));
    Span4Mux_h I__4001 (
            .O(N__25846),
            .I(N__25835));
    Span4Mux_h I__4000 (
            .O(N__25843),
            .I(N__25835));
    InMux I__3999 (
            .O(N__25842),
            .I(N__25832));
    InMux I__3998 (
            .O(N__25841),
            .I(N__25829));
    InMux I__3997 (
            .O(N__25840),
            .I(N__25826));
    Odrv4 I__3996 (
            .O(N__25835),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    LocalMux I__3995 (
            .O(N__25832),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    LocalMux I__3994 (
            .O(N__25829),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    LocalMux I__3993 (
            .O(N__25826),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    CascadeMux I__3992 (
            .O(N__25817),
            .I(N__25814));
    InMux I__3991 (
            .O(N__25814),
            .I(N__25811));
    LocalMux I__3990 (
            .O(N__25811),
            .I(N__25808));
    Odrv4 I__3989 (
            .O(N__25808),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0 ));
    CascadeMux I__3988 (
            .O(N__25805),
            .I(N__25802));
    InMux I__3987 (
            .O(N__25802),
            .I(N__25799));
    LocalMux I__3986 (
            .O(N__25799),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0 ));
    InMux I__3985 (
            .O(N__25796),
            .I(N__25792));
    InMux I__3984 (
            .O(N__25795),
            .I(N__25789));
    LocalMux I__3983 (
            .O(N__25792),
            .I(N__25786));
    LocalMux I__3982 (
            .O(N__25789),
            .I(N__25782));
    Span4Mux_v I__3981 (
            .O(N__25786),
            .I(N__25779));
    InMux I__3980 (
            .O(N__25785),
            .I(N__25776));
    Span4Mux_h I__3979 (
            .O(N__25782),
            .I(N__25769));
    Span4Mux_h I__3978 (
            .O(N__25779),
            .I(N__25769));
    LocalMux I__3977 (
            .O(N__25776),
            .I(N__25766));
    InMux I__3976 (
            .O(N__25775),
            .I(N__25761));
    InMux I__3975 (
            .O(N__25774),
            .I(N__25761));
    Odrv4 I__3974 (
            .O(N__25769),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__3973 (
            .O(N__25766),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    LocalMux I__3972 (
            .O(N__25761),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    InMux I__3971 (
            .O(N__25754),
            .I(N__25751));
    LocalMux I__3970 (
            .O(N__25751),
            .I(N__25747));
    InMux I__3969 (
            .O(N__25750),
            .I(N__25743));
    Span4Mux_v I__3968 (
            .O(N__25747),
            .I(N__25740));
    InMux I__3967 (
            .O(N__25746),
            .I(N__25737));
    LocalMux I__3966 (
            .O(N__25743),
            .I(N__25732));
    Span4Mux_h I__3965 (
            .O(N__25740),
            .I(N__25727));
    LocalMux I__3964 (
            .O(N__25737),
            .I(N__25727));
    InMux I__3963 (
            .O(N__25736),
            .I(N__25722));
    InMux I__3962 (
            .O(N__25735),
            .I(N__25722));
    Odrv4 I__3961 (
            .O(N__25732),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv4 I__3960 (
            .O(N__25727),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    LocalMux I__3959 (
            .O(N__25722),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    CascadeMux I__3958 (
            .O(N__25715),
            .I(N__25710));
    CascadeMux I__3957 (
            .O(N__25714),
            .I(N__25707));
    InMux I__3956 (
            .O(N__25713),
            .I(N__25704));
    InMux I__3955 (
            .O(N__25710),
            .I(N__25701));
    InMux I__3954 (
            .O(N__25707),
            .I(N__25698));
    LocalMux I__3953 (
            .O(N__25704),
            .I(N__25694));
    LocalMux I__3952 (
            .O(N__25701),
            .I(N__25691));
    LocalMux I__3951 (
            .O(N__25698),
            .I(N__25688));
    InMux I__3950 (
            .O(N__25697),
            .I(N__25684));
    Span4Mux_v I__3949 (
            .O(N__25694),
            .I(N__25681));
    Span4Mux_v I__3948 (
            .O(N__25691),
            .I(N__25676));
    Span4Mux_v I__3947 (
            .O(N__25688),
            .I(N__25676));
    InMux I__3946 (
            .O(N__25687),
            .I(N__25673));
    LocalMux I__3945 (
            .O(N__25684),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv4 I__3944 (
            .O(N__25681),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv4 I__3943 (
            .O(N__25676),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    LocalMux I__3942 (
            .O(N__25673),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    InMux I__3941 (
            .O(N__25664),
            .I(N__25661));
    LocalMux I__3940 (
            .O(N__25661),
            .I(N__25658));
    Odrv4 I__3939 (
            .O(N__25658),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3 ));
    InMux I__3938 (
            .O(N__25655),
            .I(N__25651));
    InMux I__3937 (
            .O(N__25654),
            .I(N__25648));
    LocalMux I__3936 (
            .O(N__25651),
            .I(N__25645));
    LocalMux I__3935 (
            .O(N__25648),
            .I(N__25642));
    Span4Mux_v I__3934 (
            .O(N__25645),
            .I(N__25639));
    Span4Mux_h I__3933 (
            .O(N__25642),
            .I(N__25636));
    Span4Mux_h I__3932 (
            .O(N__25639),
            .I(N__25633));
    Odrv4 I__3931 (
            .O(N__25636),
            .I(\current_shift_inst.PI_CTRL.N_72 ));
    Odrv4 I__3930 (
            .O(N__25633),
            .I(\current_shift_inst.PI_CTRL.N_72 ));
    CascadeMux I__3929 (
            .O(N__25628),
            .I(N__25625));
    InMux I__3928 (
            .O(N__25625),
            .I(N__25622));
    LocalMux I__3927 (
            .O(N__25622),
            .I(N__25619));
    Odrv4 I__3926 (
            .O(N__25619),
            .I(\current_shift_inst.PI_CTRL.integrator_i_25 ));
    InMux I__3925 (
            .O(N__25616),
            .I(N__25612));
    InMux I__3924 (
            .O(N__25615),
            .I(N__25609));
    LocalMux I__3923 (
            .O(N__25612),
            .I(N__25606));
    LocalMux I__3922 (
            .O(N__25609),
            .I(N__25603));
    Span4Mux_v I__3921 (
            .O(N__25606),
            .I(N__25600));
    Span4Mux_h I__3920 (
            .O(N__25603),
            .I(N__25597));
    Odrv4 I__3919 (
            .O(N__25600),
            .I(\current_shift_inst.PI_CTRL.integrator_i_0 ));
    Odrv4 I__3918 (
            .O(N__25597),
            .I(\current_shift_inst.PI_CTRL.integrator_i_0 ));
    CascadeMux I__3917 (
            .O(N__25592),
            .I(N__25589));
    InMux I__3916 (
            .O(N__25589),
            .I(N__25586));
    LocalMux I__3915 (
            .O(N__25586),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4 ));
    CascadeMux I__3914 (
            .O(N__25583),
            .I(N__25580));
    InMux I__3913 (
            .O(N__25580),
            .I(N__25577));
    LocalMux I__3912 (
            .O(N__25577),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0 ));
    CascadeMux I__3911 (
            .O(N__25574),
            .I(N__25571));
    InMux I__3910 (
            .O(N__25571),
            .I(N__25568));
    LocalMux I__3909 (
            .O(N__25568),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6 ));
    CascadeMux I__3908 (
            .O(N__25565),
            .I(N__25562));
    InMux I__3907 (
            .O(N__25562),
            .I(N__25559));
    LocalMux I__3906 (
            .O(N__25559),
            .I(N__25555));
    InMux I__3905 (
            .O(N__25558),
            .I(N__25552));
    Span4Mux_h I__3904 (
            .O(N__25555),
            .I(N__25549));
    LocalMux I__3903 (
            .O(N__25552),
            .I(N__25541));
    Span4Mux_h I__3902 (
            .O(N__25549),
            .I(N__25541));
    InMux I__3901 (
            .O(N__25548),
            .I(N__25536));
    InMux I__3900 (
            .O(N__25547),
            .I(N__25536));
    InMux I__3899 (
            .O(N__25546),
            .I(N__25533));
    Odrv4 I__3898 (
            .O(N__25541),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    LocalMux I__3897 (
            .O(N__25536),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    LocalMux I__3896 (
            .O(N__25533),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    CascadeMux I__3895 (
            .O(N__25526),
            .I(N__25523));
    InMux I__3894 (
            .O(N__25523),
            .I(N__25520));
    LocalMux I__3893 (
            .O(N__25520),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0 ));
    InMux I__3892 (
            .O(N__25517),
            .I(N__25514));
    LocalMux I__3891 (
            .O(N__25514),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0 ));
    CascadeMux I__3890 (
            .O(N__25511),
            .I(N__25506));
    CascadeMux I__3889 (
            .O(N__25510),
            .I(N__25502));
    InMux I__3888 (
            .O(N__25509),
            .I(N__25497));
    InMux I__3887 (
            .O(N__25506),
            .I(N__25497));
    InMux I__3886 (
            .O(N__25505),
            .I(N__25494));
    InMux I__3885 (
            .O(N__25502),
            .I(N__25491));
    LocalMux I__3884 (
            .O(N__25497),
            .I(N__25486));
    LocalMux I__3883 (
            .O(N__25494),
            .I(N__25481));
    LocalMux I__3882 (
            .O(N__25491),
            .I(N__25481));
    InMux I__3881 (
            .O(N__25490),
            .I(N__25476));
    InMux I__3880 (
            .O(N__25489),
            .I(N__25476));
    Odrv4 I__3879 (
            .O(N__25486),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv12 I__3878 (
            .O(N__25481),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    LocalMux I__3877 (
            .O(N__25476),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    CascadeMux I__3876 (
            .O(N__25469),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15_cascade_ ));
    CascadeMux I__3875 (
            .O(N__25466),
            .I(N__25463));
    InMux I__3874 (
            .O(N__25463),
            .I(N__25460));
    LocalMux I__3873 (
            .O(N__25460),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0 ));
    CascadeMux I__3872 (
            .O(N__25457),
            .I(N__25454));
    InMux I__3871 (
            .O(N__25454),
            .I(N__25451));
    LocalMux I__3870 (
            .O(N__25451),
            .I(N__25448));
    Odrv4 I__3869 (
            .O(N__25448),
            .I(\current_shift_inst.PI_CTRL.integrator_i_4 ));
    InMux I__3868 (
            .O(N__25445),
            .I(N__25442));
    LocalMux I__3867 (
            .O(N__25442),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    CascadeMux I__3866 (
            .O(N__25439),
            .I(N__25436));
    InMux I__3865 (
            .O(N__25436),
            .I(N__25433));
    LocalMux I__3864 (
            .O(N__25433),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    InMux I__3863 (
            .O(N__25430),
            .I(N__25427));
    LocalMux I__3862 (
            .O(N__25427),
            .I(N__25424));
    Odrv4 I__3861 (
            .O(N__25424),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    InMux I__3860 (
            .O(N__25421),
            .I(N__25418));
    LocalMux I__3859 (
            .O(N__25418),
            .I(N__25415));
    Odrv4 I__3858 (
            .O(N__25415),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ));
    InMux I__3857 (
            .O(N__25412),
            .I(N__25409));
    LocalMux I__3856 (
            .O(N__25409),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    CascadeMux I__3855 (
            .O(N__25406),
            .I(N__25403));
    InMux I__3854 (
            .O(N__25403),
            .I(N__25400));
    LocalMux I__3853 (
            .O(N__25400),
            .I(N__25397));
    Odrv12 I__3852 (
            .O(N__25397),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ));
    CascadeMux I__3851 (
            .O(N__25394),
            .I(N__25391));
    InMux I__3850 (
            .O(N__25391),
            .I(N__25388));
    LocalMux I__3849 (
            .O(N__25388),
            .I(N__25385));
    Odrv4 I__3848 (
            .O(N__25385),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7 ));
    InMux I__3847 (
            .O(N__25382),
            .I(N__25375));
    CascadeMux I__3846 (
            .O(N__25381),
            .I(N__25372));
    InMux I__3845 (
            .O(N__25380),
            .I(N__25367));
    InMux I__3844 (
            .O(N__25379),
            .I(N__25367));
    InMux I__3843 (
            .O(N__25378),
            .I(N__25364));
    LocalMux I__3842 (
            .O(N__25375),
            .I(N__25361));
    InMux I__3841 (
            .O(N__25372),
            .I(N__25358));
    LocalMux I__3840 (
            .O(N__25367),
            .I(N__25355));
    LocalMux I__3839 (
            .O(N__25364),
            .I(N__25352));
    Span4Mux_v I__3838 (
            .O(N__25361),
            .I(N__25349));
    LocalMux I__3837 (
            .O(N__25358),
            .I(N__25346));
    Span4Mux_h I__3836 (
            .O(N__25355),
            .I(N__25341));
    Span4Mux_h I__3835 (
            .O(N__25352),
            .I(N__25341));
    Odrv4 I__3834 (
            .O(N__25349),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv4 I__3833 (
            .O(N__25346),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv4 I__3832 (
            .O(N__25341),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    CascadeMux I__3831 (
            .O(N__25334),
            .I(N__25331));
    InMux I__3830 (
            .O(N__25331),
            .I(N__25328));
    LocalMux I__3829 (
            .O(N__25328),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0 ));
    InMux I__3828 (
            .O(N__25325),
            .I(N__25321));
    InMux I__3827 (
            .O(N__25324),
            .I(N__25318));
    LocalMux I__3826 (
            .O(N__25321),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__3825 (
            .O(N__25318),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__3824 (
            .O(N__25313),
            .I(N__25310));
    LocalMux I__3823 (
            .O(N__25310),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ));
    InMux I__3822 (
            .O(N__25307),
            .I(N__25304));
    LocalMux I__3821 (
            .O(N__25304),
            .I(N__25301));
    Odrv4 I__3820 (
            .O(N__25301),
            .I(\phase_controller_inst2.stoper_hc.un6_running_16 ));
    InMux I__3819 (
            .O(N__25298),
            .I(N__25294));
    InMux I__3818 (
            .O(N__25297),
            .I(N__25291));
    LocalMux I__3817 (
            .O(N__25294),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    LocalMux I__3816 (
            .O(N__25291),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    CascadeMux I__3815 (
            .O(N__25286),
            .I(N__25283));
    InMux I__3814 (
            .O(N__25283),
            .I(N__25280));
    LocalMux I__3813 (
            .O(N__25280),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_16 ));
    InMux I__3812 (
            .O(N__25277),
            .I(N__25273));
    InMux I__3811 (
            .O(N__25276),
            .I(N__25270));
    LocalMux I__3810 (
            .O(N__25273),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    LocalMux I__3809 (
            .O(N__25270),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    CascadeMux I__3808 (
            .O(N__25265),
            .I(N__25262));
    InMux I__3807 (
            .O(N__25262),
            .I(N__25259));
    LocalMux I__3806 (
            .O(N__25259),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_17 ));
    InMux I__3805 (
            .O(N__25256),
            .I(N__25253));
    LocalMux I__3804 (
            .O(N__25253),
            .I(N__25250));
    Span4Mux_v I__3803 (
            .O(N__25250),
            .I(N__25247));
    Odrv4 I__3802 (
            .O(N__25247),
            .I(\phase_controller_inst2.stoper_hc.un6_running_18 ));
    InMux I__3801 (
            .O(N__25244),
            .I(N__25240));
    InMux I__3800 (
            .O(N__25243),
            .I(N__25237));
    LocalMux I__3799 (
            .O(N__25240),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__3798 (
            .O(N__25237),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    CascadeMux I__3797 (
            .O(N__25232),
            .I(N__25229));
    InMux I__3796 (
            .O(N__25229),
            .I(N__25226));
    LocalMux I__3795 (
            .O(N__25226),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_18 ));
    InMux I__3794 (
            .O(N__25223),
            .I(N__25219));
    InMux I__3793 (
            .O(N__25222),
            .I(N__25216));
    LocalMux I__3792 (
            .O(N__25219),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__3791 (
            .O(N__25216),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    CascadeMux I__3790 (
            .O(N__25211),
            .I(N__25208));
    InMux I__3789 (
            .O(N__25208),
            .I(N__25205));
    LocalMux I__3788 (
            .O(N__25205),
            .I(N__25202));
    Odrv12 I__3787 (
            .O(N__25202),
            .I(\phase_controller_inst2.stoper_hc.un6_running_19 ));
    InMux I__3786 (
            .O(N__25199),
            .I(N__25196));
    LocalMux I__3785 (
            .O(N__25196),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_19 ));
    InMux I__3784 (
            .O(N__25193),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_19 ));
    IoInMux I__3783 (
            .O(N__25190),
            .I(N__25187));
    LocalMux I__3782 (
            .O(N__25187),
            .I(N__25184));
    Span12Mux_s1_v I__3781 (
            .O(N__25184),
            .I(N__25181));
    Odrv12 I__3780 (
            .O(N__25181),
            .I(s3_phy_c));
    InMux I__3779 (
            .O(N__25178),
            .I(N__25175));
    LocalMux I__3778 (
            .O(N__25175),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8 ));
    CascadeMux I__3777 (
            .O(N__25172),
            .I(N__25169));
    InMux I__3776 (
            .O(N__25169),
            .I(N__25166));
    LocalMux I__3775 (
            .O(N__25166),
            .I(N__25163));
    Odrv4 I__3774 (
            .O(N__25163),
            .I(\phase_controller_inst2.stoper_hc.un6_running_8 ));
    InMux I__3773 (
            .O(N__25160),
            .I(N__25156));
    InMux I__3772 (
            .O(N__25159),
            .I(N__25153));
    LocalMux I__3771 (
            .O(N__25156),
            .I(N__25150));
    LocalMux I__3770 (
            .O(N__25153),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    Odrv4 I__3769 (
            .O(N__25150),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__3768 (
            .O(N__25145),
            .I(N__25142));
    LocalMux I__3767 (
            .O(N__25142),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ));
    CascadeMux I__3766 (
            .O(N__25139),
            .I(N__25136));
    InMux I__3765 (
            .O(N__25136),
            .I(N__25133));
    LocalMux I__3764 (
            .O(N__25133),
            .I(N__25130));
    Odrv12 I__3763 (
            .O(N__25130),
            .I(\phase_controller_inst2.stoper_hc.un6_running_9 ));
    InMux I__3762 (
            .O(N__25127),
            .I(N__25123));
    InMux I__3761 (
            .O(N__25126),
            .I(N__25120));
    LocalMux I__3760 (
            .O(N__25123),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__3759 (
            .O(N__25120),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__3758 (
            .O(N__25115),
            .I(N__25112));
    LocalMux I__3757 (
            .O(N__25112),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ));
    InMux I__3756 (
            .O(N__25109),
            .I(N__25106));
    LocalMux I__3755 (
            .O(N__25106),
            .I(N__25103));
    Odrv12 I__3754 (
            .O(N__25103),
            .I(\phase_controller_inst2.stoper_hc.un6_running_10 ));
    InMux I__3753 (
            .O(N__25100),
            .I(N__25096));
    InMux I__3752 (
            .O(N__25099),
            .I(N__25093));
    LocalMux I__3751 (
            .O(N__25096),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__3750 (
            .O(N__25093),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    CascadeMux I__3749 (
            .O(N__25088),
            .I(N__25085));
    InMux I__3748 (
            .O(N__25085),
            .I(N__25082));
    LocalMux I__3747 (
            .O(N__25082),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ));
    InMux I__3746 (
            .O(N__25079),
            .I(N__25076));
    LocalMux I__3745 (
            .O(N__25076),
            .I(N__25073));
    Span4Mux_v I__3744 (
            .O(N__25073),
            .I(N__25070));
    Odrv4 I__3743 (
            .O(N__25070),
            .I(\phase_controller_inst2.stoper_hc.un6_running_11 ));
    InMux I__3742 (
            .O(N__25067),
            .I(N__25063));
    InMux I__3741 (
            .O(N__25066),
            .I(N__25060));
    LocalMux I__3740 (
            .O(N__25063),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__3739 (
            .O(N__25060),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    CascadeMux I__3738 (
            .O(N__25055),
            .I(N__25052));
    InMux I__3737 (
            .O(N__25052),
            .I(N__25049));
    LocalMux I__3736 (
            .O(N__25049),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ));
    CascadeMux I__3735 (
            .O(N__25046),
            .I(N__25043));
    InMux I__3734 (
            .O(N__25043),
            .I(N__25040));
    LocalMux I__3733 (
            .O(N__25040),
            .I(N__25037));
    Odrv12 I__3732 (
            .O(N__25037),
            .I(\phase_controller_inst2.stoper_hc.un6_running_12 ));
    InMux I__3731 (
            .O(N__25034),
            .I(N__25030));
    InMux I__3730 (
            .O(N__25033),
            .I(N__25027));
    LocalMux I__3729 (
            .O(N__25030),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    LocalMux I__3728 (
            .O(N__25027),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__3727 (
            .O(N__25022),
            .I(N__25019));
    LocalMux I__3726 (
            .O(N__25019),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ));
    InMux I__3725 (
            .O(N__25016),
            .I(N__25013));
    LocalMux I__3724 (
            .O(N__25013),
            .I(N__25010));
    Odrv12 I__3723 (
            .O(N__25010),
            .I(\phase_controller_inst2.stoper_hc.un6_running_13 ));
    InMux I__3722 (
            .O(N__25007),
            .I(N__25003));
    InMux I__3721 (
            .O(N__25006),
            .I(N__25000));
    LocalMux I__3720 (
            .O(N__25003),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    LocalMux I__3719 (
            .O(N__25000),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    CascadeMux I__3718 (
            .O(N__24995),
            .I(N__24992));
    InMux I__3717 (
            .O(N__24992),
            .I(N__24989));
    LocalMux I__3716 (
            .O(N__24989),
            .I(N__24986));
    Odrv4 I__3715 (
            .O(N__24986),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ));
    InMux I__3714 (
            .O(N__24983),
            .I(N__24980));
    LocalMux I__3713 (
            .O(N__24980),
            .I(N__24977));
    Odrv12 I__3712 (
            .O(N__24977),
            .I(\phase_controller_inst2.stoper_hc.un6_running_14 ));
    InMux I__3711 (
            .O(N__24974),
            .I(N__24970));
    InMux I__3710 (
            .O(N__24973),
            .I(N__24967));
    LocalMux I__3709 (
            .O(N__24970),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__3708 (
            .O(N__24967),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    CascadeMux I__3707 (
            .O(N__24962),
            .I(N__24959));
    InMux I__3706 (
            .O(N__24959),
            .I(N__24956));
    LocalMux I__3705 (
            .O(N__24956),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ));
    CascadeMux I__3704 (
            .O(N__24953),
            .I(N__24946));
    CascadeMux I__3703 (
            .O(N__24952),
            .I(N__24935));
    CascadeMux I__3702 (
            .O(N__24951),
            .I(N__24932));
    CascadeMux I__3701 (
            .O(N__24950),
            .I(N__24929));
    CascadeMux I__3700 (
            .O(N__24949),
            .I(N__24926));
    InMux I__3699 (
            .O(N__24946),
            .I(N__24922));
    InMux I__3698 (
            .O(N__24945),
            .I(N__24919));
    InMux I__3697 (
            .O(N__24944),
            .I(N__24910));
    InMux I__3696 (
            .O(N__24943),
            .I(N__24910));
    InMux I__3695 (
            .O(N__24942),
            .I(N__24910));
    InMux I__3694 (
            .O(N__24941),
            .I(N__24910));
    InMux I__3693 (
            .O(N__24940),
            .I(N__24897));
    InMux I__3692 (
            .O(N__24939),
            .I(N__24897));
    InMux I__3691 (
            .O(N__24938),
            .I(N__24897));
    InMux I__3690 (
            .O(N__24935),
            .I(N__24897));
    InMux I__3689 (
            .O(N__24932),
            .I(N__24897));
    InMux I__3688 (
            .O(N__24929),
            .I(N__24897));
    InMux I__3687 (
            .O(N__24926),
            .I(N__24892));
    InMux I__3686 (
            .O(N__24925),
            .I(N__24892));
    LocalMux I__3685 (
            .O(N__24922),
            .I(N__24889));
    LocalMux I__3684 (
            .O(N__24919),
            .I(N__24886));
    LocalMux I__3683 (
            .O(N__24910),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0Z0Z_6 ));
    LocalMux I__3682 (
            .O(N__24897),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0Z0Z_6 ));
    LocalMux I__3681 (
            .O(N__24892),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0Z0Z_6 ));
    Odrv4 I__3680 (
            .O(N__24889),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0Z0Z_6 ));
    Odrv12 I__3679 (
            .O(N__24886),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0Z0Z_6 ));
    CascadeMux I__3678 (
            .O(N__24875),
            .I(N__24872));
    InMux I__3677 (
            .O(N__24872),
            .I(N__24856));
    InMux I__3676 (
            .O(N__24871),
            .I(N__24856));
    InMux I__3675 (
            .O(N__24870),
            .I(N__24853));
    InMux I__3674 (
            .O(N__24869),
            .I(N__24846));
    InMux I__3673 (
            .O(N__24868),
            .I(N__24846));
    InMux I__3672 (
            .O(N__24867),
            .I(N__24846));
    InMux I__3671 (
            .O(N__24866),
            .I(N__24839));
    InMux I__3670 (
            .O(N__24865),
            .I(N__24839));
    InMux I__3669 (
            .O(N__24864),
            .I(N__24839));
    InMux I__3668 (
            .O(N__24863),
            .I(N__24836));
    InMux I__3667 (
            .O(N__24862),
            .I(N__24831));
    InMux I__3666 (
            .O(N__24861),
            .I(N__24831));
    LocalMux I__3665 (
            .O(N__24856),
            .I(\phase_controller_inst1.stoper_hc.N_327 ));
    LocalMux I__3664 (
            .O(N__24853),
            .I(\phase_controller_inst1.stoper_hc.N_327 ));
    LocalMux I__3663 (
            .O(N__24846),
            .I(\phase_controller_inst1.stoper_hc.N_327 ));
    LocalMux I__3662 (
            .O(N__24839),
            .I(\phase_controller_inst1.stoper_hc.N_327 ));
    LocalMux I__3661 (
            .O(N__24836),
            .I(\phase_controller_inst1.stoper_hc.N_327 ));
    LocalMux I__3660 (
            .O(N__24831),
            .I(\phase_controller_inst1.stoper_hc.N_327 ));
    InMux I__3659 (
            .O(N__24818),
            .I(N__24815));
    LocalMux I__3658 (
            .O(N__24815),
            .I(N__24812));
    Span4Mux_v I__3657 (
            .O(N__24812),
            .I(N__24809));
    Odrv4 I__3656 (
            .O(N__24809),
            .I(\phase_controller_inst2.stoper_hc.un6_running_1 ));
    InMux I__3655 (
            .O(N__24806),
            .I(N__24802));
    CascadeMux I__3654 (
            .O(N__24805),
            .I(N__24798));
    LocalMux I__3653 (
            .O(N__24802),
            .I(N__24795));
    InMux I__3652 (
            .O(N__24801),
            .I(N__24792));
    InMux I__3651 (
            .O(N__24798),
            .I(N__24789));
    Span4Mux_h I__3650 (
            .O(N__24795),
            .I(N__24786));
    LocalMux I__3649 (
            .O(N__24792),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__3648 (
            .O(N__24789),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__3647 (
            .O(N__24786),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    CascadeMux I__3646 (
            .O(N__24779),
            .I(N__24776));
    InMux I__3645 (
            .O(N__24776),
            .I(N__24773));
    LocalMux I__3644 (
            .O(N__24773),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ));
    InMux I__3643 (
            .O(N__24770),
            .I(N__24767));
    LocalMux I__3642 (
            .O(N__24767),
            .I(\phase_controller_inst2.stoper_hc.un6_running_2 ));
    InMux I__3641 (
            .O(N__24764),
            .I(N__24760));
    InMux I__3640 (
            .O(N__24763),
            .I(N__24757));
    LocalMux I__3639 (
            .O(N__24760),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__3638 (
            .O(N__24757),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    CascadeMux I__3637 (
            .O(N__24752),
            .I(N__24749));
    InMux I__3636 (
            .O(N__24749),
            .I(N__24746));
    LocalMux I__3635 (
            .O(N__24746),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ));
    InMux I__3634 (
            .O(N__24743),
            .I(N__24739));
    InMux I__3633 (
            .O(N__24742),
            .I(N__24736));
    LocalMux I__3632 (
            .O(N__24739),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__3631 (
            .O(N__24736),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__3630 (
            .O(N__24731),
            .I(N__24728));
    LocalMux I__3629 (
            .O(N__24728),
            .I(N__24725));
    Span4Mux_v I__3628 (
            .O(N__24725),
            .I(N__24722));
    Odrv4 I__3627 (
            .O(N__24722),
            .I(\phase_controller_inst2.stoper_hc.un6_running_3 ));
    CascadeMux I__3626 (
            .O(N__24719),
            .I(N__24716));
    InMux I__3625 (
            .O(N__24716),
            .I(N__24713));
    LocalMux I__3624 (
            .O(N__24713),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ));
    InMux I__3623 (
            .O(N__24710),
            .I(N__24707));
    LocalMux I__3622 (
            .O(N__24707),
            .I(N__24703));
    InMux I__3621 (
            .O(N__24706),
            .I(N__24700));
    Sp12to4 I__3620 (
            .O(N__24703),
            .I(N__24697));
    LocalMux I__3619 (
            .O(N__24700),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    Odrv12 I__3618 (
            .O(N__24697),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__3617 (
            .O(N__24692),
            .I(N__24689));
    LocalMux I__3616 (
            .O(N__24689),
            .I(\phase_controller_inst2.stoper_hc.un6_running_4 ));
    CascadeMux I__3615 (
            .O(N__24686),
            .I(N__24683));
    InMux I__3614 (
            .O(N__24683),
            .I(N__24680));
    LocalMux I__3613 (
            .O(N__24680),
            .I(N__24677));
    Odrv4 I__3612 (
            .O(N__24677),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ));
    InMux I__3611 (
            .O(N__24674),
            .I(N__24671));
    LocalMux I__3610 (
            .O(N__24671),
            .I(N__24668));
    Odrv4 I__3609 (
            .O(N__24668),
            .I(\phase_controller_inst2.stoper_hc.un6_running_5 ));
    InMux I__3608 (
            .O(N__24665),
            .I(N__24661));
    InMux I__3607 (
            .O(N__24664),
            .I(N__24658));
    LocalMux I__3606 (
            .O(N__24661),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__3605 (
            .O(N__24658),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    CascadeMux I__3604 (
            .O(N__24653),
            .I(N__24650));
    InMux I__3603 (
            .O(N__24650),
            .I(N__24647));
    LocalMux I__3602 (
            .O(N__24647),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ));
    InMux I__3601 (
            .O(N__24644),
            .I(N__24640));
    InMux I__3600 (
            .O(N__24643),
            .I(N__24637));
    LocalMux I__3599 (
            .O(N__24640),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__3598 (
            .O(N__24637),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    CascadeMux I__3597 (
            .O(N__24632),
            .I(N__24629));
    InMux I__3596 (
            .O(N__24629),
            .I(N__24626));
    LocalMux I__3595 (
            .O(N__24626),
            .I(N__24623));
    Odrv4 I__3594 (
            .O(N__24623),
            .I(\phase_controller_inst2.stoper_hc.un6_running_6 ));
    InMux I__3593 (
            .O(N__24620),
            .I(N__24617));
    LocalMux I__3592 (
            .O(N__24617),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ));
    CascadeMux I__3591 (
            .O(N__24614),
            .I(N__24611));
    InMux I__3590 (
            .O(N__24611),
            .I(N__24608));
    LocalMux I__3589 (
            .O(N__24608),
            .I(N__24605));
    Odrv4 I__3588 (
            .O(N__24605),
            .I(\phase_controller_inst2.stoper_hc.un6_running_7 ));
    InMux I__3587 (
            .O(N__24602),
            .I(N__24598));
    InMux I__3586 (
            .O(N__24601),
            .I(N__24595));
    LocalMux I__3585 (
            .O(N__24598),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__3584 (
            .O(N__24595),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__3583 (
            .O(N__24590),
            .I(N__24587));
    LocalMux I__3582 (
            .O(N__24587),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ));
    CascadeMux I__3581 (
            .O(N__24584),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6_cascade_ ));
    CascadeMux I__3580 (
            .O(N__24581),
            .I(N__24577));
    InMux I__3579 (
            .O(N__24580),
            .I(N__24573));
    InMux I__3578 (
            .O(N__24577),
            .I(N__24570));
    InMux I__3577 (
            .O(N__24576),
            .I(N__24567));
    LocalMux I__3576 (
            .O(N__24573),
            .I(elapsed_time_ns_1_RNIIU2KD1_0_6));
    LocalMux I__3575 (
            .O(N__24570),
            .I(elapsed_time_ns_1_RNIIU2KD1_0_6));
    LocalMux I__3574 (
            .O(N__24567),
            .I(elapsed_time_ns_1_RNIIU2KD1_0_6));
    CascadeMux I__3573 (
            .O(N__24560),
            .I(elapsed_time_ns_1_RNIIU2KD1_0_6_cascade_));
    InMux I__3572 (
            .O(N__24557),
            .I(N__24552));
    InMux I__3571 (
            .O(N__24556),
            .I(N__24547));
    InMux I__3570 (
            .O(N__24555),
            .I(N__24547));
    LocalMux I__3569 (
            .O(N__24552),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2 ));
    LocalMux I__3568 (
            .O(N__24547),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2 ));
    CascadeMux I__3567 (
            .O(N__24542),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_ ));
    CascadeMux I__3566 (
            .O(N__24539),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0Z0Z_6_cascade_ ));
    CascadeMux I__3565 (
            .O(N__24536),
            .I(N__24532));
    InMux I__3564 (
            .O(N__24535),
            .I(N__24529));
    InMux I__3563 (
            .O(N__24532),
            .I(N__24526));
    LocalMux I__3562 (
            .O(N__24529),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1 ));
    LocalMux I__3561 (
            .O(N__24526),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1 ));
    CascadeMux I__3560 (
            .O(N__24521),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_ ));
    InMux I__3559 (
            .O(N__24518),
            .I(N__24512));
    InMux I__3558 (
            .O(N__24517),
            .I(N__24509));
    InMux I__3557 (
            .O(N__24516),
            .I(N__24504));
    InMux I__3556 (
            .O(N__24515),
            .I(N__24504));
    LocalMux I__3555 (
            .O(N__24512),
            .I(elapsed_time_ns_1_RNIDP2KD1_0_1));
    LocalMux I__3554 (
            .O(N__24509),
            .I(elapsed_time_ns_1_RNIDP2KD1_0_1));
    LocalMux I__3553 (
            .O(N__24504),
            .I(elapsed_time_ns_1_RNIDP2KD1_0_1));
    InMux I__3552 (
            .O(N__24497),
            .I(N__24493));
    InMux I__3551 (
            .O(N__24496),
            .I(N__24490));
    LocalMux I__3550 (
            .O(N__24493),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2 ));
    LocalMux I__3549 (
            .O(N__24490),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2 ));
    CascadeMux I__3548 (
            .O(N__24485),
            .I(elapsed_time_ns_1_RNIQ4OD11_0_31_cascade_));
    InMux I__3547 (
            .O(N__24482),
            .I(N__24479));
    LocalMux I__3546 (
            .O(N__24479),
            .I(N__24476));
    Odrv4 I__3545 (
            .O(N__24476),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_1Z0Z_9 ));
    CascadeMux I__3544 (
            .O(N__24473),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_1Z0Z_9_cascade_ ));
    InMux I__3543 (
            .O(N__24470),
            .I(N__24462));
    InMux I__3542 (
            .O(N__24469),
            .I(N__24462));
    CascadeMux I__3541 (
            .O(N__24468),
            .I(N__24454));
    CascadeMux I__3540 (
            .O(N__24467),
            .I(N__24451));
    LocalMux I__3539 (
            .O(N__24462),
            .I(N__24446));
    InMux I__3538 (
            .O(N__24461),
            .I(N__24441));
    InMux I__3537 (
            .O(N__24460),
            .I(N__24441));
    InMux I__3536 (
            .O(N__24459),
            .I(N__24438));
    InMux I__3535 (
            .O(N__24458),
            .I(N__24431));
    InMux I__3534 (
            .O(N__24457),
            .I(N__24431));
    InMux I__3533 (
            .O(N__24454),
            .I(N__24431));
    InMux I__3532 (
            .O(N__24451),
            .I(N__24428));
    InMux I__3531 (
            .O(N__24450),
            .I(N__24423));
    InMux I__3530 (
            .O(N__24449),
            .I(N__24423));
    Sp12to4 I__3529 (
            .O(N__24446),
            .I(N__24418));
    LocalMux I__3528 (
            .O(N__24441),
            .I(N__24418));
    LocalMux I__3527 (
            .O(N__24438),
            .I(\phase_controller_inst1.stoper_hc.N_315 ));
    LocalMux I__3526 (
            .O(N__24431),
            .I(\phase_controller_inst1.stoper_hc.N_315 ));
    LocalMux I__3525 (
            .O(N__24428),
            .I(\phase_controller_inst1.stoper_hc.N_315 ));
    LocalMux I__3524 (
            .O(N__24423),
            .I(\phase_controller_inst1.stoper_hc.N_315 ));
    Odrv12 I__3523 (
            .O(N__24418),
            .I(\phase_controller_inst1.stoper_hc.N_315 ));
    CascadeMux I__3522 (
            .O(N__24407),
            .I(N__24403));
    InMux I__3521 (
            .O(N__24406),
            .I(N__24400));
    InMux I__3520 (
            .O(N__24403),
            .I(N__24397));
    LocalMux I__3519 (
            .O(N__24400),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3 ));
    LocalMux I__3518 (
            .O(N__24397),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3 ));
    CascadeMux I__3517 (
            .O(N__24392),
            .I(\phase_controller_inst1.stoper_hc.N_283_cascade_ ));
    InMux I__3516 (
            .O(N__24389),
            .I(N__24385));
    InMux I__3515 (
            .O(N__24388),
            .I(N__24382));
    LocalMux I__3514 (
            .O(N__24385),
            .I(\phase_controller_inst1.stoper_hc.N_307 ));
    LocalMux I__3513 (
            .O(N__24382),
            .I(\phase_controller_inst1.stoper_hc.N_307 ));
    InMux I__3512 (
            .O(N__24377),
            .I(N__24374));
    LocalMux I__3511 (
            .O(N__24374),
            .I(N__24371));
    Span4Mux_h I__3510 (
            .O(N__24371),
            .I(N__24368));
    Odrv4 I__3509 (
            .O(N__24368),
            .I(\phase_controller_inst1.stoper_hc.un6_running_7 ));
    CEMux I__3508 (
            .O(N__24365),
            .I(N__24357));
    InMux I__3507 (
            .O(N__24364),
            .I(N__24343));
    InMux I__3506 (
            .O(N__24363),
            .I(N__24343));
    InMux I__3505 (
            .O(N__24362),
            .I(N__24343));
    InMux I__3504 (
            .O(N__24361),
            .I(N__24343));
    InMux I__3503 (
            .O(N__24360),
            .I(N__24340));
    LocalMux I__3502 (
            .O(N__24357),
            .I(N__24337));
    CEMux I__3501 (
            .O(N__24356),
            .I(N__24333));
    InMux I__3500 (
            .O(N__24355),
            .I(N__24314));
    InMux I__3499 (
            .O(N__24354),
            .I(N__24314));
    InMux I__3498 (
            .O(N__24353),
            .I(N__24314));
    InMux I__3497 (
            .O(N__24352),
            .I(N__24314));
    LocalMux I__3496 (
            .O(N__24343),
            .I(N__24309));
    LocalMux I__3495 (
            .O(N__24340),
            .I(N__24309));
    Span4Mux_v I__3494 (
            .O(N__24337),
            .I(N__24306));
    CEMux I__3493 (
            .O(N__24336),
            .I(N__24303));
    LocalMux I__3492 (
            .O(N__24333),
            .I(N__24300));
    InMux I__3491 (
            .O(N__24332),
            .I(N__24293));
    InMux I__3490 (
            .O(N__24331),
            .I(N__24293));
    InMux I__3489 (
            .O(N__24330),
            .I(N__24293));
    InMux I__3488 (
            .O(N__24329),
            .I(N__24284));
    InMux I__3487 (
            .O(N__24328),
            .I(N__24284));
    InMux I__3486 (
            .O(N__24327),
            .I(N__24284));
    InMux I__3485 (
            .O(N__24326),
            .I(N__24284));
    InMux I__3484 (
            .O(N__24325),
            .I(N__24277));
    InMux I__3483 (
            .O(N__24324),
            .I(N__24277));
    InMux I__3482 (
            .O(N__24323),
            .I(N__24277));
    LocalMux I__3481 (
            .O(N__24314),
            .I(N__24270));
    Span4Mux_v I__3480 (
            .O(N__24309),
            .I(N__24270));
    Span4Mux_h I__3479 (
            .O(N__24306),
            .I(N__24270));
    LocalMux I__3478 (
            .O(N__24303),
            .I(N__24263));
    Span4Mux_v I__3477 (
            .O(N__24300),
            .I(N__24263));
    LocalMux I__3476 (
            .O(N__24293),
            .I(N__24263));
    LocalMux I__3475 (
            .O(N__24284),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    LocalMux I__3474 (
            .O(N__24277),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__3473 (
            .O(N__24270),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__3472 (
            .O(N__24263),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    CascadeMux I__3471 (
            .O(N__24254),
            .I(elapsed_time_ns_1_RNI62CED1_0_19_cascade_));
    CascadeMux I__3470 (
            .O(N__24251),
            .I(\phase_controller_inst1.stoper_hc.N_315_cascade_ ));
    CascadeMux I__3469 (
            .O(N__24248),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18_cascade_ ));
    InMux I__3468 (
            .O(N__24245),
            .I(N__24242));
    LocalMux I__3467 (
            .O(N__24242),
            .I(N__24239));
    Odrv4 I__3466 (
            .O(N__24239),
            .I(\phase_controller_inst1.stoper_hc.un6_running_9 ));
    CascadeMux I__3465 (
            .O(N__24236),
            .I(N__24233));
    InMux I__3464 (
            .O(N__24233),
            .I(N__24230));
    LocalMux I__3463 (
            .O(N__24230),
            .I(N__24227));
    Odrv12 I__3462 (
            .O(N__24227),
            .I(\phase_controller_inst1.stoper_hc.un6_running_13 ));
    InMux I__3461 (
            .O(N__24224),
            .I(N__24221));
    LocalMux I__3460 (
            .O(N__24221),
            .I(N__24218));
    Span4Mux_h I__3459 (
            .O(N__24218),
            .I(N__24215));
    Odrv4 I__3458 (
            .O(N__24215),
            .I(\phase_controller_inst1.stoper_hc.un6_running_19 ));
    InMux I__3457 (
            .O(N__24212),
            .I(N__24209));
    LocalMux I__3456 (
            .O(N__24209),
            .I(N__24206));
    Span4Mux_h I__3455 (
            .O(N__24206),
            .I(N__24203));
    Odrv4 I__3454 (
            .O(N__24203),
            .I(\phase_controller_inst1.stoper_hc.un6_running_18 ));
    InMux I__3453 (
            .O(N__24200),
            .I(N__24197));
    LocalMux I__3452 (
            .O(N__24197),
            .I(N__24194));
    Span4Mux_v I__3451 (
            .O(N__24194),
            .I(N__24191));
    Odrv4 I__3450 (
            .O(N__24191),
            .I(\phase_controller_inst1.stoper_hc.un6_running_17 ));
    InMux I__3449 (
            .O(N__24188),
            .I(N__24185));
    LocalMux I__3448 (
            .O(N__24185),
            .I(N__24182));
    Odrv4 I__3447 (
            .O(N__24182),
            .I(\phase_controller_inst1.stoper_hc.un6_running_16 ));
    InMux I__3446 (
            .O(N__24179),
            .I(N__24176));
    LocalMux I__3445 (
            .O(N__24176),
            .I(N__24173));
    Odrv4 I__3444 (
            .O(N__24173),
            .I(\phase_controller_inst1.stoper_hc.un6_running_15 ));
    CascadeMux I__3443 (
            .O(N__24170),
            .I(N__24167));
    InMux I__3442 (
            .O(N__24167),
            .I(N__24164));
    LocalMux I__3441 (
            .O(N__24164),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    InMux I__3440 (
            .O(N__24161),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ));
    InMux I__3439 (
            .O(N__24158),
            .I(N__24155));
    LocalMux I__3438 (
            .O(N__24155),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    InMux I__3437 (
            .O(N__24152),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ));
    InMux I__3436 (
            .O(N__24149),
            .I(bfn_9_12_0_));
    InMux I__3435 (
            .O(N__24146),
            .I(N__24143));
    LocalMux I__3434 (
            .O(N__24143),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ));
    CascadeMux I__3433 (
            .O(N__24140),
            .I(N__24137));
    InMux I__3432 (
            .O(N__24137),
            .I(N__24130));
    InMux I__3431 (
            .O(N__24136),
            .I(N__24130));
    InMux I__3430 (
            .O(N__24135),
            .I(N__24127));
    LocalMux I__3429 (
            .O(N__24130),
            .I(N__24123));
    LocalMux I__3428 (
            .O(N__24127),
            .I(N__24120));
    InMux I__3427 (
            .O(N__24126),
            .I(N__24117));
    Span4Mux_v I__3426 (
            .O(N__24123),
            .I(N__24114));
    Odrv12 I__3425 (
            .O(N__24120),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    LocalMux I__3424 (
            .O(N__24117),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv4 I__3423 (
            .O(N__24114),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    CascadeMux I__3422 (
            .O(N__24107),
            .I(N__24104));
    InMux I__3421 (
            .O(N__24104),
            .I(N__24101));
    LocalMux I__3420 (
            .O(N__24101),
            .I(\current_shift_inst.PI_CTRL.integrator_i_29 ));
    CascadeMux I__3419 (
            .O(N__24098),
            .I(N__24093));
    InMux I__3418 (
            .O(N__24097),
            .I(N__24088));
    InMux I__3417 (
            .O(N__24096),
            .I(N__24088));
    InMux I__3416 (
            .O(N__24093),
            .I(N__24085));
    LocalMux I__3415 (
            .O(N__24088),
            .I(N__24081));
    LocalMux I__3414 (
            .O(N__24085),
            .I(N__24078));
    InMux I__3413 (
            .O(N__24084),
            .I(N__24075));
    Span4Mux_h I__3412 (
            .O(N__24081),
            .I(N__24072));
    Odrv12 I__3411 (
            .O(N__24078),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__3410 (
            .O(N__24075),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__3409 (
            .O(N__24072),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    InMux I__3408 (
            .O(N__24065),
            .I(N__24062));
    LocalMux I__3407 (
            .O(N__24062),
            .I(\current_shift_inst.PI_CTRL.integrator_i_28 ));
    CascadeMux I__3406 (
            .O(N__24059),
            .I(N__24056));
    InMux I__3405 (
            .O(N__24056),
            .I(N__24053));
    LocalMux I__3404 (
            .O(N__24053),
            .I(N__24050));
    Odrv4 I__3403 (
            .O(N__24050),
            .I(\current_shift_inst.PI_CTRL.integrator_i_15 ));
    InMux I__3402 (
            .O(N__24047),
            .I(N__24042));
    InMux I__3401 (
            .O(N__24046),
            .I(N__24035));
    InMux I__3400 (
            .O(N__24045),
            .I(N__24035));
    LocalMux I__3399 (
            .O(N__24042),
            .I(N__24032));
    CascadeMux I__3398 (
            .O(N__24041),
            .I(N__24029));
    CascadeMux I__3397 (
            .O(N__24040),
            .I(N__24026));
    LocalMux I__3396 (
            .O(N__24035),
            .I(N__24023));
    Span4Mux_v I__3395 (
            .O(N__24032),
            .I(N__24020));
    InMux I__3394 (
            .O(N__24029),
            .I(N__24017));
    InMux I__3393 (
            .O(N__24026),
            .I(N__24014));
    Span4Mux_v I__3392 (
            .O(N__24023),
            .I(N__24011));
    Odrv4 I__3391 (
            .O(N__24020),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    LocalMux I__3390 (
            .O(N__24017),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    LocalMux I__3389 (
            .O(N__24014),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__3388 (
            .O(N__24011),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    InMux I__3387 (
            .O(N__24002),
            .I(N__23999));
    LocalMux I__3386 (
            .O(N__23999),
            .I(N__23996));
    Odrv4 I__3385 (
            .O(N__23996),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0 ));
    InMux I__3384 (
            .O(N__23993),
            .I(N__23990));
    LocalMux I__3383 (
            .O(N__23990),
            .I(N__23987));
    Span4Mux_h I__3382 (
            .O(N__23987),
            .I(N__23984));
    Odrv4 I__3381 (
            .O(N__23984),
            .I(\current_shift_inst.PI_CTRL.integrator_i_22 ));
    InMux I__3380 (
            .O(N__23981),
            .I(N__23978));
    LocalMux I__3379 (
            .O(N__23978),
            .I(N__23975));
    Odrv4 I__3378 (
            .O(N__23975),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    InMux I__3377 (
            .O(N__23972),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ));
    CascadeMux I__3376 (
            .O(N__23969),
            .I(N__23966));
    InMux I__3375 (
            .O(N__23966),
            .I(N__23963));
    LocalMux I__3374 (
            .O(N__23963),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    InMux I__3373 (
            .O(N__23960),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ));
    InMux I__3372 (
            .O(N__23957),
            .I(N__23954));
    LocalMux I__3371 (
            .O(N__23954),
            .I(N__23951));
    Span4Mux_v I__3370 (
            .O(N__23951),
            .I(N__23948));
    Odrv4 I__3369 (
            .O(N__23948),
            .I(\current_shift_inst.PI_CTRL.integrator_i_23 ));
    InMux I__3368 (
            .O(N__23945),
            .I(N__23942));
    LocalMux I__3367 (
            .O(N__23942),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    InMux I__3366 (
            .O(N__23939),
            .I(bfn_9_11_0_));
    InMux I__3365 (
            .O(N__23936),
            .I(N__23933));
    LocalMux I__3364 (
            .O(N__23933),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    InMux I__3363 (
            .O(N__23930),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ));
    CascadeMux I__3362 (
            .O(N__23927),
            .I(N__23924));
    InMux I__3361 (
            .O(N__23924),
            .I(N__23921));
    LocalMux I__3360 (
            .O(N__23921),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    InMux I__3359 (
            .O(N__23918),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ));
    CascadeMux I__3358 (
            .O(N__23915),
            .I(N__23912));
    InMux I__3357 (
            .O(N__23912),
            .I(N__23909));
    LocalMux I__3356 (
            .O(N__23909),
            .I(N__23906));
    Odrv12 I__3355 (
            .O(N__23906),
            .I(\current_shift_inst.PI_CTRL.integrator_i_26 ));
    InMux I__3354 (
            .O(N__23903),
            .I(N__23900));
    LocalMux I__3353 (
            .O(N__23900),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    InMux I__3352 (
            .O(N__23897),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ));
    InMux I__3351 (
            .O(N__23894),
            .I(N__23891));
    LocalMux I__3350 (
            .O(N__23891),
            .I(N__23888));
    Span4Mux_h I__3349 (
            .O(N__23888),
            .I(N__23885));
    Odrv4 I__3348 (
            .O(N__23885),
            .I(\current_shift_inst.PI_CTRL.integrator_i_27 ));
    InMux I__3347 (
            .O(N__23882),
            .I(N__23879));
    LocalMux I__3346 (
            .O(N__23879),
            .I(N__23876));
    Odrv4 I__3345 (
            .O(N__23876),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    InMux I__3344 (
            .O(N__23873),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ));
    InMux I__3343 (
            .O(N__23870),
            .I(N__23867));
    LocalMux I__3342 (
            .O(N__23867),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    InMux I__3341 (
            .O(N__23864),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ));
    InMux I__3340 (
            .O(N__23861),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ));
    InMux I__3339 (
            .O(N__23858),
            .I(N__23855));
    LocalMux I__3338 (
            .O(N__23855),
            .I(N__23852));
    Odrv4 I__3337 (
            .O(N__23852),
            .I(\current_shift_inst.PI_CTRL.integrator_i_14 ));
    InMux I__3336 (
            .O(N__23849),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ));
    InMux I__3335 (
            .O(N__23846),
            .I(N__23843));
    LocalMux I__3334 (
            .O(N__23843),
            .I(N__23840));
    Odrv4 I__3333 (
            .O(N__23840),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    InMux I__3332 (
            .O(N__23837),
            .I(bfn_9_10_0_));
    InMux I__3331 (
            .O(N__23834),
            .I(N__23831));
    LocalMux I__3330 (
            .O(N__23831),
            .I(N__23828));
    Odrv4 I__3329 (
            .O(N__23828),
            .I(\current_shift_inst.PI_CTRL.integrator_i_16 ));
    InMux I__3328 (
            .O(N__23825),
            .I(N__23822));
    LocalMux I__3327 (
            .O(N__23822),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    InMux I__3326 (
            .O(N__23819),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ));
    InMux I__3325 (
            .O(N__23816),
            .I(N__23813));
    LocalMux I__3324 (
            .O(N__23813),
            .I(N__23810));
    Odrv4 I__3323 (
            .O(N__23810),
            .I(\current_shift_inst.PI_CTRL.integrator_i_17 ));
    InMux I__3322 (
            .O(N__23807),
            .I(N__23804));
    LocalMux I__3321 (
            .O(N__23804),
            .I(N__23801));
    Odrv4 I__3320 (
            .O(N__23801),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    InMux I__3319 (
            .O(N__23798),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ));
    InMux I__3318 (
            .O(N__23795),
            .I(N__23792));
    LocalMux I__3317 (
            .O(N__23792),
            .I(N__23789));
    Odrv4 I__3316 (
            .O(N__23789),
            .I(\current_shift_inst.PI_CTRL.integrator_i_18 ));
    InMux I__3315 (
            .O(N__23786),
            .I(N__23783));
    LocalMux I__3314 (
            .O(N__23783),
            .I(N__23780));
    Odrv4 I__3313 (
            .O(N__23780),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    InMux I__3312 (
            .O(N__23777),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ));
    InMux I__3311 (
            .O(N__23774),
            .I(N__23771));
    LocalMux I__3310 (
            .O(N__23771),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    InMux I__3309 (
            .O(N__23768),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ));
    InMux I__3308 (
            .O(N__23765),
            .I(N__23762));
    LocalMux I__3307 (
            .O(N__23762),
            .I(N__23759));
    Odrv12 I__3306 (
            .O(N__23759),
            .I(\current_shift_inst.PI_CTRL.integrator_i_20 ));
    CascadeMux I__3305 (
            .O(N__23756),
            .I(N__23753));
    InMux I__3304 (
            .O(N__23753),
            .I(N__23750));
    LocalMux I__3303 (
            .O(N__23750),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    InMux I__3302 (
            .O(N__23747),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ));
    InMux I__3301 (
            .O(N__23744),
            .I(N__23741));
    LocalMux I__3300 (
            .O(N__23741),
            .I(\current_shift_inst.PI_CTRL.integrator_i_5 ));
    CascadeMux I__3299 (
            .O(N__23738),
            .I(N__23735));
    InMux I__3298 (
            .O(N__23735),
            .I(N__23732));
    LocalMux I__3297 (
            .O(N__23732),
            .I(N__23729));
    Odrv4 I__3296 (
            .O(N__23729),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9 ));
    CascadeMux I__3295 (
            .O(N__23726),
            .I(N__23723));
    InMux I__3294 (
            .O(N__23723),
            .I(N__23720));
    LocalMux I__3293 (
            .O(N__23720),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    InMux I__3292 (
            .O(N__23717),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ));
    InMux I__3291 (
            .O(N__23714),
            .I(N__23711));
    LocalMux I__3290 (
            .O(N__23711),
            .I(N__23708));
    Span4Mux_v I__3289 (
            .O(N__23708),
            .I(N__23705));
    Odrv4 I__3288 (
            .O(N__23705),
            .I(\current_shift_inst.PI_CTRL.integrator_i_6 ));
    InMux I__3287 (
            .O(N__23702),
            .I(N__23699));
    LocalMux I__3286 (
            .O(N__23699),
            .I(N__23696));
    Odrv4 I__3285 (
            .O(N__23696),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    InMux I__3284 (
            .O(N__23693),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ));
    InMux I__3283 (
            .O(N__23690),
            .I(N__23687));
    LocalMux I__3282 (
            .O(N__23687),
            .I(\current_shift_inst.PI_CTRL.integrator_i_7 ));
    CascadeMux I__3281 (
            .O(N__23684),
            .I(N__23681));
    InMux I__3280 (
            .O(N__23681),
            .I(N__23678));
    LocalMux I__3279 (
            .O(N__23678),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11 ));
    InMux I__3278 (
            .O(N__23675),
            .I(N__23672));
    LocalMux I__3277 (
            .O(N__23672),
            .I(N__23669));
    Odrv4 I__3276 (
            .O(N__23669),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    InMux I__3275 (
            .O(N__23666),
            .I(bfn_9_9_0_));
    InMux I__3274 (
            .O(N__23663),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ));
    InMux I__3273 (
            .O(N__23660),
            .I(N__23657));
    LocalMux I__3272 (
            .O(N__23657),
            .I(N__23654));
    Span4Mux_h I__3271 (
            .O(N__23654),
            .I(N__23651));
    Odrv4 I__3270 (
            .O(N__23651),
            .I(\current_shift_inst.PI_CTRL.integrator_i_9 ));
    InMux I__3269 (
            .O(N__23648),
            .I(N__23645));
    LocalMux I__3268 (
            .O(N__23645),
            .I(N__23642));
    Odrv4 I__3267 (
            .O(N__23642),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    InMux I__3266 (
            .O(N__23639),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ));
    InMux I__3265 (
            .O(N__23636),
            .I(N__23633));
    LocalMux I__3264 (
            .O(N__23633),
            .I(N__23630));
    Span4Mux_h I__3263 (
            .O(N__23630),
            .I(N__23627));
    Odrv4 I__3262 (
            .O(N__23627),
            .I(\current_shift_inst.PI_CTRL.integrator_i_10 ));
    InMux I__3261 (
            .O(N__23624),
            .I(N__23621));
    LocalMux I__3260 (
            .O(N__23621),
            .I(N__23618));
    Odrv4 I__3259 (
            .O(N__23618),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    InMux I__3258 (
            .O(N__23615),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ));
    InMux I__3257 (
            .O(N__23612),
            .I(N__23609));
    LocalMux I__3256 (
            .O(N__23609),
            .I(\current_shift_inst.PI_CTRL.integrator_i_11 ));
    InMux I__3255 (
            .O(N__23606),
            .I(N__23603));
    LocalMux I__3254 (
            .O(N__23603),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    InMux I__3253 (
            .O(N__23600),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ));
    InMux I__3252 (
            .O(N__23597),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ));
    IoInMux I__3251 (
            .O(N__23594),
            .I(N__23591));
    LocalMux I__3250 (
            .O(N__23591),
            .I(N__23588));
    Span4Mux_s2_v I__3249 (
            .O(N__23588),
            .I(N__23585));
    Span4Mux_v I__3248 (
            .O(N__23585),
            .I(N__23582));
    Odrv4 I__3247 (
            .O(N__23582),
            .I(\delay_measurement_inst.delay_tr_timer.N_434_i ));
    CascadeMux I__3246 (
            .O(N__23579),
            .I(N__23576));
    InMux I__3245 (
            .O(N__23576),
            .I(N__23573));
    LocalMux I__3244 (
            .O(N__23573),
            .I(N__23568));
    InMux I__3243 (
            .O(N__23572),
            .I(N__23565));
    InMux I__3242 (
            .O(N__23571),
            .I(N__23562));
    Span4Mux_v I__3241 (
            .O(N__23568),
            .I(N__23557));
    LocalMux I__3240 (
            .O(N__23565),
            .I(N__23557));
    LocalMux I__3239 (
            .O(N__23562),
            .I(N__23554));
    Span4Mux_h I__3238 (
            .O(N__23557),
            .I(N__23551));
    Span4Mux_h I__3237 (
            .O(N__23554),
            .I(N__23548));
    Span4Mux_v I__3236 (
            .O(N__23551),
            .I(N__23545));
    Odrv4 I__3235 (
            .O(N__23548),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    Odrv4 I__3234 (
            .O(N__23545),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    InMux I__3233 (
            .O(N__23540),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ));
    InMux I__3232 (
            .O(N__23537),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ));
    InMux I__3231 (
            .O(N__23534),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ));
    InMux I__3230 (
            .O(N__23531),
            .I(N__23528));
    LocalMux I__3229 (
            .O(N__23528),
            .I(\current_shift_inst.PI_CTRL.integrator_i_3 ));
    InMux I__3228 (
            .O(N__23525),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ));
    InMux I__3227 (
            .O(N__23522),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ));
    InMux I__3226 (
            .O(N__23519),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ));
    InMux I__3225 (
            .O(N__23516),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ));
    InMux I__3224 (
            .O(N__23513),
            .I(bfn_8_21_0_));
    InMux I__3223 (
            .O(N__23510),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ));
    InMux I__3222 (
            .O(N__23507),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ));
    InMux I__3221 (
            .O(N__23504),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__3220 (
            .O(N__23501),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__3219 (
            .O(N__23498),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__3218 (
            .O(N__23495),
            .I(bfn_8_20_0_));
    InMux I__3217 (
            .O(N__23492),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__3216 (
            .O(N__23489),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__3215 (
            .O(N__23486),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__3214 (
            .O(N__23483),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__3213 (
            .O(N__23480),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__3212 (
            .O(N__23477),
            .I(N__23474));
    LocalMux I__3211 (
            .O(N__23474),
            .I(N__23471));
    Span4Mux_v I__3210 (
            .O(N__23471),
            .I(N__23468));
    Odrv4 I__3209 (
            .O(N__23468),
            .I(\phase_controller_inst1.stoper_hc.un6_running_5 ));
    InMux I__3208 (
            .O(N__23465),
            .I(N__23462));
    LocalMux I__3207 (
            .O(N__23462),
            .I(N__23459));
    Span4Mux_v I__3206 (
            .O(N__23459),
            .I(N__23456));
    Odrv4 I__3205 (
            .O(N__23456),
            .I(\phase_controller_inst1.stoper_hc.un6_running_8 ));
    InMux I__3204 (
            .O(N__23453),
            .I(N__23450));
    LocalMux I__3203 (
            .O(N__23450),
            .I(N__23447));
    Span4Mux_v I__3202 (
            .O(N__23447),
            .I(N__23444));
    Odrv4 I__3201 (
            .O(N__23444),
            .I(\phase_controller_inst1.stoper_hc.un6_running_3 ));
    InMux I__3200 (
            .O(N__23441),
            .I(N__23438));
    LocalMux I__3199 (
            .O(N__23438),
            .I(N__23435));
    Span4Mux_v I__3198 (
            .O(N__23435),
            .I(N__23432));
    Odrv4 I__3197 (
            .O(N__23432),
            .I(\phase_controller_inst1.stoper_hc.un6_running_1 ));
    InMux I__3196 (
            .O(N__23429),
            .I(N__23426));
    LocalMux I__3195 (
            .O(N__23426),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ));
    InMux I__3194 (
            .O(N__23423),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ));
    CascadeMux I__3193 (
            .O(N__23420),
            .I(N__23417));
    InMux I__3192 (
            .O(N__23417),
            .I(N__23414));
    LocalMux I__3191 (
            .O(N__23414),
            .I(N__23411));
    Odrv4 I__3190 (
            .O(N__23411),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNINJBZ0Z21 ));
    InMux I__3189 (
            .O(N__23408),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__3188 (
            .O(N__23405),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__3187 (
            .O(N__23402),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__3186 (
            .O(N__23399),
            .I(N__23396));
    LocalMux I__3185 (
            .O(N__23396),
            .I(N__23393));
    Span4Mux_v I__3184 (
            .O(N__23393),
            .I(N__23390));
    Odrv4 I__3183 (
            .O(N__23390),
            .I(\phase_controller_inst1.stoper_hc.un6_running_6 ));
    InMux I__3182 (
            .O(N__23387),
            .I(N__23384));
    LocalMux I__3181 (
            .O(N__23384),
            .I(N__23381));
    Span4Mux_v I__3180 (
            .O(N__23381),
            .I(N__23378));
    Odrv4 I__3179 (
            .O(N__23378),
            .I(\phase_controller_inst1.stoper_hc.un6_running_2 ));
    InMux I__3178 (
            .O(N__23375),
            .I(N__23372));
    LocalMux I__3177 (
            .O(N__23372),
            .I(N__23369));
    Span4Mux_v I__3176 (
            .O(N__23369),
            .I(N__23366));
    Odrv4 I__3175 (
            .O(N__23366),
            .I(\phase_controller_inst1.stoper_hc.un6_running_4 ));
    InMux I__3174 (
            .O(N__23363),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ));
    InMux I__3173 (
            .O(N__23360),
            .I(N__23356));
    InMux I__3172 (
            .O(N__23359),
            .I(N__23353));
    LocalMux I__3171 (
            .O(N__23356),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__3170 (
            .O(N__23353),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    CascadeMux I__3169 (
            .O(N__23348),
            .I(N__23344));
    CascadeMux I__3168 (
            .O(N__23347),
            .I(N__23340));
    InMux I__3167 (
            .O(N__23344),
            .I(N__23337));
    InMux I__3166 (
            .O(N__23343),
            .I(N__23334));
    InMux I__3165 (
            .O(N__23340),
            .I(N__23331));
    LocalMux I__3164 (
            .O(N__23337),
            .I(N__23326));
    LocalMux I__3163 (
            .O(N__23334),
            .I(N__23326));
    LocalMux I__3162 (
            .O(N__23331),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__3161 (
            .O(N__23326),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__3160 (
            .O(N__23321),
            .I(N__23317));
    InMux I__3159 (
            .O(N__23320),
            .I(N__23314));
    LocalMux I__3158 (
            .O(N__23317),
            .I(\phase_controller_inst1.stoper_hc.running_1_sqmuxa ));
    LocalMux I__3157 (
            .O(N__23314),
            .I(\phase_controller_inst1.stoper_hc.running_1_sqmuxa ));
    InMux I__3156 (
            .O(N__23309),
            .I(N__23306));
    LocalMux I__3155 (
            .O(N__23306),
            .I(N__23303));
    Odrv4 I__3154 (
            .O(N__23303),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ));
    InMux I__3153 (
            .O(N__23300),
            .I(N__23296));
    InMux I__3152 (
            .O(N__23299),
            .I(N__23293));
    LocalMux I__3151 (
            .O(N__23296),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_CO ));
    LocalMux I__3150 (
            .O(N__23293),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_CO ));
    InMux I__3149 (
            .O(N__23288),
            .I(N__23284));
    InMux I__3148 (
            .O(N__23287),
            .I(N__23281));
    LocalMux I__3147 (
            .O(N__23284),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ));
    LocalMux I__3146 (
            .O(N__23281),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ));
    CascadeMux I__3145 (
            .O(N__23276),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ));
    InMux I__3144 (
            .O(N__23273),
            .I(N__23270));
    LocalMux I__3143 (
            .O(N__23270),
            .I(N__23267));
    Odrv4 I__3142 (
            .O(N__23267),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNIQVTIZ0Z1 ));
    InMux I__3141 (
            .O(N__23264),
            .I(N__23259));
    InMux I__3140 (
            .O(N__23263),
            .I(N__23254));
    InMux I__3139 (
            .O(N__23262),
            .I(N__23254));
    LocalMux I__3138 (
            .O(N__23259),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    LocalMux I__3137 (
            .O(N__23254),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    InMux I__3136 (
            .O(N__23249),
            .I(N__23243));
    InMux I__3135 (
            .O(N__23248),
            .I(N__23240));
    InMux I__3134 (
            .O(N__23247),
            .I(N__23235));
    InMux I__3133 (
            .O(N__23246),
            .I(N__23235));
    LocalMux I__3132 (
            .O(N__23243),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    LocalMux I__3131 (
            .O(N__23240),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    LocalMux I__3130 (
            .O(N__23235),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    InMux I__3129 (
            .O(N__23228),
            .I(N__23224));
    InMux I__3128 (
            .O(N__23227),
            .I(N__23221));
    LocalMux I__3127 (
            .O(N__23224),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__3126 (
            .O(N__23221),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__3125 (
            .O(N__23216),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__3124 (
            .O(N__23213),
            .I(N__23209));
    InMux I__3123 (
            .O(N__23212),
            .I(N__23206));
    LocalMux I__3122 (
            .O(N__23209),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__3121 (
            .O(N__23206),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__3120 (
            .O(N__23201),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__3119 (
            .O(N__23198),
            .I(N__23194));
    InMux I__3118 (
            .O(N__23197),
            .I(N__23191));
    LocalMux I__3117 (
            .O(N__23194),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    LocalMux I__3116 (
            .O(N__23191),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__3115 (
            .O(N__23186),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__3114 (
            .O(N__23183),
            .I(N__23179));
    InMux I__3113 (
            .O(N__23182),
            .I(N__23176));
    LocalMux I__3112 (
            .O(N__23179),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    LocalMux I__3111 (
            .O(N__23176),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__3110 (
            .O(N__23171),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__3109 (
            .O(N__23168),
            .I(N__23164));
    InMux I__3108 (
            .O(N__23167),
            .I(N__23161));
    LocalMux I__3107 (
            .O(N__23164),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__3106 (
            .O(N__23161),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__3105 (
            .O(N__23156),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__3104 (
            .O(N__23153),
            .I(N__23149));
    InMux I__3103 (
            .O(N__23152),
            .I(N__23146));
    LocalMux I__3102 (
            .O(N__23149),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__3101 (
            .O(N__23146),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__3100 (
            .O(N__23141),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ));
    InMux I__3099 (
            .O(N__23138),
            .I(N__23134));
    InMux I__3098 (
            .O(N__23137),
            .I(N__23131));
    LocalMux I__3097 (
            .O(N__23134),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    LocalMux I__3096 (
            .O(N__23131),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__3095 (
            .O(N__23126),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ));
    InMux I__3094 (
            .O(N__23123),
            .I(N__23119));
    InMux I__3093 (
            .O(N__23122),
            .I(N__23116));
    LocalMux I__3092 (
            .O(N__23119),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    LocalMux I__3091 (
            .O(N__23116),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__3090 (
            .O(N__23111),
            .I(bfn_8_15_0_));
    InMux I__3089 (
            .O(N__23108),
            .I(N__23104));
    InMux I__3088 (
            .O(N__23107),
            .I(N__23101));
    LocalMux I__3087 (
            .O(N__23104),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__3086 (
            .O(N__23101),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__3085 (
            .O(N__23096),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ));
    InMux I__3084 (
            .O(N__23093),
            .I(N__23089));
    InMux I__3083 (
            .O(N__23092),
            .I(N__23086));
    LocalMux I__3082 (
            .O(N__23089),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__3081 (
            .O(N__23086),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__3080 (
            .O(N__23081),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ));
    CascadeMux I__3079 (
            .O(N__23078),
            .I(N__23075));
    InMux I__3078 (
            .O(N__23075),
            .I(N__23071));
    InMux I__3077 (
            .O(N__23074),
            .I(N__23068));
    LocalMux I__3076 (
            .O(N__23071),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__3075 (
            .O(N__23068),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__3074 (
            .O(N__23063),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__3073 (
            .O(N__23060),
            .I(N__23056));
    InMux I__3072 (
            .O(N__23059),
            .I(N__23053));
    LocalMux I__3071 (
            .O(N__23056),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__3070 (
            .O(N__23053),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__3069 (
            .O(N__23048),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__3068 (
            .O(N__23045),
            .I(N__23041));
    InMux I__3067 (
            .O(N__23044),
            .I(N__23038));
    LocalMux I__3066 (
            .O(N__23041),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__3065 (
            .O(N__23038),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__3064 (
            .O(N__23033),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__3063 (
            .O(N__23030),
            .I(N__23026));
    InMux I__3062 (
            .O(N__23029),
            .I(N__23023));
    LocalMux I__3061 (
            .O(N__23026),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__3060 (
            .O(N__23023),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__3059 (
            .O(N__23018),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__3058 (
            .O(N__23015),
            .I(N__23011));
    InMux I__3057 (
            .O(N__23014),
            .I(N__23008));
    LocalMux I__3056 (
            .O(N__23011),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__3055 (
            .O(N__23008),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__3054 (
            .O(N__23003),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__3053 (
            .O(N__23000),
            .I(N__22996));
    InMux I__3052 (
            .O(N__22999),
            .I(N__22993));
    LocalMux I__3051 (
            .O(N__22996),
            .I(N__22988));
    LocalMux I__3050 (
            .O(N__22993),
            .I(N__22988));
    Odrv4 I__3049 (
            .O(N__22988),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__3048 (
            .O(N__22985),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__3047 (
            .O(N__22982),
            .I(N__22978));
    InMux I__3046 (
            .O(N__22981),
            .I(N__22975));
    LocalMux I__3045 (
            .O(N__22978),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__3044 (
            .O(N__22975),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__3043 (
            .O(N__22970),
            .I(bfn_8_14_0_));
    InMux I__3042 (
            .O(N__22967),
            .I(N__22964));
    LocalMux I__3041 (
            .O(N__22964),
            .I(N__22961));
    Span4Mux_h I__3040 (
            .O(N__22961),
            .I(N__22958));
    Odrv4 I__3039 (
            .O(N__22958),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    CascadeMux I__3038 (
            .O(N__22955),
            .I(N__22946));
    CascadeMux I__3037 (
            .O(N__22954),
            .I(N__22942));
    CascadeMux I__3036 (
            .O(N__22953),
            .I(N__22938));
    CascadeMux I__3035 (
            .O(N__22952),
            .I(N__22930));
    CascadeMux I__3034 (
            .O(N__22951),
            .I(N__22926));
    InMux I__3033 (
            .O(N__22950),
            .I(N__22908));
    InMux I__3032 (
            .O(N__22949),
            .I(N__22908));
    InMux I__3031 (
            .O(N__22946),
            .I(N__22908));
    InMux I__3030 (
            .O(N__22945),
            .I(N__22908));
    InMux I__3029 (
            .O(N__22942),
            .I(N__22908));
    InMux I__3028 (
            .O(N__22941),
            .I(N__22908));
    InMux I__3027 (
            .O(N__22938),
            .I(N__22908));
    InMux I__3026 (
            .O(N__22937),
            .I(N__22908));
    CascadeMux I__3025 (
            .O(N__22936),
            .I(N__22905));
    CascadeMux I__3024 (
            .O(N__22935),
            .I(N__22901));
    CascadeMux I__3023 (
            .O(N__22934),
            .I(N__22897));
    CascadeMux I__3022 (
            .O(N__22933),
            .I(N__22893));
    InMux I__3021 (
            .O(N__22930),
            .I(N__22883));
    InMux I__3020 (
            .O(N__22929),
            .I(N__22883));
    InMux I__3019 (
            .O(N__22926),
            .I(N__22883));
    InMux I__3018 (
            .O(N__22925),
            .I(N__22883));
    LocalMux I__3017 (
            .O(N__22908),
            .I(N__22880));
    InMux I__3016 (
            .O(N__22905),
            .I(N__22863));
    InMux I__3015 (
            .O(N__22904),
            .I(N__22863));
    InMux I__3014 (
            .O(N__22901),
            .I(N__22863));
    InMux I__3013 (
            .O(N__22900),
            .I(N__22863));
    InMux I__3012 (
            .O(N__22897),
            .I(N__22863));
    InMux I__3011 (
            .O(N__22896),
            .I(N__22863));
    InMux I__3010 (
            .O(N__22893),
            .I(N__22863));
    InMux I__3009 (
            .O(N__22892),
            .I(N__22863));
    LocalMux I__3008 (
            .O(N__22883),
            .I(N__22860));
    Span4Mux_v I__3007 (
            .O(N__22880),
            .I(N__22855));
    LocalMux I__3006 (
            .O(N__22863),
            .I(N__22855));
    Span4Mux_h I__3005 (
            .O(N__22860),
            .I(N__22852));
    Odrv4 I__3004 (
            .O(N__22855),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    Odrv4 I__3003 (
            .O(N__22852),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    InMux I__3002 (
            .O(N__22847),
            .I(N__22843));
    InMux I__3001 (
            .O(N__22846),
            .I(N__22840));
    LocalMux I__3000 (
            .O(N__22843),
            .I(\current_shift_inst.PI_CTRL.N_74_16 ));
    LocalMux I__2999 (
            .O(N__22840),
            .I(\current_shift_inst.PI_CTRL.N_74_16 ));
    CascadeMux I__2998 (
            .O(N__22835),
            .I(N__22832));
    InMux I__2997 (
            .O(N__22832),
            .I(N__22828));
    InMux I__2996 (
            .O(N__22831),
            .I(N__22825));
    LocalMux I__2995 (
            .O(N__22828),
            .I(N__22822));
    LocalMux I__2994 (
            .O(N__22825),
            .I(\current_shift_inst.PI_CTRL.N_74_21 ));
    Odrv4 I__2993 (
            .O(N__22822),
            .I(\current_shift_inst.PI_CTRL.N_74_21 ));
    CascadeMux I__2992 (
            .O(N__22817),
            .I(\current_shift_inst.PI_CTRL.N_103_cascade_ ));
    InMux I__2991 (
            .O(N__22814),
            .I(N__22811));
    LocalMux I__2990 (
            .O(N__22811),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ));
    CascadeMux I__2989 (
            .O(N__22808),
            .I(N__22805));
    InMux I__2988 (
            .O(N__22805),
            .I(N__22799));
    InMux I__2987 (
            .O(N__22804),
            .I(N__22799));
    LocalMux I__2986 (
            .O(N__22799),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ));
    CascadeMux I__2985 (
            .O(N__22796),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ));
    InMux I__2984 (
            .O(N__22793),
            .I(N__22786));
    InMux I__2983 (
            .O(N__22792),
            .I(N__22786));
    InMux I__2982 (
            .O(N__22791),
            .I(N__22783));
    LocalMux I__2981 (
            .O(N__22786),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    LocalMux I__2980 (
            .O(N__22783),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    InMux I__2979 (
            .O(N__22778),
            .I(N__22775));
    LocalMux I__2978 (
            .O(N__22775),
            .I(N__22772));
    Odrv12 I__2977 (
            .O(N__22772),
            .I(il_max_comp1_c));
    CascadeMux I__2976 (
            .O(N__22769),
            .I(N__22766));
    InMux I__2975 (
            .O(N__22766),
            .I(N__22763));
    LocalMux I__2974 (
            .O(N__22763),
            .I(N__22758));
    InMux I__2973 (
            .O(N__22762),
            .I(N__22753));
    InMux I__2972 (
            .O(N__22761),
            .I(N__22753));
    Span4Mux_h I__2971 (
            .O(N__22758),
            .I(N__22748));
    LocalMux I__2970 (
            .O(N__22753),
            .I(N__22745));
    InMux I__2969 (
            .O(N__22752),
            .I(N__22740));
    InMux I__2968 (
            .O(N__22751),
            .I(N__22740));
    Odrv4 I__2967 (
            .O(N__22748),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv4 I__2966 (
            .O(N__22745),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    LocalMux I__2965 (
            .O(N__22740),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    CascadeMux I__2964 (
            .O(N__22733),
            .I(\phase_controller_inst2.start_timer_hc_0_sqmuxa_cascade_ ));
    InMux I__2963 (
            .O(N__22730),
            .I(N__22727));
    LocalMux I__2962 (
            .O(N__22727),
            .I(\phase_controller_inst2.start_timer_hc_RNOZ0Z_0 ));
    CascadeMux I__2961 (
            .O(N__22724),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0_cascade_ ));
    CascadeMux I__2960 (
            .O(N__22721),
            .I(N__22718));
    InMux I__2959 (
            .O(N__22718),
            .I(N__22715));
    LocalMux I__2958 (
            .O(N__22715),
            .I(N__22712));
    Odrv4 I__2957 (
            .O(N__22712),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    CascadeMux I__2956 (
            .O(N__22709),
            .I(N__22706));
    InMux I__2955 (
            .O(N__22706),
            .I(N__22703));
    LocalMux I__2954 (
            .O(N__22703),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ));
    CascadeMux I__2953 (
            .O(N__22700),
            .I(N__22697));
    InMux I__2952 (
            .O(N__22697),
            .I(N__22694));
    LocalMux I__2951 (
            .O(N__22694),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ));
    CascadeMux I__2950 (
            .O(N__22691),
            .I(N__22688));
    InMux I__2949 (
            .O(N__22688),
            .I(N__22685));
    LocalMux I__2948 (
            .O(N__22685),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ));
    CascadeMux I__2947 (
            .O(N__22682),
            .I(N__22679));
    InMux I__2946 (
            .O(N__22679),
            .I(N__22676));
    LocalMux I__2945 (
            .O(N__22676),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ));
    InMux I__2944 (
            .O(N__22673),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_19 ));
    CascadeMux I__2943 (
            .O(N__22670),
            .I(N__22667));
    InMux I__2942 (
            .O(N__22667),
            .I(N__22664));
    LocalMux I__2941 (
            .O(N__22664),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    CascadeMux I__2940 (
            .O(N__22661),
            .I(N__22658));
    InMux I__2939 (
            .O(N__22658),
            .I(N__22655));
    LocalMux I__2938 (
            .O(N__22655),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    CascadeMux I__2937 (
            .O(N__22652),
            .I(N__22649));
    InMux I__2936 (
            .O(N__22649),
            .I(N__22646));
    LocalMux I__2935 (
            .O(N__22646),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    InMux I__2934 (
            .O(N__22643),
            .I(N__22640));
    LocalMux I__2933 (
            .O(N__22640),
            .I(N__22637));
    Span4Mux_v I__2932 (
            .O(N__22637),
            .I(N__22634));
    Odrv4 I__2931 (
            .O(N__22634),
            .I(\phase_controller_inst1.stoper_hc.un6_running_10 ));
    CascadeMux I__2930 (
            .O(N__22631),
            .I(N__22628));
    InMux I__2929 (
            .O(N__22628),
            .I(N__22625));
    LocalMux I__2928 (
            .O(N__22625),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    InMux I__2927 (
            .O(N__22622),
            .I(N__22619));
    LocalMux I__2926 (
            .O(N__22619),
            .I(N__22616));
    Span4Mux_h I__2925 (
            .O(N__22616),
            .I(N__22613));
    Odrv4 I__2924 (
            .O(N__22613),
            .I(\phase_controller_inst1.stoper_hc.un6_running_11 ));
    CascadeMux I__2923 (
            .O(N__22610),
            .I(N__22607));
    InMux I__2922 (
            .O(N__22607),
            .I(N__22604));
    LocalMux I__2921 (
            .O(N__22604),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    InMux I__2920 (
            .O(N__22601),
            .I(N__22598));
    LocalMux I__2919 (
            .O(N__22598),
            .I(N__22595));
    Span4Mux_h I__2918 (
            .O(N__22595),
            .I(N__22592));
    Odrv4 I__2917 (
            .O(N__22592),
            .I(\phase_controller_inst1.stoper_hc.un6_running_12 ));
    CascadeMux I__2916 (
            .O(N__22589),
            .I(N__22586));
    InMux I__2915 (
            .O(N__22586),
            .I(N__22583));
    LocalMux I__2914 (
            .O(N__22583),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    InMux I__2913 (
            .O(N__22580),
            .I(N__22577));
    LocalMux I__2912 (
            .O(N__22577),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    InMux I__2911 (
            .O(N__22574),
            .I(N__22571));
    LocalMux I__2910 (
            .O(N__22571),
            .I(N__22568));
    Span4Mux_v I__2909 (
            .O(N__22568),
            .I(N__22565));
    Odrv4 I__2908 (
            .O(N__22565),
            .I(\phase_controller_inst1.stoper_hc.un6_running_14 ));
    CascadeMux I__2907 (
            .O(N__22562),
            .I(N__22559));
    InMux I__2906 (
            .O(N__22559),
            .I(N__22556));
    LocalMux I__2905 (
            .O(N__22556),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    CascadeMux I__2904 (
            .O(N__22553),
            .I(N__22550));
    InMux I__2903 (
            .O(N__22550),
            .I(N__22547));
    LocalMux I__2902 (
            .O(N__22547),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    CascadeMux I__2901 (
            .O(N__22544),
            .I(N__22541));
    InMux I__2900 (
            .O(N__22541),
            .I(N__22538));
    LocalMux I__2899 (
            .O(N__22538),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    CascadeMux I__2898 (
            .O(N__22535),
            .I(N__22532));
    InMux I__2897 (
            .O(N__22532),
            .I(N__22529));
    LocalMux I__2896 (
            .O(N__22529),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    CascadeMux I__2895 (
            .O(N__22526),
            .I(N__22523));
    InMux I__2894 (
            .O(N__22523),
            .I(N__22520));
    LocalMux I__2893 (
            .O(N__22520),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    CascadeMux I__2892 (
            .O(N__22517),
            .I(N__22514));
    InMux I__2891 (
            .O(N__22514),
            .I(N__22511));
    LocalMux I__2890 (
            .O(N__22511),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    CascadeMux I__2889 (
            .O(N__22508),
            .I(N__22505));
    InMux I__2888 (
            .O(N__22505),
            .I(N__22502));
    LocalMux I__2887 (
            .O(N__22502),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    InMux I__2886 (
            .O(N__22499),
            .I(N__22496));
    LocalMux I__2885 (
            .O(N__22496),
            .I(N__22493));
    Odrv4 I__2884 (
            .O(N__22493),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    CascadeMux I__2883 (
            .O(N__22490),
            .I(N__22487));
    InMux I__2882 (
            .O(N__22487),
            .I(N__22484));
    LocalMux I__2881 (
            .O(N__22484),
            .I(N__22481));
    Odrv4 I__2880 (
            .O(N__22481),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    InMux I__2879 (
            .O(N__22478),
            .I(N__22475));
    LocalMux I__2878 (
            .O(N__22475),
            .I(N__22472));
    Span4Mux_h I__2877 (
            .O(N__22472),
            .I(N__22469));
    Odrv4 I__2876 (
            .O(N__22469),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ));
    InMux I__2875 (
            .O(N__22466),
            .I(N__22463));
    LocalMux I__2874 (
            .O(N__22463),
            .I(N__22460));
    Odrv12 I__2873 (
            .O(N__22460),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    InMux I__2872 (
            .O(N__22457),
            .I(N__22454));
    LocalMux I__2871 (
            .O(N__22454),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0 ));
    InMux I__2870 (
            .O(N__22451),
            .I(N__22448));
    LocalMux I__2869 (
            .O(N__22448),
            .I(N__22445));
    Span4Mux_v I__2868 (
            .O(N__22445),
            .I(N__22442));
    Odrv4 I__2867 (
            .O(N__22442),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ));
    InMux I__2866 (
            .O(N__22439),
            .I(N__22436));
    LocalMux I__2865 (
            .O(N__22436),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_1 ));
    InMux I__2864 (
            .O(N__22433),
            .I(N__22430));
    LocalMux I__2863 (
            .O(N__22430),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31 ));
    InMux I__2862 (
            .O(N__22427),
            .I(N__22424));
    LocalMux I__2861 (
            .O(N__22424),
            .I(\current_shift_inst.PI_CTRL.N_62 ));
    CascadeMux I__2860 (
            .O(N__22421),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_7_cascade_ ));
    InMux I__2859 (
            .O(N__22418),
            .I(N__22415));
    LocalMux I__2858 (
            .O(N__22415),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ));
    InMux I__2857 (
            .O(N__22412),
            .I(N__22409));
    LocalMux I__2856 (
            .O(N__22409),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_18 ));
    CascadeMux I__2855 (
            .O(N__22406),
            .I(N__22403));
    InMux I__2854 (
            .O(N__22403),
            .I(N__22400));
    LocalMux I__2853 (
            .O(N__22400),
            .I(N__22397));
    Span4Mux_v I__2852 (
            .O(N__22397),
            .I(N__22394));
    Odrv4 I__2851 (
            .O(N__22394),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    InMux I__2850 (
            .O(N__22391),
            .I(N__22388));
    LocalMux I__2849 (
            .O(N__22388),
            .I(N__22385));
    Odrv4 I__2848 (
            .O(N__22385),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31 ));
    InMux I__2847 (
            .O(N__22382),
            .I(N__22379));
    LocalMux I__2846 (
            .O(N__22379),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ));
    InMux I__2845 (
            .O(N__22376),
            .I(N__22373));
    LocalMux I__2844 (
            .O(N__22373),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12 ));
    CascadeMux I__2843 (
            .O(N__22370),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_16_cascade_ ));
    CascadeMux I__2842 (
            .O(N__22367),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_20_cascade_ ));
    CascadeMux I__2841 (
            .O(N__22364),
            .I(\current_shift_inst.PI_CTRL.N_75_cascade_ ));
    InMux I__2840 (
            .O(N__22361),
            .I(N__22355));
    InMux I__2839 (
            .O(N__22360),
            .I(N__22355));
    LocalMux I__2838 (
            .O(N__22355),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    InMux I__2837 (
            .O(N__22352),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ));
    CascadeMux I__2836 (
            .O(N__22349),
            .I(N__22346));
    InMux I__2835 (
            .O(N__22346),
            .I(N__22340));
    InMux I__2834 (
            .O(N__22345),
            .I(N__22340));
    LocalMux I__2833 (
            .O(N__22340),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    InMux I__2832 (
            .O(N__22337),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    InMux I__2831 (
            .O(N__22334),
            .I(N__22331));
    LocalMux I__2830 (
            .O(N__22331),
            .I(N__22327));
    InMux I__2829 (
            .O(N__22330),
            .I(N__22324));
    Odrv4 I__2828 (
            .O(N__22327),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    LocalMux I__2827 (
            .O(N__22324),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    InMux I__2826 (
            .O(N__22319),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    CascadeMux I__2825 (
            .O(N__22316),
            .I(N__22313));
    InMux I__2824 (
            .O(N__22313),
            .I(N__22307));
    InMux I__2823 (
            .O(N__22312),
            .I(N__22307));
    LocalMux I__2822 (
            .O(N__22307),
            .I(N__22304));
    Odrv4 I__2821 (
            .O(N__22304),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    InMux I__2820 (
            .O(N__22301),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ));
    InMux I__2819 (
            .O(N__22298),
            .I(N__22295));
    LocalMux I__2818 (
            .O(N__22295),
            .I(N__22291));
    InMux I__2817 (
            .O(N__22294),
            .I(N__22288));
    Odrv4 I__2816 (
            .O(N__22291),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    LocalMux I__2815 (
            .O(N__22288),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    InMux I__2814 (
            .O(N__22283),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    InMux I__2813 (
            .O(N__22280),
            .I(N__22277));
    LocalMux I__2812 (
            .O(N__22277),
            .I(N__22273));
    CascadeMux I__2811 (
            .O(N__22276),
            .I(N__22270));
    Span4Mux_h I__2810 (
            .O(N__22273),
            .I(N__22267));
    InMux I__2809 (
            .O(N__22270),
            .I(N__22264));
    Odrv4 I__2808 (
            .O(N__22267),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    LocalMux I__2807 (
            .O(N__22264),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    InMux I__2806 (
            .O(N__22259),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    InMux I__2805 (
            .O(N__22256),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    InMux I__2804 (
            .O(N__22253),
            .I(N__22249));
    CascadeMux I__2803 (
            .O(N__22252),
            .I(N__22245));
    LocalMux I__2802 (
            .O(N__22249),
            .I(N__22236));
    InMux I__2801 (
            .O(N__22248),
            .I(N__22227));
    InMux I__2800 (
            .O(N__22245),
            .I(N__22227));
    InMux I__2799 (
            .O(N__22244),
            .I(N__22227));
    InMux I__2798 (
            .O(N__22243),
            .I(N__22227));
    InMux I__2797 (
            .O(N__22242),
            .I(N__22224));
    InMux I__2796 (
            .O(N__22241),
            .I(N__22221));
    InMux I__2795 (
            .O(N__22240),
            .I(N__22216));
    InMux I__2794 (
            .O(N__22239),
            .I(N__22216));
    Span4Mux_v I__2793 (
            .O(N__22236),
            .I(N__22204));
    LocalMux I__2792 (
            .O(N__22227),
            .I(N__22204));
    LocalMux I__2791 (
            .O(N__22224),
            .I(N__22204));
    LocalMux I__2790 (
            .O(N__22221),
            .I(N__22204));
    LocalMux I__2789 (
            .O(N__22216),
            .I(N__22204));
    InMux I__2788 (
            .O(N__22215),
            .I(N__22201));
    Span4Mux_v I__2787 (
            .O(N__22204),
            .I(N__22196));
    LocalMux I__2786 (
            .O(N__22201),
            .I(N__22196));
    Span4Mux_h I__2785 (
            .O(N__22196),
            .I(N__22193));
    Odrv4 I__2784 (
            .O(N__22193),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    InMux I__2783 (
            .O(N__22190),
            .I(N__22187));
    LocalMux I__2782 (
            .O(N__22187),
            .I(N__22184));
    Span4Mux_v I__2781 (
            .O(N__22184),
            .I(N__22181));
    Odrv4 I__2780 (
            .O(N__22181),
            .I(il_max_comp2_D1));
    CascadeMux I__2779 (
            .O(N__22178),
            .I(N__22175));
    InMux I__2778 (
            .O(N__22175),
            .I(N__22171));
    InMux I__2777 (
            .O(N__22174),
            .I(N__22168));
    LocalMux I__2776 (
            .O(N__22171),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    LocalMux I__2775 (
            .O(N__22168),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    InMux I__2774 (
            .O(N__22163),
            .I(bfn_5_11_0_));
    InMux I__2773 (
            .O(N__22160),
            .I(N__22157));
    LocalMux I__2772 (
            .O(N__22157),
            .I(N__22153));
    InMux I__2771 (
            .O(N__22156),
            .I(N__22150));
    Odrv4 I__2770 (
            .O(N__22153),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    LocalMux I__2769 (
            .O(N__22150),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    InMux I__2768 (
            .O(N__22145),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ));
    InMux I__2767 (
            .O(N__22142),
            .I(N__22139));
    LocalMux I__2766 (
            .O(N__22139),
            .I(N__22135));
    InMux I__2765 (
            .O(N__22138),
            .I(N__22132));
    Odrv4 I__2764 (
            .O(N__22135),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    LocalMux I__2763 (
            .O(N__22132),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    InMux I__2762 (
            .O(N__22127),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    InMux I__2761 (
            .O(N__22124),
            .I(N__22118));
    InMux I__2760 (
            .O(N__22123),
            .I(N__22118));
    LocalMux I__2759 (
            .O(N__22118),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    InMux I__2758 (
            .O(N__22115),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    CascadeMux I__2757 (
            .O(N__22112),
            .I(N__22108));
    InMux I__2756 (
            .O(N__22111),
            .I(N__22103));
    InMux I__2755 (
            .O(N__22108),
            .I(N__22103));
    LocalMux I__2754 (
            .O(N__22103),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    InMux I__2753 (
            .O(N__22100),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ));
    CascadeMux I__2752 (
            .O(N__22097),
            .I(N__22093));
    InMux I__2751 (
            .O(N__22096),
            .I(N__22088));
    InMux I__2750 (
            .O(N__22093),
            .I(N__22088));
    LocalMux I__2749 (
            .O(N__22088),
            .I(N__22085));
    Odrv4 I__2748 (
            .O(N__22085),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    InMux I__2747 (
            .O(N__22082),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    InMux I__2746 (
            .O(N__22079),
            .I(N__22073));
    InMux I__2745 (
            .O(N__22078),
            .I(N__22073));
    LocalMux I__2744 (
            .O(N__22073),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    InMux I__2743 (
            .O(N__22070),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    InMux I__2742 (
            .O(N__22067),
            .I(N__22063));
    InMux I__2741 (
            .O(N__22066),
            .I(N__22060));
    LocalMux I__2740 (
            .O(N__22063),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    LocalMux I__2739 (
            .O(N__22060),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    InMux I__2738 (
            .O(N__22055),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    CascadeMux I__2737 (
            .O(N__22052),
            .I(N__22049));
    InMux I__2736 (
            .O(N__22049),
            .I(N__22046));
    LocalMux I__2735 (
            .O(N__22046),
            .I(N__22042));
    InMux I__2734 (
            .O(N__22045),
            .I(N__22039));
    Odrv4 I__2733 (
            .O(N__22042),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    LocalMux I__2732 (
            .O(N__22039),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    InMux I__2731 (
            .O(N__22034),
            .I(bfn_5_12_0_));
    InMux I__2730 (
            .O(N__22031),
            .I(N__22026));
    InMux I__2729 (
            .O(N__22030),
            .I(N__22023));
    InMux I__2728 (
            .O(N__22029),
            .I(N__22020));
    LocalMux I__2727 (
            .O(N__22026),
            .I(N__22017));
    LocalMux I__2726 (
            .O(N__22023),
            .I(N__22012));
    LocalMux I__2725 (
            .O(N__22020),
            .I(N__22012));
    Span4Mux_h I__2724 (
            .O(N__22017),
            .I(N__22009));
    Odrv12 I__2723 (
            .O(N__22012),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    Odrv4 I__2722 (
            .O(N__22009),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    InMux I__2721 (
            .O(N__22004),
            .I(bfn_5_10_0_));
    InMux I__2720 (
            .O(N__22001),
            .I(N__21998));
    LocalMux I__2719 (
            .O(N__21998),
            .I(N__21993));
    InMux I__2718 (
            .O(N__21997),
            .I(N__21990));
    InMux I__2717 (
            .O(N__21996),
            .I(N__21987));
    Span4Mux_h I__2716 (
            .O(N__21993),
            .I(N__21984));
    LocalMux I__2715 (
            .O(N__21990),
            .I(N__21979));
    LocalMux I__2714 (
            .O(N__21987),
            .I(N__21979));
    Odrv4 I__2713 (
            .O(N__21984),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    Odrv12 I__2712 (
            .O(N__21979),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    InMux I__2711 (
            .O(N__21974),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ));
    InMux I__2710 (
            .O(N__21971),
            .I(N__21965));
    InMux I__2709 (
            .O(N__21970),
            .I(N__21965));
    LocalMux I__2708 (
            .O(N__21965),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    InMux I__2707 (
            .O(N__21962),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    InMux I__2706 (
            .O(N__21959),
            .I(N__21956));
    LocalMux I__2705 (
            .O(N__21956),
            .I(N__21952));
    InMux I__2704 (
            .O(N__21955),
            .I(N__21949));
    Odrv4 I__2703 (
            .O(N__21952),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    LocalMux I__2702 (
            .O(N__21949),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    InMux I__2701 (
            .O(N__21944),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    CascadeMux I__2700 (
            .O(N__21941),
            .I(N__21938));
    InMux I__2699 (
            .O(N__21938),
            .I(N__21935));
    LocalMux I__2698 (
            .O(N__21935),
            .I(N__21931));
    InMux I__2697 (
            .O(N__21934),
            .I(N__21928));
    Odrv4 I__2696 (
            .O(N__21931),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    LocalMux I__2695 (
            .O(N__21928),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    InMux I__2694 (
            .O(N__21923),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ));
    InMux I__2693 (
            .O(N__21920),
            .I(N__21916));
    InMux I__2692 (
            .O(N__21919),
            .I(N__21913));
    LocalMux I__2691 (
            .O(N__21916),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    LocalMux I__2690 (
            .O(N__21913),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    InMux I__2689 (
            .O(N__21908),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    InMux I__2688 (
            .O(N__21905),
            .I(N__21901));
    InMux I__2687 (
            .O(N__21904),
            .I(N__21898));
    LocalMux I__2686 (
            .O(N__21901),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    LocalMux I__2685 (
            .O(N__21898),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    InMux I__2684 (
            .O(N__21893),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    InMux I__2683 (
            .O(N__21890),
            .I(N__21886));
    InMux I__2682 (
            .O(N__21889),
            .I(N__21883));
    LocalMux I__2681 (
            .O(N__21886),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    LocalMux I__2680 (
            .O(N__21883),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    InMux I__2679 (
            .O(N__21878),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    InMux I__2678 (
            .O(N__21875),
            .I(N__21872));
    LocalMux I__2677 (
            .O(N__21872),
            .I(N__21869));
    Odrv12 I__2676 (
            .O(N__21869),
            .I(il_max_comp2_c));
    InMux I__2675 (
            .O(N__21866),
            .I(N__21863));
    LocalMux I__2674 (
            .O(N__21863),
            .I(N__21860));
    Odrv12 I__2673 (
            .O(N__21860),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    InMux I__2672 (
            .O(N__21857),
            .I(N__21854));
    LocalMux I__2671 (
            .O(N__21854),
            .I(N__21851));
    Odrv12 I__2670 (
            .O(N__21851),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    InMux I__2669 (
            .O(N__21848),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ));
    InMux I__2668 (
            .O(N__21845),
            .I(N__21842));
    LocalMux I__2667 (
            .O(N__21842),
            .I(N__21839));
    Odrv12 I__2666 (
            .O(N__21839),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__2665 (
            .O(N__21836),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ));
    InMux I__2664 (
            .O(N__21833),
            .I(N__21828));
    InMux I__2663 (
            .O(N__21832),
            .I(N__21825));
    InMux I__2662 (
            .O(N__21831),
            .I(N__21822));
    LocalMux I__2661 (
            .O(N__21828),
            .I(N__21817));
    LocalMux I__2660 (
            .O(N__21825),
            .I(N__21817));
    LocalMux I__2659 (
            .O(N__21822),
            .I(N__21812));
    Span4Mux_v I__2658 (
            .O(N__21817),
            .I(N__21812));
    Odrv4 I__2657 (
            .O(N__21812),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__2656 (
            .O(N__21809),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ));
    InMux I__2655 (
            .O(N__21806),
            .I(N__21802));
    InMux I__2654 (
            .O(N__21805),
            .I(N__21798));
    LocalMux I__2653 (
            .O(N__21802),
            .I(N__21794));
    InMux I__2652 (
            .O(N__21801),
            .I(N__21791));
    LocalMux I__2651 (
            .O(N__21798),
            .I(N__21788));
    InMux I__2650 (
            .O(N__21797),
            .I(N__21785));
    Span4Mux_v I__2649 (
            .O(N__21794),
            .I(N__21780));
    LocalMux I__2648 (
            .O(N__21791),
            .I(N__21780));
    Span4Mux_v I__2647 (
            .O(N__21788),
            .I(N__21777));
    LocalMux I__2646 (
            .O(N__21785),
            .I(N__21774));
    Span4Mux_h I__2645 (
            .O(N__21780),
            .I(N__21771));
    Odrv4 I__2644 (
            .O(N__21777),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    Odrv4 I__2643 (
            .O(N__21774),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    Odrv4 I__2642 (
            .O(N__21771),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    InMux I__2641 (
            .O(N__21764),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ));
    CascadeMux I__2640 (
            .O(N__21761),
            .I(N__21758));
    InMux I__2639 (
            .O(N__21758),
            .I(N__21753));
    InMux I__2638 (
            .O(N__21757),
            .I(N__21750));
    InMux I__2637 (
            .O(N__21756),
            .I(N__21747));
    LocalMux I__2636 (
            .O(N__21753),
            .I(N__21740));
    LocalMux I__2635 (
            .O(N__21750),
            .I(N__21740));
    LocalMux I__2634 (
            .O(N__21747),
            .I(N__21740));
    Span4Mux_v I__2633 (
            .O(N__21740),
            .I(N__21737));
    Odrv4 I__2632 (
            .O(N__21737),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    InMux I__2631 (
            .O(N__21734),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    InMux I__2630 (
            .O(N__21731),
            .I(N__21726));
    InMux I__2629 (
            .O(N__21730),
            .I(N__21723));
    InMux I__2628 (
            .O(N__21729),
            .I(N__21720));
    LocalMux I__2627 (
            .O(N__21726),
            .I(N__21715));
    LocalMux I__2626 (
            .O(N__21723),
            .I(N__21715));
    LocalMux I__2625 (
            .O(N__21720),
            .I(N__21712));
    Span4Mux_h I__2624 (
            .O(N__21715),
            .I(N__21709));
    Span4Mux_h I__2623 (
            .O(N__21712),
            .I(N__21706));
    Odrv4 I__2622 (
            .O(N__21709),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    Odrv4 I__2621 (
            .O(N__21706),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    InMux I__2620 (
            .O(N__21701),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    InMux I__2619 (
            .O(N__21698),
            .I(N__21693));
    InMux I__2618 (
            .O(N__21697),
            .I(N__21690));
    InMux I__2617 (
            .O(N__21696),
            .I(N__21687));
    LocalMux I__2616 (
            .O(N__21693),
            .I(N__21684));
    LocalMux I__2615 (
            .O(N__21690),
            .I(N__21679));
    LocalMux I__2614 (
            .O(N__21687),
            .I(N__21679));
    Span4Mux_h I__2613 (
            .O(N__21684),
            .I(N__21676));
    Span4Mux_h I__2612 (
            .O(N__21679),
            .I(N__21673));
    Odrv4 I__2611 (
            .O(N__21676),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    Odrv4 I__2610 (
            .O(N__21673),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    InMux I__2609 (
            .O(N__21668),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    InMux I__2608 (
            .O(N__21665),
            .I(N__21662));
    LocalMux I__2607 (
            .O(N__21662),
            .I(N__21659));
    Odrv4 I__2606 (
            .O(N__21659),
            .I(\pwm_generator_inst.thresholdZ0Z_9 ));
    InMux I__2605 (
            .O(N__21656),
            .I(N__21653));
    LocalMux I__2604 (
            .O(N__21653),
            .I(N__21650));
    Span4Mux_h I__2603 (
            .O(N__21650),
            .I(N__21647));
    Odrv4 I__2602 (
            .O(N__21647),
            .I(\pwm_generator_inst.thresholdZ0Z_3 ));
    CascadeMux I__2601 (
            .O(N__21644),
            .I(N__21641));
    InMux I__2600 (
            .O(N__21641),
            .I(N__21638));
    LocalMux I__2599 (
            .O(N__21638),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ));
    InMux I__2598 (
            .O(N__21635),
            .I(N__21632));
    LocalMux I__2597 (
            .O(N__21632),
            .I(N__21629));
    Odrv4 I__2596 (
            .O(N__21629),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_2 ));
    InMux I__2595 (
            .O(N__21626),
            .I(N__21623));
    LocalMux I__2594 (
            .O(N__21623),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ));
    InMux I__2593 (
            .O(N__21620),
            .I(N__21617));
    LocalMux I__2592 (
            .O(N__21617),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_3 ));
    InMux I__2591 (
            .O(N__21614),
            .I(N__21611));
    LocalMux I__2590 (
            .O(N__21611),
            .I(N__21608));
    Span4Mux_h I__2589 (
            .O(N__21608),
            .I(N__21605));
    Odrv4 I__2588 (
            .O(N__21605),
            .I(\pwm_generator_inst.thresholdZ0Z_8 ));
    InMux I__2587 (
            .O(N__21602),
            .I(N__21599));
    LocalMux I__2586 (
            .O(N__21599),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ));
    InMux I__2585 (
            .O(N__21596),
            .I(N__21593));
    LocalMux I__2584 (
            .O(N__21593),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_8 ));
    InMux I__2583 (
            .O(N__21590),
            .I(N__21577));
    InMux I__2582 (
            .O(N__21589),
            .I(N__21577));
    InMux I__2581 (
            .O(N__21588),
            .I(N__21572));
    InMux I__2580 (
            .O(N__21587),
            .I(N__21572));
    InMux I__2579 (
            .O(N__21586),
            .I(N__21561));
    InMux I__2578 (
            .O(N__21585),
            .I(N__21561));
    InMux I__2577 (
            .O(N__21584),
            .I(N__21561));
    InMux I__2576 (
            .O(N__21583),
            .I(N__21561));
    InMux I__2575 (
            .O(N__21582),
            .I(N__21561));
    LocalMux I__2574 (
            .O(N__21577),
            .I(N__21558));
    LocalMux I__2573 (
            .O(N__21572),
            .I(N__21555));
    LocalMux I__2572 (
            .O(N__21561),
            .I(N__21551));
    Span4Mux_v I__2571 (
            .O(N__21558),
            .I(N__21546));
    Span4Mux_v I__2570 (
            .O(N__21555),
            .I(N__21546));
    InMux I__2569 (
            .O(N__21554),
            .I(N__21543));
    Span4Mux_v I__2568 (
            .O(N__21551),
            .I(N__21540));
    Span4Mux_v I__2567 (
            .O(N__21546),
            .I(N__21537));
    LocalMux I__2566 (
            .O(N__21543),
            .I(\pwm_generator_inst.N_16 ));
    Odrv4 I__2565 (
            .O(N__21540),
            .I(\pwm_generator_inst.N_16 ));
    Odrv4 I__2564 (
            .O(N__21537),
            .I(\pwm_generator_inst.N_16 ));
    InMux I__2563 (
            .O(N__21530),
            .I(N__21522));
    InMux I__2562 (
            .O(N__21529),
            .I(N__21522));
    InMux I__2561 (
            .O(N__21528),
            .I(N__21517));
    InMux I__2560 (
            .O(N__21527),
            .I(N__21517));
    LocalMux I__2559 (
            .O(N__21522),
            .I(N__21509));
    LocalMux I__2558 (
            .O(N__21517),
            .I(N__21506));
    InMux I__2557 (
            .O(N__21516),
            .I(N__21495));
    InMux I__2556 (
            .O(N__21515),
            .I(N__21495));
    InMux I__2555 (
            .O(N__21514),
            .I(N__21495));
    InMux I__2554 (
            .O(N__21513),
            .I(N__21495));
    InMux I__2553 (
            .O(N__21512),
            .I(N__21495));
    Span4Mux_v I__2552 (
            .O(N__21509),
            .I(N__21490));
    Span4Mux_v I__2551 (
            .O(N__21506),
            .I(N__21490));
    LocalMux I__2550 (
            .O(N__21495),
            .I(N__21487));
    Span4Mux_v I__2549 (
            .O(N__21490),
            .I(N__21483));
    Span4Mux_v I__2548 (
            .O(N__21487),
            .I(N__21480));
    InMux I__2547 (
            .O(N__21486),
            .I(N__21477));
    Odrv4 I__2546 (
            .O(N__21483),
            .I(\pwm_generator_inst.N_17 ));
    Odrv4 I__2545 (
            .O(N__21480),
            .I(\pwm_generator_inst.N_17 ));
    LocalMux I__2544 (
            .O(N__21477),
            .I(\pwm_generator_inst.N_17 ));
    CascadeMux I__2543 (
            .O(N__21470),
            .I(N__21465));
    CascadeMux I__2542 (
            .O(N__21469),
            .I(N__21461));
    CascadeMux I__2541 (
            .O(N__21468),
            .I(N__21458));
    InMux I__2540 (
            .O(N__21465),
            .I(N__21453));
    InMux I__2539 (
            .O(N__21464),
            .I(N__21453));
    InMux I__2538 (
            .O(N__21461),
            .I(N__21448));
    InMux I__2537 (
            .O(N__21458),
            .I(N__21448));
    LocalMux I__2536 (
            .O(N__21453),
            .I(N__21445));
    LocalMux I__2535 (
            .O(N__21448),
            .I(N__21442));
    Span4Mux_v I__2534 (
            .O(N__21445),
            .I(N__21431));
    Span4Mux_h I__2533 (
            .O(N__21442),
            .I(N__21428));
    InMux I__2532 (
            .O(N__21441),
            .I(N__21423));
    InMux I__2531 (
            .O(N__21440),
            .I(N__21423));
    CascadeMux I__2530 (
            .O(N__21439),
            .I(N__21420));
    CascadeMux I__2529 (
            .O(N__21438),
            .I(N__21417));
    CascadeMux I__2528 (
            .O(N__21437),
            .I(N__21414));
    CascadeMux I__2527 (
            .O(N__21436),
            .I(N__21411));
    CascadeMux I__2526 (
            .O(N__21435),
            .I(N__21408));
    CascadeMux I__2525 (
            .O(N__21434),
            .I(N__21405));
    Span4Mux_h I__2524 (
            .O(N__21431),
            .I(N__21398));
    Span4Mux_v I__2523 (
            .O(N__21428),
            .I(N__21398));
    LocalMux I__2522 (
            .O(N__21423),
            .I(N__21398));
    InMux I__2521 (
            .O(N__21420),
            .I(N__21392));
    InMux I__2520 (
            .O(N__21417),
            .I(N__21385));
    InMux I__2519 (
            .O(N__21414),
            .I(N__21385));
    InMux I__2518 (
            .O(N__21411),
            .I(N__21385));
    InMux I__2517 (
            .O(N__21408),
            .I(N__21380));
    InMux I__2516 (
            .O(N__21405),
            .I(N__21380));
    Span4Mux_v I__2515 (
            .O(N__21398),
            .I(N__21376));
    InMux I__2514 (
            .O(N__21397),
            .I(N__21369));
    InMux I__2513 (
            .O(N__21396),
            .I(N__21369));
    InMux I__2512 (
            .O(N__21395),
            .I(N__21369));
    LocalMux I__2511 (
            .O(N__21392),
            .I(N__21362));
    LocalMux I__2510 (
            .O(N__21385),
            .I(N__21362));
    LocalMux I__2509 (
            .O(N__21380),
            .I(N__21362));
    CascadeMux I__2508 (
            .O(N__21379),
            .I(N__21359));
    Span4Mux_s1_h I__2507 (
            .O(N__21376),
            .I(N__21338));
    LocalMux I__2506 (
            .O(N__21369),
            .I(N__21338));
    Span12Mux_v I__2505 (
            .O(N__21362),
            .I(N__21335));
    InMux I__2504 (
            .O(N__21359),
            .I(N__21332));
    InMux I__2503 (
            .O(N__21358),
            .I(N__21329));
    InMux I__2502 (
            .O(N__21357),
            .I(N__21312));
    InMux I__2501 (
            .O(N__21356),
            .I(N__21312));
    InMux I__2500 (
            .O(N__21355),
            .I(N__21312));
    InMux I__2499 (
            .O(N__21354),
            .I(N__21312));
    InMux I__2498 (
            .O(N__21353),
            .I(N__21312));
    InMux I__2497 (
            .O(N__21352),
            .I(N__21312));
    InMux I__2496 (
            .O(N__21351),
            .I(N__21312));
    InMux I__2495 (
            .O(N__21350),
            .I(N__21312));
    InMux I__2494 (
            .O(N__21349),
            .I(N__21297));
    InMux I__2493 (
            .O(N__21348),
            .I(N__21297));
    InMux I__2492 (
            .O(N__21347),
            .I(N__21297));
    InMux I__2491 (
            .O(N__21346),
            .I(N__21297));
    InMux I__2490 (
            .O(N__21345),
            .I(N__21297));
    InMux I__2489 (
            .O(N__21344),
            .I(N__21297));
    InMux I__2488 (
            .O(N__21343),
            .I(N__21297));
    Span4Mux_v I__2487 (
            .O(N__21338),
            .I(N__21294));
    Odrv12 I__2486 (
            .O(N__21335),
            .I(N_19_1));
    LocalMux I__2485 (
            .O(N__21332),
            .I(N_19_1));
    LocalMux I__2484 (
            .O(N__21329),
            .I(N_19_1));
    LocalMux I__2483 (
            .O(N__21312),
            .I(N_19_1));
    LocalMux I__2482 (
            .O(N__21297),
            .I(N_19_1));
    Odrv4 I__2481 (
            .O(N__21294),
            .I(N_19_1));
    InMux I__2480 (
            .O(N__21281),
            .I(N__21278));
    LocalMux I__2479 (
            .O(N__21278),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ));
    InMux I__2478 (
            .O(N__21275),
            .I(N__21272));
    LocalMux I__2477 (
            .O(N__21272),
            .I(N__21269));
    Odrv4 I__2476 (
            .O(N__21269),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_9 ));
    InMux I__2475 (
            .O(N__21266),
            .I(N__21263));
    LocalMux I__2474 (
            .O(N__21263),
            .I(N__21260));
    Odrv4 I__2473 (
            .O(N__21260),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ));
    InMux I__2472 (
            .O(N__21257),
            .I(N__21254));
    LocalMux I__2471 (
            .O(N__21254),
            .I(N__21250));
    InMux I__2470 (
            .O(N__21253),
            .I(N__21247));
    Span4Mux_h I__2469 (
            .O(N__21250),
            .I(N__21241));
    LocalMux I__2468 (
            .O(N__21247),
            .I(N__21241));
    InMux I__2467 (
            .O(N__21246),
            .I(N__21238));
    Span4Mux_v I__2466 (
            .O(N__21241),
            .I(N__21235));
    LocalMux I__2465 (
            .O(N__21238),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    Odrv4 I__2464 (
            .O(N__21235),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    CascadeMux I__2463 (
            .O(N__21230),
            .I(N__21227));
    InMux I__2462 (
            .O(N__21227),
            .I(N__21224));
    LocalMux I__2461 (
            .O(N__21224),
            .I(N__21221));
    Span4Mux_h I__2460 (
            .O(N__21221),
            .I(N__21217));
    InMux I__2459 (
            .O(N__21220),
            .I(N__21214));
    Odrv4 I__2458 (
            .O(N__21217),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ));
    LocalMux I__2457 (
            .O(N__21214),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ));
    CascadeMux I__2456 (
            .O(N__21209),
            .I(N__21205));
    CascadeMux I__2455 (
            .O(N__21208),
            .I(N__21198));
    InMux I__2454 (
            .O(N__21205),
            .I(N__21194));
    InMux I__2453 (
            .O(N__21204),
            .I(N__21191));
    InMux I__2452 (
            .O(N__21203),
            .I(N__21186));
    InMux I__2451 (
            .O(N__21202),
            .I(N__21186));
    InMux I__2450 (
            .O(N__21201),
            .I(N__21183));
    InMux I__2449 (
            .O(N__21198),
            .I(N__21180));
    InMux I__2448 (
            .O(N__21197),
            .I(N__21177));
    LocalMux I__2447 (
            .O(N__21194),
            .I(N__21173));
    LocalMux I__2446 (
            .O(N__21191),
            .I(N__21170));
    LocalMux I__2445 (
            .O(N__21186),
            .I(N__21164));
    LocalMux I__2444 (
            .O(N__21183),
            .I(N__21157));
    LocalMux I__2443 (
            .O(N__21180),
            .I(N__21157));
    LocalMux I__2442 (
            .O(N__21177),
            .I(N__21157));
    InMux I__2441 (
            .O(N__21176),
            .I(N__21154));
    Span4Mux_v I__2440 (
            .O(N__21173),
            .I(N__21151));
    Span4Mux_v I__2439 (
            .O(N__21170),
            .I(N__21148));
    InMux I__2438 (
            .O(N__21169),
            .I(N__21145));
    InMux I__2437 (
            .O(N__21168),
            .I(N__21142));
    InMux I__2436 (
            .O(N__21167),
            .I(N__21139));
    Span4Mux_s2_h I__2435 (
            .O(N__21164),
            .I(N__21132));
    Span4Mux_h I__2434 (
            .O(N__21157),
            .I(N__21132));
    LocalMux I__2433 (
            .O(N__21154),
            .I(N__21132));
    Odrv4 I__2432 (
            .O(N__21151),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    Odrv4 I__2431 (
            .O(N__21148),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    LocalMux I__2430 (
            .O(N__21145),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    LocalMux I__2429 (
            .O(N__21142),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    LocalMux I__2428 (
            .O(N__21139),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    Odrv4 I__2427 (
            .O(N__21132),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    InMux I__2426 (
            .O(N__21119),
            .I(N__21116));
    LocalMux I__2425 (
            .O(N__21116),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_3 ));
    InMux I__2424 (
            .O(N__21113),
            .I(N__21108));
    InMux I__2423 (
            .O(N__21112),
            .I(N__21105));
    InMux I__2422 (
            .O(N__21111),
            .I(N__21102));
    LocalMux I__2421 (
            .O(N__21108),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__2420 (
            .O(N__21105),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__2419 (
            .O(N__21102),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    InMux I__2418 (
            .O(N__21095),
            .I(\pwm_generator_inst.counter_cry_2 ));
    InMux I__2417 (
            .O(N__21092),
            .I(N__21087));
    InMux I__2416 (
            .O(N__21091),
            .I(N__21084));
    InMux I__2415 (
            .O(N__21090),
            .I(N__21081));
    LocalMux I__2414 (
            .O(N__21087),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__2413 (
            .O(N__21084),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__2412 (
            .O(N__21081),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    InMux I__2411 (
            .O(N__21074),
            .I(\pwm_generator_inst.counter_cry_3 ));
    InMux I__2410 (
            .O(N__21071),
            .I(N__21066));
    InMux I__2409 (
            .O(N__21070),
            .I(N__21063));
    InMux I__2408 (
            .O(N__21069),
            .I(N__21060));
    LocalMux I__2407 (
            .O(N__21066),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__2406 (
            .O(N__21063),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__2405 (
            .O(N__21060),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    InMux I__2404 (
            .O(N__21053),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__2403 (
            .O(N__21050),
            .I(N__21045));
    InMux I__2402 (
            .O(N__21049),
            .I(N__21042));
    InMux I__2401 (
            .O(N__21048),
            .I(N__21039));
    LocalMux I__2400 (
            .O(N__21045),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__2399 (
            .O(N__21042),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__2398 (
            .O(N__21039),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    InMux I__2397 (
            .O(N__21032),
            .I(\pwm_generator_inst.counter_cry_5 ));
    InMux I__2396 (
            .O(N__21029),
            .I(N__21024));
    InMux I__2395 (
            .O(N__21028),
            .I(N__21021));
    InMux I__2394 (
            .O(N__21027),
            .I(N__21018));
    LocalMux I__2393 (
            .O(N__21024),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__2392 (
            .O(N__21021),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__2391 (
            .O(N__21018),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    InMux I__2390 (
            .O(N__21011),
            .I(\pwm_generator_inst.counter_cry_6 ));
    InMux I__2389 (
            .O(N__21008),
            .I(N__21003));
    InMux I__2388 (
            .O(N__21007),
            .I(N__21000));
    InMux I__2387 (
            .O(N__21006),
            .I(N__20997));
    LocalMux I__2386 (
            .O(N__21003),
            .I(N__20994));
    LocalMux I__2385 (
            .O(N__21000),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__2384 (
            .O(N__20997),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    Odrv4 I__2383 (
            .O(N__20994),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    InMux I__2382 (
            .O(N__20987),
            .I(bfn_4_14_0_));
    InMux I__2381 (
            .O(N__20984),
            .I(N__20970));
    InMux I__2380 (
            .O(N__20983),
            .I(N__20970));
    InMux I__2379 (
            .O(N__20982),
            .I(N__20970));
    InMux I__2378 (
            .O(N__20981),
            .I(N__20970));
    InMux I__2377 (
            .O(N__20980),
            .I(N__20961));
    InMux I__2376 (
            .O(N__20979),
            .I(N__20961));
    LocalMux I__2375 (
            .O(N__20970),
            .I(N__20958));
    InMux I__2374 (
            .O(N__20969),
            .I(N__20949));
    InMux I__2373 (
            .O(N__20968),
            .I(N__20949));
    InMux I__2372 (
            .O(N__20967),
            .I(N__20949));
    InMux I__2371 (
            .O(N__20966),
            .I(N__20949));
    LocalMux I__2370 (
            .O(N__20961),
            .I(N__20946));
    Odrv4 I__2369 (
            .O(N__20958),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__2368 (
            .O(N__20949),
            .I(\pwm_generator_inst.un1_counter_0 ));
    Odrv4 I__2367 (
            .O(N__20946),
            .I(\pwm_generator_inst.un1_counter_0 ));
    InMux I__2366 (
            .O(N__20939),
            .I(\pwm_generator_inst.counter_cry_8 ));
    InMux I__2365 (
            .O(N__20936),
            .I(N__20931));
    InMux I__2364 (
            .O(N__20935),
            .I(N__20928));
    InMux I__2363 (
            .O(N__20934),
            .I(N__20925));
    LocalMux I__2362 (
            .O(N__20931),
            .I(N__20922));
    LocalMux I__2361 (
            .O(N__20928),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__2360 (
            .O(N__20925),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    Odrv4 I__2359 (
            .O(N__20922),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    CascadeMux I__2358 (
            .O(N__20915),
            .I(N__20912));
    InMux I__2357 (
            .O(N__20912),
            .I(N__20909));
    LocalMux I__2356 (
            .O(N__20909),
            .I(N__20906));
    Odrv4 I__2355 (
            .O(N__20906),
            .I(\pwm_generator_inst.thresholdZ0Z_2 ));
    InMux I__2354 (
            .O(N__20903),
            .I(N__20900));
    LocalMux I__2353 (
            .O(N__20900),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ));
    InMux I__2352 (
            .O(N__20897),
            .I(N__20894));
    LocalMux I__2351 (
            .O(N__20894),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ));
    CascadeMux I__2350 (
            .O(N__20891),
            .I(\pwm_generator_inst.un1_counterlto2_0_cascade_ ));
    CascadeMux I__2349 (
            .O(N__20888),
            .I(\pwm_generator_inst.un1_counterlto9_2_cascade_ ));
    InMux I__2348 (
            .O(N__20885),
            .I(N__20882));
    LocalMux I__2347 (
            .O(N__20882),
            .I(\pwm_generator_inst.un1_counterlt9 ));
    InMux I__2346 (
            .O(N__20879),
            .I(N__20874));
    InMux I__2345 (
            .O(N__20878),
            .I(N__20871));
    InMux I__2344 (
            .O(N__20877),
            .I(N__20868));
    LocalMux I__2343 (
            .O(N__20874),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__2342 (
            .O(N__20871),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__2341 (
            .O(N__20868),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__2340 (
            .O(N__20861),
            .I(bfn_4_13_0_));
    InMux I__2339 (
            .O(N__20858),
            .I(N__20853));
    InMux I__2338 (
            .O(N__20857),
            .I(N__20850));
    InMux I__2337 (
            .O(N__20856),
            .I(N__20847));
    LocalMux I__2336 (
            .O(N__20853),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__2335 (
            .O(N__20850),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__2334 (
            .O(N__20847),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    InMux I__2333 (
            .O(N__20840),
            .I(\pwm_generator_inst.counter_cry_0 ));
    InMux I__2332 (
            .O(N__20837),
            .I(N__20832));
    InMux I__2331 (
            .O(N__20836),
            .I(N__20829));
    InMux I__2330 (
            .O(N__20835),
            .I(N__20826));
    LocalMux I__2329 (
            .O(N__20832),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__2328 (
            .O(N__20829),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__2327 (
            .O(N__20826),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    InMux I__2326 (
            .O(N__20819),
            .I(\pwm_generator_inst.counter_cry_1 ));
    CascadeMux I__2325 (
            .O(N__20816),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ));
    InMux I__2324 (
            .O(N__20813),
            .I(N__20810));
    LocalMux I__2323 (
            .O(N__20810),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ));
    InMux I__2322 (
            .O(N__20807),
            .I(N__20804));
    LocalMux I__2321 (
            .O(N__20804),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ));
    InMux I__2320 (
            .O(N__20801),
            .I(N__20798));
    LocalMux I__2319 (
            .O(N__20798),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    CascadeMux I__2318 (
            .O(N__20795),
            .I(N__20792));
    InMux I__2317 (
            .O(N__20792),
            .I(N__20789));
    LocalMux I__2316 (
            .O(N__20789),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ));
    CascadeMux I__2315 (
            .O(N__20786),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ));
    InMux I__2314 (
            .O(N__20783),
            .I(N__20780));
    LocalMux I__2313 (
            .O(N__20780),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ));
    InMux I__2312 (
            .O(N__20777),
            .I(N__20774));
    LocalMux I__2311 (
            .O(N__20774),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9 ));
    InMux I__2310 (
            .O(N__20771),
            .I(N__20768));
    LocalMux I__2309 (
            .O(N__20768),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ));
    InMux I__2308 (
            .O(N__20765),
            .I(N__20762));
    LocalMux I__2307 (
            .O(N__20762),
            .I(N__20759));
    Odrv4 I__2306 (
            .O(N__20759),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_5 ));
    InMux I__2305 (
            .O(N__20756),
            .I(N__20753));
    LocalMux I__2304 (
            .O(N__20753),
            .I(N__20750));
    Span12Mux_s9_v I__2303 (
            .O(N__20750),
            .I(N__20747));
    Odrv12 I__2302 (
            .O(N__20747),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ));
    InMux I__2301 (
            .O(N__20744),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_4 ));
    InMux I__2300 (
            .O(N__20741),
            .I(N__20738));
    LocalMux I__2299 (
            .O(N__20738),
            .I(N__20735));
    Odrv4 I__2298 (
            .O(N__20735),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_6 ));
    InMux I__2297 (
            .O(N__20732),
            .I(N__20729));
    LocalMux I__2296 (
            .O(N__20729),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ));
    InMux I__2295 (
            .O(N__20726),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_5 ));
    InMux I__2294 (
            .O(N__20723),
            .I(N__20720));
    LocalMux I__2293 (
            .O(N__20720),
            .I(N__20717));
    Odrv4 I__2292 (
            .O(N__20717),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_7 ));
    InMux I__2291 (
            .O(N__20714),
            .I(N__20711));
    LocalMux I__2290 (
            .O(N__20711),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ));
    InMux I__2289 (
            .O(N__20708),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_6 ));
    InMux I__2288 (
            .O(N__20705),
            .I(bfn_3_18_0_));
    InMux I__2287 (
            .O(N__20702),
            .I(N__20699));
    LocalMux I__2286 (
            .O(N__20699),
            .I(N__20696));
    Span4Mux_v I__2285 (
            .O(N__20696),
            .I(N__20693));
    Odrv4 I__2284 (
            .O(N__20693),
            .I(\pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ));
    InMux I__2283 (
            .O(N__20690),
            .I(N__20687));
    LocalMux I__2282 (
            .O(N__20687),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ));
    InMux I__2281 (
            .O(N__20684),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_8 ));
    InMux I__2280 (
            .O(N__20681),
            .I(N__20678));
    LocalMux I__2279 (
            .O(N__20678),
            .I(N__20675));
    Span4Mux_v I__2278 (
            .O(N__20675),
            .I(N__20671));
    InMux I__2277 (
            .O(N__20674),
            .I(N__20668));
    Odrv4 I__2276 (
            .O(N__20671),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ));
    LocalMux I__2275 (
            .O(N__20668),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ));
    CascadeMux I__2274 (
            .O(N__20663),
            .I(N__20659));
    InMux I__2273 (
            .O(N__20662),
            .I(N__20655));
    InMux I__2272 (
            .O(N__20659),
            .I(N__20652));
    InMux I__2271 (
            .O(N__20658),
            .I(N__20649));
    LocalMux I__2270 (
            .O(N__20655),
            .I(N__20644));
    LocalMux I__2269 (
            .O(N__20652),
            .I(N__20644));
    LocalMux I__2268 (
            .O(N__20649),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    Odrv4 I__2267 (
            .O(N__20644),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    InMux I__2266 (
            .O(N__20639),
            .I(N__20636));
    LocalMux I__2265 (
            .O(N__20636),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ));
    InMux I__2264 (
            .O(N__20633),
            .I(N__20630));
    LocalMux I__2263 (
            .O(N__20630),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_8 ));
    InMux I__2262 (
            .O(N__20627),
            .I(N__20624));
    LocalMux I__2261 (
            .O(N__20624),
            .I(N__20621));
    Glb2LocalMux I__2260 (
            .O(N__20621),
            .I(N__20618));
    GlobalMux I__2259 (
            .O(N__20618),
            .I(clk_12mhz));
    IoInMux I__2258 (
            .O(N__20615),
            .I(N__20612));
    LocalMux I__2257 (
            .O(N__20612),
            .I(N__20609));
    Span4Mux_s0_v I__2256 (
            .O(N__20609),
            .I(N__20606));
    Sp12to4 I__2255 (
            .O(N__20606),
            .I(N__20603));
    Odrv12 I__2254 (
            .O(N__20603),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__2253 (
            .O(N__20600),
            .I(N__20597));
    LocalMux I__2252 (
            .O(N__20597),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ));
    InMux I__2251 (
            .O(N__20594),
            .I(N__20591));
    LocalMux I__2250 (
            .O(N__20591),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_7 ));
    InMux I__2249 (
            .O(N__20588),
            .I(N__20585));
    LocalMux I__2248 (
            .O(N__20585),
            .I(N__20582));
    Odrv12 I__2247 (
            .O(N__20582),
            .I(\pwm_generator_inst.thresholdZ0Z_7 ));
    InMux I__2246 (
            .O(N__20579),
            .I(N__20576));
    LocalMux I__2245 (
            .O(N__20576),
            .I(N__20573));
    Odrv4 I__2244 (
            .O(N__20573),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_4 ));
    InMux I__2243 (
            .O(N__20570),
            .I(N__20567));
    LocalMux I__2242 (
            .O(N__20567),
            .I(N__20564));
    Odrv12 I__2241 (
            .O(N__20564),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_1 ));
    InMux I__2240 (
            .O(N__20561),
            .I(N__20558));
    LocalMux I__2239 (
            .O(N__20558),
            .I(N__20555));
    Odrv4 I__2238 (
            .O(N__20555),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_0 ));
    InMux I__2237 (
            .O(N__20552),
            .I(N__20549));
    LocalMux I__2236 (
            .O(N__20549),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ));
    InMux I__2235 (
            .O(N__20546),
            .I(N__20543));
    LocalMux I__2234 (
            .O(N__20543),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_1 ));
    InMux I__2233 (
            .O(N__20540),
            .I(N__20537));
    LocalMux I__2232 (
            .O(N__20537),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ));
    InMux I__2231 (
            .O(N__20534),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_0 ));
    InMux I__2230 (
            .O(N__20531),
            .I(N__20528));
    LocalMux I__2229 (
            .O(N__20528),
            .I(N__20525));
    Odrv4 I__2228 (
            .O(N__20525),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_2 ));
    InMux I__2227 (
            .O(N__20522),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_1 ));
    InMux I__2226 (
            .O(N__20519),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_2 ));
    InMux I__2225 (
            .O(N__20516),
            .I(N__20513));
    LocalMux I__2224 (
            .O(N__20513),
            .I(N__20510));
    Odrv4 I__2223 (
            .O(N__20510),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_4 ));
    InMux I__2222 (
            .O(N__20507),
            .I(N__20504));
    LocalMux I__2221 (
            .O(N__20504),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ));
    InMux I__2220 (
            .O(N__20501),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_3 ));
    CascadeMux I__2219 (
            .O(N__20498),
            .I(N__20495));
    InMux I__2218 (
            .O(N__20495),
            .I(N__20492));
    LocalMux I__2217 (
            .O(N__20492),
            .I(N__20489));
    Odrv4 I__2216 (
            .O(N__20489),
            .I(\pwm_generator_inst.thresholdZ0Z_4 ));
    InMux I__2215 (
            .O(N__20486),
            .I(N__20483));
    LocalMux I__2214 (
            .O(N__20483),
            .I(N__20480));
    Odrv4 I__2213 (
            .O(N__20480),
            .I(\pwm_generator_inst.thresholdZ0Z_6 ));
    InMux I__2212 (
            .O(N__20477),
            .I(N__20473));
    InMux I__2211 (
            .O(N__20476),
            .I(N__20470));
    LocalMux I__2210 (
            .O(N__20473),
            .I(N__20467));
    LocalMux I__2209 (
            .O(N__20470),
            .I(N__20464));
    Span4Mux_v I__2208 (
            .O(N__20467),
            .I(N__20461));
    Span4Mux_v I__2207 (
            .O(N__20464),
            .I(N__20458));
    Odrv4 I__2206 (
            .O(N__20461),
            .I(\pwm_generator_inst.O_10 ));
    Odrv4 I__2205 (
            .O(N__20458),
            .I(\pwm_generator_inst.O_10 ));
    InMux I__2204 (
            .O(N__20453),
            .I(N__20450));
    LocalMux I__2203 (
            .O(N__20450),
            .I(N__20446));
    InMux I__2202 (
            .O(N__20449),
            .I(N__20442));
    Span4Mux_h I__2201 (
            .O(N__20446),
            .I(N__20439));
    InMux I__2200 (
            .O(N__20445),
            .I(N__20436));
    LocalMux I__2199 (
            .O(N__20442),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    Odrv4 I__2198 (
            .O(N__20439),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    LocalMux I__2197 (
            .O(N__20436),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    CascadeMux I__2196 (
            .O(N__20429),
            .I(N__20426));
    InMux I__2195 (
            .O(N__20426),
            .I(N__20423));
    LocalMux I__2194 (
            .O(N__20423),
            .I(N__20420));
    Odrv4 I__2193 (
            .O(N__20420),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ));
    InMux I__2192 (
            .O(N__20417),
            .I(N__20414));
    LocalMux I__2191 (
            .O(N__20414),
            .I(N__20411));
    Odrv4 I__2190 (
            .O(N__20411),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_0 ));
    InMux I__2189 (
            .O(N__20408),
            .I(N__20405));
    LocalMux I__2188 (
            .O(N__20405),
            .I(N__20402));
    Odrv4 I__2187 (
            .O(N__20402),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_6 ));
    InMux I__2186 (
            .O(N__20399),
            .I(N__20396));
    LocalMux I__2185 (
            .O(N__20396),
            .I(\pwm_generator_inst.counter_i_4 ));
    CascadeMux I__2184 (
            .O(N__20393),
            .I(N__20390));
    InMux I__2183 (
            .O(N__20390),
            .I(N__20387));
    LocalMux I__2182 (
            .O(N__20387),
            .I(N__20384));
    Span4Mux_h I__2181 (
            .O(N__20384),
            .I(N__20381));
    Odrv4 I__2180 (
            .O(N__20381),
            .I(\pwm_generator_inst.thresholdZ0Z_5 ));
    InMux I__2179 (
            .O(N__20378),
            .I(N__20375));
    LocalMux I__2178 (
            .O(N__20375),
            .I(\pwm_generator_inst.counter_i_5 ));
    CascadeMux I__2177 (
            .O(N__20372),
            .I(N__20369));
    InMux I__2176 (
            .O(N__20369),
            .I(N__20366));
    LocalMux I__2175 (
            .O(N__20366),
            .I(\pwm_generator_inst.counter_i_6 ));
    CascadeMux I__2174 (
            .O(N__20363),
            .I(N__20360));
    InMux I__2173 (
            .O(N__20360),
            .I(N__20357));
    LocalMux I__2172 (
            .O(N__20357),
            .I(\pwm_generator_inst.counter_i_7 ));
    CascadeMux I__2171 (
            .O(N__20354),
            .I(N__20351));
    InMux I__2170 (
            .O(N__20351),
            .I(N__20348));
    LocalMux I__2169 (
            .O(N__20348),
            .I(\pwm_generator_inst.counter_i_8 ));
    CascadeMux I__2168 (
            .O(N__20345),
            .I(N__20342));
    InMux I__2167 (
            .O(N__20342),
            .I(N__20339));
    LocalMux I__2166 (
            .O(N__20339),
            .I(\pwm_generator_inst.counter_i_9 ));
    InMux I__2165 (
            .O(N__20336),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    IoInMux I__2164 (
            .O(N__20333),
            .I(N__20330));
    LocalMux I__2163 (
            .O(N__20330),
            .I(N__20327));
    Span4Mux_s2_v I__2162 (
            .O(N__20327),
            .I(N__20324));
    Sp12to4 I__2161 (
            .O(N__20324),
            .I(N__20321));
    Span12Mux_s10_h I__2160 (
            .O(N__20321),
            .I(N__20318));
    Span12Mux_h I__2159 (
            .O(N__20318),
            .I(N__20315));
    Odrv12 I__2158 (
            .O(N__20315),
            .I(pwm_output_c));
    InMux I__2157 (
            .O(N__20312),
            .I(N__20309));
    LocalMux I__2156 (
            .O(N__20309),
            .I(N__20306));
    Odrv4 I__2155 (
            .O(N__20306),
            .I(\pwm_generator_inst.thresholdZ0Z_0 ));
    InMux I__2154 (
            .O(N__20303),
            .I(N__20300));
    LocalMux I__2153 (
            .O(N__20300),
            .I(N__20297));
    Odrv4 I__2152 (
            .O(N__20297),
            .I(\pwm_generator_inst.thresholdZ0Z_1 ));
    InMux I__2151 (
            .O(N__20294),
            .I(N__20291));
    LocalMux I__2150 (
            .O(N__20291),
            .I(N__20287));
    InMux I__2149 (
            .O(N__20290),
            .I(N__20283));
    Span4Mux_h I__2148 (
            .O(N__20287),
            .I(N__20280));
    InMux I__2147 (
            .O(N__20286),
            .I(N__20277));
    LocalMux I__2146 (
            .O(N__20283),
            .I(pwm_duty_input_5));
    Odrv4 I__2145 (
            .O(N__20280),
            .I(pwm_duty_input_5));
    LocalMux I__2144 (
            .O(N__20277),
            .I(pwm_duty_input_5));
    InMux I__2143 (
            .O(N__20270),
            .I(N__20267));
    LocalMux I__2142 (
            .O(N__20267),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0 ));
    CascadeMux I__2141 (
            .O(N__20264),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_ ));
    CascadeMux I__2140 (
            .O(N__20261),
            .I(N__20254));
    InMux I__2139 (
            .O(N__20260),
            .I(N__20250));
    InMux I__2138 (
            .O(N__20259),
            .I(N__20239));
    InMux I__2137 (
            .O(N__20258),
            .I(N__20239));
    InMux I__2136 (
            .O(N__20257),
            .I(N__20239));
    InMux I__2135 (
            .O(N__20254),
            .I(N__20239));
    InMux I__2134 (
            .O(N__20253),
            .I(N__20239));
    LocalMux I__2133 (
            .O(N__20250),
            .I(N__20236));
    LocalMux I__2132 (
            .O(N__20239),
            .I(N__20228));
    Span4Mux_v I__2131 (
            .O(N__20236),
            .I(N__20228));
    InMux I__2130 (
            .O(N__20235),
            .I(N__20225));
    InMux I__2129 (
            .O(N__20234),
            .I(N__20220));
    InMux I__2128 (
            .O(N__20233),
            .I(N__20220));
    Odrv4 I__2127 (
            .O(N__20228),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    LocalMux I__2126 (
            .O(N__20225),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    LocalMux I__2125 (
            .O(N__20220),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    InMux I__2124 (
            .O(N__20213),
            .I(N__20210));
    LocalMux I__2123 (
            .O(N__20210),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ));
    CascadeMux I__2122 (
            .O(N__20207),
            .I(N__20201));
    CascadeMux I__2121 (
            .O(N__20206),
            .I(N__20198));
    CascadeMux I__2120 (
            .O(N__20205),
            .I(N__20195));
    CascadeMux I__2119 (
            .O(N__20204),
            .I(N__20192));
    InMux I__2118 (
            .O(N__20201),
            .I(N__20179));
    InMux I__2117 (
            .O(N__20198),
            .I(N__20179));
    InMux I__2116 (
            .O(N__20195),
            .I(N__20179));
    InMux I__2115 (
            .O(N__20192),
            .I(N__20179));
    InMux I__2114 (
            .O(N__20191),
            .I(N__20179));
    InMux I__2113 (
            .O(N__20190),
            .I(N__20176));
    LocalMux I__2112 (
            .O(N__20179),
            .I(N__20173));
    LocalMux I__2111 (
            .O(N__20176),
            .I(N__20169));
    Span4Mux_s3_h I__2110 (
            .O(N__20173),
            .I(N__20166));
    InMux I__2109 (
            .O(N__20172),
            .I(N__20163));
    Odrv4 I__2108 (
            .O(N__20169),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    Odrv4 I__2107 (
            .O(N__20166),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    LocalMux I__2106 (
            .O(N__20163),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    CascadeMux I__2105 (
            .O(N__20156),
            .I(N__20153));
    InMux I__2104 (
            .O(N__20153),
            .I(N__20150));
    LocalMux I__2103 (
            .O(N__20150),
            .I(\pwm_generator_inst.counter_i_0 ));
    CascadeMux I__2102 (
            .O(N__20147),
            .I(N__20144));
    InMux I__2101 (
            .O(N__20144),
            .I(N__20141));
    LocalMux I__2100 (
            .O(N__20141),
            .I(N__20138));
    Odrv4 I__2099 (
            .O(N__20138),
            .I(\pwm_generator_inst.counter_i_1 ));
    InMux I__2098 (
            .O(N__20135),
            .I(N__20132));
    LocalMux I__2097 (
            .O(N__20132),
            .I(\pwm_generator_inst.counter_i_2 ));
    CascadeMux I__2096 (
            .O(N__20129),
            .I(N__20126));
    InMux I__2095 (
            .O(N__20126),
            .I(N__20123));
    LocalMux I__2094 (
            .O(N__20123),
            .I(\pwm_generator_inst.counter_i_3 ));
    InMux I__2093 (
            .O(N__20120),
            .I(N__20116));
    InMux I__2092 (
            .O(N__20119),
            .I(N__20113));
    LocalMux I__2091 (
            .O(N__20116),
            .I(N__20110));
    LocalMux I__2090 (
            .O(N__20113),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    Odrv4 I__2089 (
            .O(N__20110),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    InMux I__2088 (
            .O(N__20105),
            .I(N__20102));
    LocalMux I__2087 (
            .O(N__20102),
            .I(N__20099));
    Odrv4 I__2086 (
            .O(N__20099),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ));
    InMux I__2085 (
            .O(N__20096),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ));
    InMux I__2084 (
            .O(N__20093),
            .I(N__20089));
    InMux I__2083 (
            .O(N__20092),
            .I(N__20086));
    LocalMux I__2082 (
            .O(N__20089),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    LocalMux I__2081 (
            .O(N__20086),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    InMux I__2080 (
            .O(N__20081),
            .I(N__20078));
    LocalMux I__2079 (
            .O(N__20078),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ));
    InMux I__2078 (
            .O(N__20075),
            .I(bfn_2_18_0_));
    InMux I__2077 (
            .O(N__20072),
            .I(N__20068));
    InMux I__2076 (
            .O(N__20071),
            .I(N__20065));
    LocalMux I__2075 (
            .O(N__20068),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    LocalMux I__2074 (
            .O(N__20065),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    InMux I__2073 (
            .O(N__20060),
            .I(N__20057));
    LocalMux I__2072 (
            .O(N__20057),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ));
    InMux I__2071 (
            .O(N__20054),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ));
    InMux I__2070 (
            .O(N__20051),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ));
    InMux I__2069 (
            .O(N__20048),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_18 ));
    InMux I__2068 (
            .O(N__20045),
            .I(N__20042));
    LocalMux I__2067 (
            .O(N__20042),
            .I(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ));
    InMux I__2066 (
            .O(N__20039),
            .I(N__20036));
    LocalMux I__2065 (
            .O(N__20036),
            .I(N__20033));
    Odrv4 I__2064 (
            .O(N__20033),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_5 ));
    InMux I__2063 (
            .O(N__20030),
            .I(N__20027));
    LocalMux I__2062 (
            .O(N__20027),
            .I(N__20022));
    InMux I__2061 (
            .O(N__20026),
            .I(N__20019));
    InMux I__2060 (
            .O(N__20025),
            .I(N__20016));
    Span4Mux_h I__2059 (
            .O(N__20022),
            .I(N__20013));
    LocalMux I__2058 (
            .O(N__20019),
            .I(N__20010));
    LocalMux I__2057 (
            .O(N__20016),
            .I(N__20007));
    Odrv4 I__2056 (
            .O(N__20013),
            .I(pwm_duty_input_8));
    Odrv4 I__2055 (
            .O(N__20010),
            .I(pwm_duty_input_8));
    Odrv4 I__2054 (
            .O(N__20007),
            .I(pwm_duty_input_8));
    InMux I__2053 (
            .O(N__20000),
            .I(N__19995));
    InMux I__2052 (
            .O(N__19999),
            .I(N__19992));
    InMux I__2051 (
            .O(N__19998),
            .I(N__19989));
    LocalMux I__2050 (
            .O(N__19995),
            .I(N__19986));
    LocalMux I__2049 (
            .O(N__19992),
            .I(N__19983));
    LocalMux I__2048 (
            .O(N__19989),
            .I(N__19980));
    Span4Mux_h I__2047 (
            .O(N__19986),
            .I(N__19977));
    Span4Mux_h I__2046 (
            .O(N__19983),
            .I(N__19974));
    Span4Mux_s1_h I__2045 (
            .O(N__19980),
            .I(N__19971));
    Odrv4 I__2044 (
            .O(N__19977),
            .I(pwm_duty_input_9));
    Odrv4 I__2043 (
            .O(N__19974),
            .I(pwm_duty_input_9));
    Odrv4 I__2042 (
            .O(N__19971),
            .I(pwm_duty_input_9));
    CascadeMux I__2041 (
            .O(N__19964),
            .I(N__19960));
    CascadeMux I__2040 (
            .O(N__19963),
            .I(N__19957));
    InMux I__2039 (
            .O(N__19960),
            .I(N__19953));
    InMux I__2038 (
            .O(N__19957),
            .I(N__19950));
    InMux I__2037 (
            .O(N__19956),
            .I(N__19947));
    LocalMux I__2036 (
            .O(N__19953),
            .I(N__19942));
    LocalMux I__2035 (
            .O(N__19950),
            .I(N__19942));
    LocalMux I__2034 (
            .O(N__19947),
            .I(N__19939));
    Span4Mux_v I__2033 (
            .O(N__19942),
            .I(N__19936));
    Span4Mux_s1_h I__2032 (
            .O(N__19939),
            .I(N__19933));
    Odrv4 I__2031 (
            .O(N__19936),
            .I(pwm_duty_input_6));
    Odrv4 I__2030 (
            .O(N__19933),
            .I(pwm_duty_input_6));
    InMux I__2029 (
            .O(N__19928),
            .I(N__19925));
    LocalMux I__2028 (
            .O(N__19925),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ));
    InMux I__2027 (
            .O(N__19922),
            .I(N__19918));
    InMux I__2026 (
            .O(N__19921),
            .I(N__19914));
    LocalMux I__2025 (
            .O(N__19918),
            .I(N__19911));
    InMux I__2024 (
            .O(N__19917),
            .I(N__19908));
    LocalMux I__2023 (
            .O(N__19914),
            .I(N__19905));
    Span4Mux_h I__2022 (
            .O(N__19911),
            .I(N__19900));
    LocalMux I__2021 (
            .O(N__19908),
            .I(N__19900));
    Odrv12 I__2020 (
            .O(N__19905),
            .I(pwm_duty_input_7));
    Odrv4 I__2019 (
            .O(N__19900),
            .I(pwm_duty_input_7));
    InMux I__2018 (
            .O(N__19895),
            .I(N__19892));
    LocalMux I__2017 (
            .O(N__19892),
            .I(N__19889));
    Span4Mux_h I__2016 (
            .O(N__19889),
            .I(N__19886));
    Span4Mux_v I__2015 (
            .O(N__19886),
            .I(N__19883));
    Odrv4 I__2014 (
            .O(N__19883),
            .I(\pwm_generator_inst.O_7 ));
    InMux I__2013 (
            .O(N__19880),
            .I(N__19877));
    LocalMux I__2012 (
            .O(N__19877),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_7 ));
    InMux I__2011 (
            .O(N__19874),
            .I(N__19871));
    LocalMux I__2010 (
            .O(N__19871),
            .I(N__19868));
    Span4Mux_h I__2009 (
            .O(N__19868),
            .I(N__19865));
    Span4Mux_v I__2008 (
            .O(N__19865),
            .I(N__19862));
    Odrv4 I__2007 (
            .O(N__19862),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__2006 (
            .O(N__19859),
            .I(N__19856));
    LocalMux I__2005 (
            .O(N__19856),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_8 ));
    InMux I__2004 (
            .O(N__19853),
            .I(N__19850));
    LocalMux I__2003 (
            .O(N__19850),
            .I(N__19847));
    Span4Mux_h I__2002 (
            .O(N__19847),
            .I(N__19844));
    Span4Mux_v I__2001 (
            .O(N__19844),
            .I(N__19841));
    Odrv4 I__2000 (
            .O(N__19841),
            .I(\pwm_generator_inst.O_9 ));
    InMux I__1999 (
            .O(N__19838),
            .I(N__19835));
    LocalMux I__1998 (
            .O(N__19835),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_9 ));
    InMux I__1997 (
            .O(N__19832),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ));
    InMux I__1996 (
            .O(N__19829),
            .I(N__19826));
    LocalMux I__1995 (
            .O(N__19826),
            .I(N__19823));
    Span4Mux_v I__1994 (
            .O(N__19823),
            .I(N__19819));
    InMux I__1993 (
            .O(N__19822),
            .I(N__19816));
    Span4Mux_v I__1992 (
            .O(N__19819),
            .I(N__19813));
    LocalMux I__1991 (
            .O(N__19816),
            .I(N__19810));
    Odrv4 I__1990 (
            .O(N__19813),
            .I(\pwm_generator_inst.un3_threshold_acc ));
    Odrv4 I__1989 (
            .O(N__19810),
            .I(\pwm_generator_inst.un3_threshold_acc ));
    InMux I__1988 (
            .O(N__19805),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ));
    InMux I__1987 (
            .O(N__19802),
            .I(N__19797));
    InMux I__1986 (
            .O(N__19801),
            .I(N__19794));
    InMux I__1985 (
            .O(N__19800),
            .I(N__19791));
    LocalMux I__1984 (
            .O(N__19797),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    LocalMux I__1983 (
            .O(N__19794),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    LocalMux I__1982 (
            .O(N__19791),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    InMux I__1981 (
            .O(N__19784),
            .I(N__19781));
    LocalMux I__1980 (
            .O(N__19781),
            .I(N__19778));
    Odrv4 I__1979 (
            .O(N__19778),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ));
    InMux I__1978 (
            .O(N__19775),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ));
    InMux I__1977 (
            .O(N__19772),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ));
    InMux I__1976 (
            .O(N__19769),
            .I(N__19765));
    InMux I__1975 (
            .O(N__19768),
            .I(N__19762));
    LocalMux I__1974 (
            .O(N__19765),
            .I(N__19759));
    LocalMux I__1973 (
            .O(N__19762),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    Odrv4 I__1972 (
            .O(N__19759),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    InMux I__1971 (
            .O(N__19754),
            .I(N__19751));
    LocalMux I__1970 (
            .O(N__19751),
            .I(N__19748));
    Span4Mux_h I__1969 (
            .O(N__19748),
            .I(N__19745));
    Odrv4 I__1968 (
            .O(N__19745),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ));
    InMux I__1967 (
            .O(N__19742),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ));
    InMux I__1966 (
            .O(N__19739),
            .I(N__19733));
    InMux I__1965 (
            .O(N__19738),
            .I(N__19733));
    LocalMux I__1964 (
            .O(N__19733),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ));
    CascadeMux I__1963 (
            .O(N__19730),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14_cascade_ ));
    InMux I__1962 (
            .O(N__19727),
            .I(N__19724));
    LocalMux I__1961 (
            .O(N__19724),
            .I(N__19721));
    Span4Mux_h I__1960 (
            .O(N__19721),
            .I(N__19718));
    Span4Mux_v I__1959 (
            .O(N__19718),
            .I(N__19715));
    Odrv4 I__1958 (
            .O(N__19715),
            .I(\pwm_generator_inst.O_0 ));
    InMux I__1957 (
            .O(N__19712),
            .I(N__19709));
    LocalMux I__1956 (
            .O(N__19709),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_0 ));
    InMux I__1955 (
            .O(N__19706),
            .I(N__19703));
    LocalMux I__1954 (
            .O(N__19703),
            .I(N__19700));
    Span4Mux_h I__1953 (
            .O(N__19700),
            .I(N__19697));
    Span4Mux_v I__1952 (
            .O(N__19697),
            .I(N__19694));
    Odrv4 I__1951 (
            .O(N__19694),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__1950 (
            .O(N__19691),
            .I(N__19688));
    LocalMux I__1949 (
            .O(N__19688),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_1 ));
    InMux I__1948 (
            .O(N__19685),
            .I(N__19682));
    LocalMux I__1947 (
            .O(N__19682),
            .I(N__19679));
    Span4Mux_v I__1946 (
            .O(N__19679),
            .I(N__19676));
    Span4Mux_v I__1945 (
            .O(N__19676),
            .I(N__19673));
    Odrv4 I__1944 (
            .O(N__19673),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__1943 (
            .O(N__19670),
            .I(N__19667));
    LocalMux I__1942 (
            .O(N__19667),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_2 ));
    InMux I__1941 (
            .O(N__19664),
            .I(N__19661));
    LocalMux I__1940 (
            .O(N__19661),
            .I(N__19658));
    Span4Mux_v I__1939 (
            .O(N__19658),
            .I(N__19655));
    Span4Mux_v I__1938 (
            .O(N__19655),
            .I(N__19652));
    Odrv4 I__1937 (
            .O(N__19652),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__1936 (
            .O(N__19649),
            .I(N__19646));
    LocalMux I__1935 (
            .O(N__19646),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_3 ));
    InMux I__1934 (
            .O(N__19643),
            .I(N__19640));
    LocalMux I__1933 (
            .O(N__19640),
            .I(N__19637));
    Span4Mux_h I__1932 (
            .O(N__19637),
            .I(N__19634));
    Span4Mux_v I__1931 (
            .O(N__19634),
            .I(N__19631));
    Odrv4 I__1930 (
            .O(N__19631),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__1929 (
            .O(N__19628),
            .I(N__19625));
    LocalMux I__1928 (
            .O(N__19625),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_4 ));
    InMux I__1927 (
            .O(N__19622),
            .I(N__19619));
    LocalMux I__1926 (
            .O(N__19619),
            .I(N__19616));
    Span4Mux_h I__1925 (
            .O(N__19616),
            .I(N__19613));
    Span4Mux_v I__1924 (
            .O(N__19613),
            .I(N__19610));
    Odrv4 I__1923 (
            .O(N__19610),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__1922 (
            .O(N__19607),
            .I(N__19604));
    LocalMux I__1921 (
            .O(N__19604),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_5 ));
    InMux I__1920 (
            .O(N__19601),
            .I(N__19598));
    LocalMux I__1919 (
            .O(N__19598),
            .I(N__19595));
    Span12Mux_h I__1918 (
            .O(N__19595),
            .I(N__19592));
    Odrv12 I__1917 (
            .O(N__19592),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__1916 (
            .O(N__19589),
            .I(N__19586));
    LocalMux I__1915 (
            .O(N__19586),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_6 ));
    CascadeMux I__1914 (
            .O(N__19583),
            .I(N__19580));
    InMux I__1913 (
            .O(N__19580),
            .I(N__19577));
    LocalMux I__1912 (
            .O(N__19577),
            .I(N__19574));
    Span12Mux_v I__1911 (
            .O(N__19574),
            .I(N__19571));
    Odrv12 I__1910 (
            .O(N__19571),
            .I(\pwm_generator_inst.un2_threshold_acc_2_14 ));
    InMux I__1909 (
            .O(N__19568),
            .I(N__19565));
    LocalMux I__1908 (
            .O(N__19565),
            .I(N__19562));
    Odrv4 I__1907 (
            .O(N__19562),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ));
    InMux I__1906 (
            .O(N__19559),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ));
    InMux I__1905 (
            .O(N__19556),
            .I(N__19553));
    LocalMux I__1904 (
            .O(N__19553),
            .I(N__19550));
    Span4Mux_v I__1903 (
            .O(N__19550),
            .I(N__19547));
    Span4Mux_v I__1902 (
            .O(N__19547),
            .I(N__19544));
    Odrv4 I__1901 (
            .O(N__19544),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ));
    InMux I__1900 (
            .O(N__19541),
            .I(N__19532));
    InMux I__1899 (
            .O(N__19540),
            .I(N__19529));
    CascadeMux I__1898 (
            .O(N__19539),
            .I(N__19526));
    CascadeMux I__1897 (
            .O(N__19538),
            .I(N__19522));
    CascadeMux I__1896 (
            .O(N__19537),
            .I(N__19519));
    CascadeMux I__1895 (
            .O(N__19536),
            .I(N__19516));
    CascadeMux I__1894 (
            .O(N__19535),
            .I(N__19513));
    LocalMux I__1893 (
            .O(N__19532),
            .I(N__19510));
    LocalMux I__1892 (
            .O(N__19529),
            .I(N__19507));
    InMux I__1891 (
            .O(N__19526),
            .I(N__19498));
    InMux I__1890 (
            .O(N__19525),
            .I(N__19498));
    InMux I__1889 (
            .O(N__19522),
            .I(N__19498));
    InMux I__1888 (
            .O(N__19519),
            .I(N__19498));
    InMux I__1887 (
            .O(N__19516),
            .I(N__19493));
    InMux I__1886 (
            .O(N__19513),
            .I(N__19493));
    Span4Mux_v I__1885 (
            .O(N__19510),
            .I(N__19490));
    Span4Mux_h I__1884 (
            .O(N__19507),
            .I(N__19487));
    LocalMux I__1883 (
            .O(N__19498),
            .I(N__19482));
    LocalMux I__1882 (
            .O(N__19493),
            .I(N__19482));
    Span4Mux_v I__1881 (
            .O(N__19490),
            .I(N__19479));
    Span4Mux_v I__1880 (
            .O(N__19487),
            .I(N__19476));
    Span4Mux_h I__1879 (
            .O(N__19482),
            .I(N__19473));
    Odrv4 I__1878 (
            .O(N__19479),
            .I(\pwm_generator_inst.un2_threshold_acc_1_25 ));
    Odrv4 I__1877 (
            .O(N__19476),
            .I(\pwm_generator_inst.un2_threshold_acc_1_25 ));
    Odrv4 I__1876 (
            .O(N__19473),
            .I(\pwm_generator_inst.un2_threshold_acc_1_25 ));
    CascadeMux I__1875 (
            .O(N__19466),
            .I(N__19463));
    InMux I__1874 (
            .O(N__19463),
            .I(N__19460));
    LocalMux I__1873 (
            .O(N__19460),
            .I(N__19457));
    Odrv4 I__1872 (
            .O(N__19457),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ));
    InMux I__1871 (
            .O(N__19454),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ));
    InMux I__1870 (
            .O(N__19451),
            .I(N__19448));
    LocalMux I__1869 (
            .O(N__19448),
            .I(N__19445));
    Span4Mux_h I__1868 (
            .O(N__19445),
            .I(N__19442));
    Odrv4 I__1867 (
            .O(N__19442),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ));
    InMux I__1866 (
            .O(N__19439),
            .I(N__19436));
    LocalMux I__1865 (
            .O(N__19436),
            .I(N__19433));
    Span12Mux_v I__1864 (
            .O(N__19433),
            .I(N__19430));
    Odrv12 I__1863 (
            .O(N__19430),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ));
    InMux I__1862 (
            .O(N__19427),
            .I(bfn_2_15_0_));
    InMux I__1861 (
            .O(N__19424),
            .I(N__19420));
    InMux I__1860 (
            .O(N__19423),
            .I(N__19417));
    LocalMux I__1859 (
            .O(N__19420),
            .I(N__19414));
    LocalMux I__1858 (
            .O(N__19417),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ));
    Odrv4 I__1857 (
            .O(N__19414),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ));
    CascadeMux I__1856 (
            .O(N__19409),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_ ));
    InMux I__1855 (
            .O(N__19406),
            .I(N__19400));
    InMux I__1854 (
            .O(N__19405),
            .I(N__19400));
    LocalMux I__1853 (
            .O(N__19400),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ));
    CascadeMux I__1852 (
            .O(N__19397),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_ ));
    InMux I__1851 (
            .O(N__19394),
            .I(N__19391));
    LocalMux I__1850 (
            .O(N__19391),
            .I(N__19388));
    Span4Mux_v I__1849 (
            .O(N__19388),
            .I(N__19385));
    Odrv4 I__1848 (
            .O(N__19385),
            .I(\pwm_generator_inst.un2_threshold_acc_1_21 ));
    CascadeMux I__1847 (
            .O(N__19382),
            .I(N__19379));
    InMux I__1846 (
            .O(N__19379),
            .I(N__19376));
    LocalMux I__1845 (
            .O(N__19376),
            .I(N__19373));
    Span12Mux_v I__1844 (
            .O(N__19373),
            .I(N__19370));
    Odrv12 I__1843 (
            .O(N__19370),
            .I(\pwm_generator_inst.un2_threshold_acc_2_6 ));
    InMux I__1842 (
            .O(N__19367),
            .I(N__19364));
    LocalMux I__1841 (
            .O(N__19364),
            .I(N__19361));
    Odrv4 I__1840 (
            .O(N__19361),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ));
    InMux I__1839 (
            .O(N__19358),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ));
    InMux I__1838 (
            .O(N__19355),
            .I(N__19352));
    LocalMux I__1837 (
            .O(N__19352),
            .I(N__19349));
    Span4Mux_v I__1836 (
            .O(N__19349),
            .I(N__19346));
    Span4Mux_v I__1835 (
            .O(N__19346),
            .I(N__19343));
    Odrv4 I__1834 (
            .O(N__19343),
            .I(\pwm_generator_inst.un2_threshold_acc_2_7 ));
    CascadeMux I__1833 (
            .O(N__19340),
            .I(N__19337));
    InMux I__1832 (
            .O(N__19337),
            .I(N__19334));
    LocalMux I__1831 (
            .O(N__19334),
            .I(N__19331));
    Span4Mux_h I__1830 (
            .O(N__19331),
            .I(N__19328));
    Odrv4 I__1829 (
            .O(N__19328),
            .I(\pwm_generator_inst.un2_threshold_acc_1_22 ));
    CascadeMux I__1828 (
            .O(N__19325),
            .I(N__19322));
    InMux I__1827 (
            .O(N__19322),
            .I(N__19319));
    LocalMux I__1826 (
            .O(N__19319),
            .I(N__19316));
    Odrv4 I__1825 (
            .O(N__19316),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ));
    InMux I__1824 (
            .O(N__19313),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ));
    InMux I__1823 (
            .O(N__19310),
            .I(N__19307));
    LocalMux I__1822 (
            .O(N__19307),
            .I(N__19304));
    Span12Mux_h I__1821 (
            .O(N__19304),
            .I(N__19301));
    Odrv12 I__1820 (
            .O(N__19301),
            .I(\pwm_generator_inst.un2_threshold_acc_2_8 ));
    CascadeMux I__1819 (
            .O(N__19298),
            .I(N__19295));
    InMux I__1818 (
            .O(N__19295),
            .I(N__19292));
    LocalMux I__1817 (
            .O(N__19292),
            .I(N__19289));
    Span4Mux_h I__1816 (
            .O(N__19289),
            .I(N__19286));
    Odrv4 I__1815 (
            .O(N__19286),
            .I(\pwm_generator_inst.un2_threshold_acc_1_23 ));
    InMux I__1814 (
            .O(N__19283),
            .I(N__19280));
    LocalMux I__1813 (
            .O(N__19280),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ));
    InMux I__1812 (
            .O(N__19277),
            .I(bfn_2_14_0_));
    InMux I__1811 (
            .O(N__19274),
            .I(N__19271));
    LocalMux I__1810 (
            .O(N__19271),
            .I(N__19268));
    Span4Mux_v I__1809 (
            .O(N__19268),
            .I(N__19265));
    Span4Mux_v I__1808 (
            .O(N__19265),
            .I(N__19262));
    Odrv4 I__1807 (
            .O(N__19262),
            .I(\pwm_generator_inst.un2_threshold_acc_2_9 ));
    CascadeMux I__1806 (
            .O(N__19259),
            .I(N__19256));
    InMux I__1805 (
            .O(N__19256),
            .I(N__19253));
    LocalMux I__1804 (
            .O(N__19253),
            .I(N__19250));
    Span4Mux_h I__1803 (
            .O(N__19250),
            .I(N__19247));
    Odrv4 I__1802 (
            .O(N__19247),
            .I(\pwm_generator_inst.un2_threshold_acc_1_24 ));
    InMux I__1801 (
            .O(N__19244),
            .I(N__19241));
    LocalMux I__1800 (
            .O(N__19241),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ));
    InMux I__1799 (
            .O(N__19238),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ));
    InMux I__1798 (
            .O(N__19235),
            .I(N__19232));
    LocalMux I__1797 (
            .O(N__19232),
            .I(N__19229));
    Span4Mux_v I__1796 (
            .O(N__19229),
            .I(N__19226));
    Span4Mux_v I__1795 (
            .O(N__19226),
            .I(N__19223));
    Odrv4 I__1794 (
            .O(N__19223),
            .I(\pwm_generator_inst.un2_threshold_acc_2_10 ));
    InMux I__1793 (
            .O(N__19220),
            .I(N__19217));
    LocalMux I__1792 (
            .O(N__19217),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ));
    InMux I__1791 (
            .O(N__19214),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ));
    InMux I__1790 (
            .O(N__19211),
            .I(N__19208));
    LocalMux I__1789 (
            .O(N__19208),
            .I(N__19205));
    Span4Mux_v I__1788 (
            .O(N__19205),
            .I(N__19202));
    Span4Mux_v I__1787 (
            .O(N__19202),
            .I(N__19199));
    Odrv4 I__1786 (
            .O(N__19199),
            .I(\pwm_generator_inst.un2_threshold_acc_2_11 ));
    InMux I__1785 (
            .O(N__19196),
            .I(N__19193));
    LocalMux I__1784 (
            .O(N__19193),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ));
    InMux I__1783 (
            .O(N__19190),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ));
    InMux I__1782 (
            .O(N__19187),
            .I(N__19184));
    LocalMux I__1781 (
            .O(N__19184),
            .I(N__19181));
    Span4Mux_v I__1780 (
            .O(N__19181),
            .I(N__19178));
    Span4Mux_v I__1779 (
            .O(N__19178),
            .I(N__19175));
    Odrv4 I__1778 (
            .O(N__19175),
            .I(\pwm_generator_inst.un2_threshold_acc_2_12 ));
    InMux I__1777 (
            .O(N__19172),
            .I(N__19169));
    LocalMux I__1776 (
            .O(N__19169),
            .I(N__19166));
    Odrv4 I__1775 (
            .O(N__19166),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ));
    InMux I__1774 (
            .O(N__19163),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ));
    InMux I__1773 (
            .O(N__19160),
            .I(N__19157));
    LocalMux I__1772 (
            .O(N__19157),
            .I(N__19154));
    Span4Mux_v I__1771 (
            .O(N__19154),
            .I(N__19151));
    Span4Mux_v I__1770 (
            .O(N__19151),
            .I(N__19148));
    Odrv4 I__1769 (
            .O(N__19148),
            .I(\pwm_generator_inst.un2_threshold_acc_2_13 ));
    CascadeMux I__1768 (
            .O(N__19145),
            .I(N__19142));
    InMux I__1767 (
            .O(N__19142),
            .I(N__19139));
    LocalMux I__1766 (
            .O(N__19139),
            .I(N__19136));
    Odrv4 I__1765 (
            .O(N__19136),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ));
    InMux I__1764 (
            .O(N__19133),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ));
    CascadeMux I__1763 (
            .O(N__19130),
            .I(N__19125));
    InMux I__1762 (
            .O(N__19129),
            .I(N__19116));
    InMux I__1761 (
            .O(N__19128),
            .I(N__19116));
    InMux I__1760 (
            .O(N__19125),
            .I(N__19116));
    InMux I__1759 (
            .O(N__19124),
            .I(N__19113));
    InMux I__1758 (
            .O(N__19123),
            .I(N__19110));
    LocalMux I__1757 (
            .O(N__19116),
            .I(N__19105));
    LocalMux I__1756 (
            .O(N__19113),
            .I(N__19105));
    LocalMux I__1755 (
            .O(N__19110),
            .I(\current_shift_inst.PI_CTRL.N_153 ));
    Odrv4 I__1754 (
            .O(N__19105),
            .I(\current_shift_inst.PI_CTRL.N_153 ));
    InMux I__1753 (
            .O(N__19100),
            .I(N__19097));
    LocalMux I__1752 (
            .O(N__19097),
            .I(\current_shift_inst.PI_CTRL.N_155 ));
    InMux I__1751 (
            .O(N__19094),
            .I(N__19091));
    LocalMux I__1750 (
            .O(N__19091),
            .I(N__19088));
    Span12Mux_h I__1749 (
            .O(N__19088),
            .I(N__19085));
    Odrv12 I__1748 (
            .O(N__19085),
            .I(\pwm_generator_inst.un2_threshold_acc_2_0 ));
    CascadeMux I__1747 (
            .O(N__19082),
            .I(N__19079));
    InMux I__1746 (
            .O(N__19079),
            .I(N__19076));
    LocalMux I__1745 (
            .O(N__19076),
            .I(N__19073));
    Span4Mux_h I__1744 (
            .O(N__19073),
            .I(N__19070));
    Odrv4 I__1743 (
            .O(N__19070),
            .I(\pwm_generator_inst.un2_threshold_acc_1_15 ));
    InMux I__1742 (
            .O(N__19067),
            .I(N__19064));
    LocalMux I__1741 (
            .O(N__19064),
            .I(\pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ));
    InMux I__1740 (
            .O(N__19061),
            .I(N__19058));
    LocalMux I__1739 (
            .O(N__19058),
            .I(N__19055));
    Span4Mux_v I__1738 (
            .O(N__19055),
            .I(N__19052));
    Span4Mux_v I__1737 (
            .O(N__19052),
            .I(N__19049));
    Odrv4 I__1736 (
            .O(N__19049),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1 ));
    CascadeMux I__1735 (
            .O(N__19046),
            .I(N__19043));
    InMux I__1734 (
            .O(N__19043),
            .I(N__19040));
    LocalMux I__1733 (
            .O(N__19040),
            .I(N__19037));
    Span4Mux_h I__1732 (
            .O(N__19037),
            .I(N__19034));
    Odrv4 I__1731 (
            .O(N__19034),
            .I(\pwm_generator_inst.un2_threshold_acc_1_16 ));
    CascadeMux I__1730 (
            .O(N__19031),
            .I(N__19028));
    InMux I__1729 (
            .O(N__19028),
            .I(N__19025));
    LocalMux I__1728 (
            .O(N__19025),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ));
    InMux I__1727 (
            .O(N__19022),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ));
    InMux I__1726 (
            .O(N__19019),
            .I(N__19016));
    LocalMux I__1725 (
            .O(N__19016),
            .I(N__19013));
    Span4Mux_v I__1724 (
            .O(N__19013),
            .I(N__19010));
    Span4Mux_v I__1723 (
            .O(N__19010),
            .I(N__19007));
    Odrv4 I__1722 (
            .O(N__19007),
            .I(\pwm_generator_inst.un2_threshold_acc_2_2 ));
    CascadeMux I__1721 (
            .O(N__19004),
            .I(N__19001));
    InMux I__1720 (
            .O(N__19001),
            .I(N__18998));
    LocalMux I__1719 (
            .O(N__18998),
            .I(N__18995));
    Span4Mux_v I__1718 (
            .O(N__18995),
            .I(N__18992));
    Odrv4 I__1717 (
            .O(N__18992),
            .I(\pwm_generator_inst.un2_threshold_acc_1_17 ));
    InMux I__1716 (
            .O(N__18989),
            .I(N__18986));
    LocalMux I__1715 (
            .O(N__18986),
            .I(N__18983));
    Odrv4 I__1714 (
            .O(N__18983),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ));
    InMux I__1713 (
            .O(N__18980),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ));
    InMux I__1712 (
            .O(N__18977),
            .I(N__18974));
    LocalMux I__1711 (
            .O(N__18974),
            .I(N__18971));
    Span4Mux_v I__1710 (
            .O(N__18971),
            .I(N__18968));
    Span4Mux_v I__1709 (
            .O(N__18968),
            .I(N__18965));
    Odrv4 I__1708 (
            .O(N__18965),
            .I(\pwm_generator_inst.un2_threshold_acc_2_3 ));
    CascadeMux I__1707 (
            .O(N__18962),
            .I(N__18959));
    InMux I__1706 (
            .O(N__18959),
            .I(N__18956));
    LocalMux I__1705 (
            .O(N__18956),
            .I(N__18953));
    Span4Mux_h I__1704 (
            .O(N__18953),
            .I(N__18950));
    Odrv4 I__1703 (
            .O(N__18950),
            .I(\pwm_generator_inst.un2_threshold_acc_1_18 ));
    CascadeMux I__1702 (
            .O(N__18947),
            .I(N__18944));
    InMux I__1701 (
            .O(N__18944),
            .I(N__18941));
    LocalMux I__1700 (
            .O(N__18941),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ));
    InMux I__1699 (
            .O(N__18938),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ));
    InMux I__1698 (
            .O(N__18935),
            .I(N__18932));
    LocalMux I__1697 (
            .O(N__18932),
            .I(N__18929));
    Span4Mux_v I__1696 (
            .O(N__18929),
            .I(N__18926));
    Span4Mux_v I__1695 (
            .O(N__18926),
            .I(N__18923));
    Odrv4 I__1694 (
            .O(N__18923),
            .I(\pwm_generator_inst.un2_threshold_acc_2_4 ));
    CascadeMux I__1693 (
            .O(N__18920),
            .I(N__18917));
    InMux I__1692 (
            .O(N__18917),
            .I(N__18914));
    LocalMux I__1691 (
            .O(N__18914),
            .I(N__18911));
    Span4Mux_h I__1690 (
            .O(N__18911),
            .I(N__18908));
    Odrv4 I__1689 (
            .O(N__18908),
            .I(\pwm_generator_inst.un2_threshold_acc_1_19 ));
    InMux I__1688 (
            .O(N__18905),
            .I(N__18902));
    LocalMux I__1687 (
            .O(N__18902),
            .I(N__18899));
    Odrv4 I__1686 (
            .O(N__18899),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ));
    InMux I__1685 (
            .O(N__18896),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ));
    InMux I__1684 (
            .O(N__18893),
            .I(N__18890));
    LocalMux I__1683 (
            .O(N__18890),
            .I(N__18887));
    Span4Mux_v I__1682 (
            .O(N__18887),
            .I(N__18884));
    Span4Mux_v I__1681 (
            .O(N__18884),
            .I(N__18881));
    Odrv4 I__1680 (
            .O(N__18881),
            .I(\pwm_generator_inst.un2_threshold_acc_2_5 ));
    CascadeMux I__1679 (
            .O(N__18878),
            .I(N__18875));
    InMux I__1678 (
            .O(N__18875),
            .I(N__18872));
    LocalMux I__1677 (
            .O(N__18872),
            .I(N__18869));
    Span4Mux_v I__1676 (
            .O(N__18869),
            .I(N__18866));
    Span4Mux_h I__1675 (
            .O(N__18866),
            .I(N__18863));
    Odrv4 I__1674 (
            .O(N__18863),
            .I(\pwm_generator_inst.un2_threshold_acc_1_20 ));
    CascadeMux I__1673 (
            .O(N__18860),
            .I(N__18857));
    InMux I__1672 (
            .O(N__18857),
            .I(N__18854));
    LocalMux I__1671 (
            .O(N__18854),
            .I(N__18851));
    Odrv4 I__1670 (
            .O(N__18851),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ));
    InMux I__1669 (
            .O(N__18848),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ));
    InMux I__1668 (
            .O(N__18845),
            .I(N__18840));
    InMux I__1667 (
            .O(N__18844),
            .I(N__18835));
    InMux I__1666 (
            .O(N__18843),
            .I(N__18835));
    LocalMux I__1665 (
            .O(N__18840),
            .I(N__18832));
    LocalMux I__1664 (
            .O(N__18835),
            .I(pwm_duty_input_4));
    Odrv4 I__1663 (
            .O(N__18832),
            .I(pwm_duty_input_4));
    CascadeMux I__1662 (
            .O(N__18827),
            .I(N__18822));
    CascadeMux I__1661 (
            .O(N__18826),
            .I(N__18819));
    InMux I__1660 (
            .O(N__18825),
            .I(N__18816));
    InMux I__1659 (
            .O(N__18822),
            .I(N__18811));
    InMux I__1658 (
            .O(N__18819),
            .I(N__18811));
    LocalMux I__1657 (
            .O(N__18816),
            .I(N__18808));
    LocalMux I__1656 (
            .O(N__18811),
            .I(N__18805));
    Span4Mux_s1_h I__1655 (
            .O(N__18808),
            .I(N__18802));
    Odrv4 I__1654 (
            .O(N__18805),
            .I(pwm_duty_input_3));
    Odrv4 I__1653 (
            .O(N__18802),
            .I(pwm_duty_input_3));
    InMux I__1652 (
            .O(N__18797),
            .I(N__18793));
    InMux I__1651 (
            .O(N__18796),
            .I(N__18790));
    LocalMux I__1650 (
            .O(N__18793),
            .I(N__18787));
    LocalMux I__1649 (
            .O(N__18790),
            .I(pwm_duty_input_0));
    Odrv4 I__1648 (
            .O(N__18787),
            .I(pwm_duty_input_0));
    InMux I__1647 (
            .O(N__18782),
            .I(N__18779));
    LocalMux I__1646 (
            .O(N__18779),
            .I(N__18775));
    InMux I__1645 (
            .O(N__18778),
            .I(N__18772));
    Span4Mux_v I__1644 (
            .O(N__18775),
            .I(N__18769));
    LocalMux I__1643 (
            .O(N__18772),
            .I(pwm_duty_input_1));
    Odrv4 I__1642 (
            .O(N__18769),
            .I(pwm_duty_input_1));
    InMux I__1641 (
            .O(N__18764),
            .I(N__18761));
    LocalMux I__1640 (
            .O(N__18761),
            .I(N__18757));
    InMux I__1639 (
            .O(N__18760),
            .I(N__18754));
    Span4Mux_s1_h I__1638 (
            .O(N__18757),
            .I(N__18751));
    LocalMux I__1637 (
            .O(N__18754),
            .I(pwm_duty_input_2));
    Odrv4 I__1636 (
            .O(N__18751),
            .I(pwm_duty_input_2));
    InMux I__1635 (
            .O(N__18746),
            .I(N__18743));
    LocalMux I__1634 (
            .O(N__18743),
            .I(\pwm_generator_inst.un1_duty_inputlt3 ));
    CascadeMux I__1633 (
            .O(N__18740),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ));
    CascadeMux I__1632 (
            .O(N__18737),
            .I(N__18734));
    InMux I__1631 (
            .O(N__18734),
            .I(N__18728));
    InMux I__1630 (
            .O(N__18733),
            .I(N__18728));
    LocalMux I__1629 (
            .O(N__18728),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    CascadeMux I__1628 (
            .O(N__18725),
            .I(\current_shift_inst.PI_CTRL.N_31_cascade_ ));
    InMux I__1627 (
            .O(N__18722),
            .I(N__18719));
    LocalMux I__1626 (
            .O(N__18719),
            .I(N__18716));
    Odrv4 I__1625 (
            .O(N__18716),
            .I(\current_shift_inst.PI_CTRL.N_149 ));
    CascadeMux I__1624 (
            .O(N__18713),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ));
    InMux I__1623 (
            .O(N__18710),
            .I(N__18707));
    LocalMux I__1622 (
            .O(N__18707),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    CascadeMux I__1621 (
            .O(N__18704),
            .I(\current_shift_inst.PI_CTRL.N_27_cascade_ ));
    InMux I__1620 (
            .O(N__18701),
            .I(N__18695));
    InMux I__1619 (
            .O(N__18700),
            .I(N__18695));
    LocalMux I__1618 (
            .O(N__18695),
            .I(N__18692));
    Odrv4 I__1617 (
            .O(N__18692),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ));
    CascadeMux I__1616 (
            .O(N__18689),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_ ));
    InMux I__1615 (
            .O(N__18686),
            .I(N__18683));
    LocalMux I__1614 (
            .O(N__18683),
            .I(N_38_i_i));
    InMux I__1613 (
            .O(N__18680),
            .I(N__18677));
    LocalMux I__1612 (
            .O(N__18677),
            .I(rgb_drv_RNOZ0));
    InMux I__1611 (
            .O(N__18674),
            .I(N__18671));
    LocalMux I__1610 (
            .O(N__18671),
            .I(N__18668));
    Span4Mux_h I__1609 (
            .O(N__18668),
            .I(N__18664));
    InMux I__1608 (
            .O(N__18667),
            .I(N__18661));
    Odrv4 I__1607 (
            .O(N__18664),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_15 ));
    LocalMux I__1606 (
            .O(N__18661),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_15 ));
    InMux I__1605 (
            .O(N__18656),
            .I(N__18653));
    LocalMux I__1604 (
            .O(N__18653),
            .I(N__18650));
    Odrv4 I__1603 (
            .O(N__18650),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_16 ));
    InMux I__1602 (
            .O(N__18647),
            .I(N__18638));
    InMux I__1601 (
            .O(N__18646),
            .I(N__18638));
    InMux I__1600 (
            .O(N__18645),
            .I(N__18638));
    LocalMux I__1599 (
            .O(N__18638),
            .I(\current_shift_inst.PI_CTRL.N_154 ));
    InMux I__1598 (
            .O(N__18635),
            .I(N__18632));
    LocalMux I__1597 (
            .O(N__18632),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ));
    CascadeMux I__1596 (
            .O(N__18629),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3_cascade_ ));
    CascadeMux I__1595 (
            .O(N__18626),
            .I(N__18622));
    CascadeMux I__1594 (
            .O(N__18625),
            .I(N__18619));
    InMux I__1593 (
            .O(N__18622),
            .I(N__18613));
    InMux I__1592 (
            .O(N__18619),
            .I(N__18613));
    InMux I__1591 (
            .O(N__18618),
            .I(N__18610));
    LocalMux I__1590 (
            .O(N__18613),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_3 ));
    LocalMux I__1589 (
            .O(N__18610),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_3 ));
    InMux I__1588 (
            .O(N__18605),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_19 ));
    InMux I__1587 (
            .O(N__18602),
            .I(N__18596));
    InMux I__1586 (
            .O(N__18601),
            .I(N__18596));
    LocalMux I__1585 (
            .O(N__18596),
            .I(N__18593));
    Odrv4 I__1584 (
            .O(N__18593),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ));
    CascadeMux I__1583 (
            .O(N__18590),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_ ));
    InMux I__1582 (
            .O(N__18587),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4 ));
    InMux I__1581 (
            .O(N__18584),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5 ));
    InMux I__1580 (
            .O(N__18581),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6 ));
    InMux I__1579 (
            .O(N__18578),
            .I(bfn_1_15_0_));
    IoInMux I__1578 (
            .O(N__18575),
            .I(N__18572));
    LocalMux I__1577 (
            .O(N__18572),
            .I(N__18569));
    IoSpan4Mux I__1576 (
            .O(N__18569),
            .I(N__18566));
    Sp12to4 I__1575 (
            .O(N__18566),
            .I(N__18563));
    Span12Mux_s6_v I__1574 (
            .O(N__18563),
            .I(N__18560));
    Span12Mux_h I__1573 (
            .O(N__18560),
            .I(N__18557));
    Odrv12 I__1572 (
            .O(N__18557),
            .I(\pll_inst.red_c_i ));
    InMux I__1571 (
            .O(N__18554),
            .I(N__18551));
    LocalMux I__1570 (
            .O(N__18551),
            .I(N__18548));
    Odrv4 I__1569 (
            .O(N__18548),
            .I(\pwm_generator_inst.O_12 ));
    InMux I__1568 (
            .O(N__18545),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0 ));
    InMux I__1567 (
            .O(N__18542),
            .I(N__18539));
    LocalMux I__1566 (
            .O(N__18539),
            .I(N__18536));
    Odrv4 I__1565 (
            .O(N__18536),
            .I(\pwm_generator_inst.O_13 ));
    InMux I__1564 (
            .O(N__18533),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1 ));
    InMux I__1563 (
            .O(N__18530),
            .I(N__18527));
    LocalMux I__1562 (
            .O(N__18527),
            .I(N__18524));
    Span4Mux_h I__1561 (
            .O(N__18524),
            .I(N__18521));
    Odrv4 I__1560 (
            .O(N__18521),
            .I(\pwm_generator_inst.O_14 ));
    InMux I__1559 (
            .O(N__18518),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2 ));
    InMux I__1558 (
            .O(N__18515),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3 ));
    IoInMux I__1557 (
            .O(N__18512),
            .I(N__18509));
    LocalMux I__1556 (
            .O(N__18509),
            .I(N__18506));
    Span4Mux_s3_v I__1555 (
            .O(N__18506),
            .I(N__18503));
    Span4Mux_h I__1554 (
            .O(N__18503),
            .I(N__18500));
    Sp12to4 I__1553 (
            .O(N__18500),
            .I(N__18497));
    Span12Mux_v I__1552 (
            .O(N__18497),
            .I(N__18494));
    Span12Mux_v I__1551 (
            .O(N__18494),
            .I(N__18491));
    Odrv12 I__1550 (
            .O(N__18491),
            .I(delay_tr_input_ibuf_gb_io_gb_input));
    IoInMux I__1549 (
            .O(N__18488),
            .I(N__18485));
    LocalMux I__1548 (
            .O(N__18485),
            .I(N__18482));
    IoSpan4Mux I__1547 (
            .O(N__18482),
            .I(N__18479));
    IoSpan4Mux I__1546 (
            .O(N__18479),
            .I(N__18476));
    Odrv4 I__1545 (
            .O(N__18476),
            .I(delay_hc_input_ibuf_gb_io_gb_input));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_6 ),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_14 ),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_22 ),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_9_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_30 ),
            .carryinitout(bfn_9_12_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_acc_cry_7 ),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_1_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_16_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_acc_cry_15 ),
            .carryinitout(bfn_1_16_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_15_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_14_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_15_14_0_));
    defparam IN_MUX_bfv_15_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_15_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_15_15_0_));
    defparam IN_MUX_bfv_8_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_19_0_));
    defparam IN_MUX_bfv_8_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_20_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_8_20_0_));
    defparam IN_MUX_bfv_8_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_21_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_8_21_0_));
    defparam IN_MUX_bfv_18_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_11_0_));
    defparam IN_MUX_bfv_18_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_12_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_18_12_0_));
    defparam IN_MUX_bfv_18_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_13_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_18_13_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_8_15_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_14_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_19_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .carryinitout(bfn_14_19_0_));
    defparam IN_MUX_bfv_14_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_20_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .carryinitout(bfn_14_20_0_));
    defparam IN_MUX_bfv_14_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_21_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .carryinitout(bfn_14_21_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_16_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_16_0_));
    defparam IN_MUX_bfv_16_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_17_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_7 ),
            .carryinitout(bfn_16_17_0_));
    defparam IN_MUX_bfv_16_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_18_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_15 ),
            .carryinitout(bfn_16_18_0_));
    defparam IN_MUX_bfv_16_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_19_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_23 ),
            .carryinitout(bfn_16_19_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_13_0_));
    defparam IN_MUX_bfv_2_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_14_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ),
            .carryinitout(bfn_2_14_0_));
    defparam IN_MUX_bfv_2_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_15_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ),
            .carryinitout(bfn_2_15_0_));
    defparam IN_MUX_bfv_2_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_16_0_));
    defparam IN_MUX_bfv_2_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_17_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_acc_1_cry_7 ),
            .carryinitout(bfn_2_17_0_));
    defparam IN_MUX_bfv_2_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_18_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_acc_1_cry_15 ),
            .carryinitout(bfn_2_18_0_));
    defparam IN_MUX_bfv_3_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_12_0_));
    defparam IN_MUX_bfv_3_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_13_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_3_13_0_));
    defparam IN_MUX_bfv_3_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_17_0_));
    defparam IN_MUX_bfv_3_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_18_0_ (
            .carryinitin(\pwm_generator_inst.un19_threshold_acc_cry_7 ),
            .carryinitout(bfn_3_18_0_));
    defparam IN_MUX_bfv_4_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_13_0_));
    defparam IN_MUX_bfv_4_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_14_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_4_14_0_));
    defparam IN_MUX_bfv_15_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_10_0_));
    defparam IN_MUX_bfv_15_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_11_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un6_running_cry_8 ),
            .carryinitout(bfn_15_11_0_));
    defparam IN_MUX_bfv_15_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_12_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un6_running_cry_16 ),
            .carryinitout(bfn_15_12_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_9_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_20_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un6_running_cry_8 ),
            .carryinitout(bfn_9_20_0_));
    defparam IN_MUX_bfv_9_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_21_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un6_running_cry_16 ),
            .carryinitout(bfn_9_21_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un6_running_cry_8 ),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_17_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_12_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un6_running_cry_16 ),
            .carryinitout(bfn_17_12_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un6_running_cry_8 ),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un6_running_cry_16 ),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_13_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_9_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_13_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_11_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_13_11_0_));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_13_12_0_));
    defparam IN_MUX_bfv_13_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_5_0_));
    defparam IN_MUX_bfv_13_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_6_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_13_6_0_));
    defparam IN_MUX_bfv_13_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_7_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_13_7_0_));
    defparam IN_MUX_bfv_13_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_13_8_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_11_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_16_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_11_16_0_));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_11_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_19_0_));
    defparam IN_MUX_bfv_11_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_20_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_11_20_0_));
    defparam IN_MUX_bfv_11_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_21_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_11_21_0_));
    defparam IN_MUX_bfv_11_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_22_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_11_22_0_));
    defparam IN_MUX_bfv_18_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_19_0_));
    defparam IN_MUX_bfv_18_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_20_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_18_20_0_));
    defparam IN_MUX_bfv_18_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_21_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_18_21_0_));
    defparam IN_MUX_bfv_18_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_22_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_18_22_0_));
    defparam IN_MUX_bfv_17_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_15_0_));
    defparam IN_MUX_bfv_17_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_16_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_8 ),
            .carryinitout(bfn_17_16_0_));
    defparam IN_MUX_bfv_17_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_17_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_16 ),
            .carryinitout(bfn_17_17_0_));
    defparam IN_MUX_bfv_17_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_18_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_24 ),
            .carryinitout(bfn_17_18_0_));
    defparam IN_MUX_bfv_16_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_21_0_));
    defparam IN_MUX_bfv_16_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_22_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_16_22_0_));
    defparam IN_MUX_bfv_16_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_23_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_16_23_0_));
    defparam IN_MUX_bfv_16_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_24_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_16_24_0_));
    defparam IN_MUX_bfv_15_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_16_0_));
    defparam IN_MUX_bfv_15_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_17_0_ (
            .carryinitin(\current_shift_inst.control_input_1_cry_7 ),
            .carryinitout(bfn_15_17_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_11_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ),
            .carryinitout(bfn_11_12_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_5_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_9_0_));
    defparam IN_MUX_bfv_5_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_10_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryinitout(bfn_5_10_0_));
    defparam IN_MUX_bfv_5_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_11_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryinitout(bfn_5_11_0_));
    defparam IN_MUX_bfv_5_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryinitout(bfn_5_12_0_));
    defparam IN_MUX_bfv_12_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_11_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .carryinitout(bfn_12_12_0_));
    ICE_GB delay_tr_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__18512),
            .GLOBALBUFFEROUTPUT(delay_tr_input_c_g));
    ICE_GB delay_hc_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__18488),
            .GLOBALBUFFEROUTPUT(delay_hc_input_c_g));
    ICE_GB \current_shift_inst.timer_s1.running_RNII51H_0  (
            .USERSIGNALTOGLOBALBUFFER(N__37628),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_166_i_g ));
    ICE_GB \delay_measurement_inst.delay_tr_timer.running_RNICNBI_0  (
            .USERSIGNALTOGLOBALBUFFER(N__23594),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_tr_timer.N_434_i_g ));
    ICE_GB \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0  (
            .USERSIGNALTOGLOBALBUFFER(N__30617),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_hc_timer.N_432_i_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__39048),
            .CLKHFEN(N__39068),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__39067),
            .RGB2PWM(N__18686),
            .RGB1(rgb_g),
            .CURREN(N__38975),
            .RGB2(rgb_b),
            .RGB1PWM(N__18680),
            .RGB0PWM(N__47483),
            .RGB0(rgb_r));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_5_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_5_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_5_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_5_0  (
            .in0(N__19541),
            .in1(N__18667),
            .in2(_gnd_net_),
            .in3(N__21358),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22253),
            .lcout(N_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47876),
            .ce(),
            .sr(N__47362));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_9_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_9_1 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_1_9_1  (
            .in0(N__18618),
            .in1(N__21857),
            .in2(N__19130),
            .in3(N__18646),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47874),
            .ce(),
            .sr(N__47386));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_9_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_9_4 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_1_9_4  (
            .in0(N__18647),
            .in1(N__21845),
            .in2(N__18626),
            .in3(N__19129),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47874),
            .ce(),
            .sr(N__47386));
    defparam \pwm_generator_inst.threshold_5_LC_1_9_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_5_LC_1_9_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_5_LC_1_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_5_LC_1_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20039),
            .lcout(\pwm_generator_inst.thresholdZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47874),
            .ce(),
            .sr(N__47386));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_9_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_9_6 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_1_9_6  (
            .in0(N__18645),
            .in1(N__21866),
            .in2(N__18625),
            .in3(N__19128),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47874),
            .ce(),
            .sr(N__47386));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_10_1 .LUT_INIT=16'b1010000011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_1_10_1  (
            .in0(N__21731),
            .in1(N__20257),
            .in2(N__20205),
            .in3(N__22243),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47873),
            .ce(),
            .sr(N__47389));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_10_3 .LUT_INIT=16'b1010000011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_1_10_3  (
            .in0(N__21697),
            .in1(N__20258),
            .in2(N__20206),
            .in3(N__22244),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47873),
            .ce(),
            .sr(N__47389));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_10_4 .LUT_INIT=16'b1100111100001010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_1_10_4  (
            .in0(N__20253),
            .in1(N__20191),
            .in2(N__22252),
            .in3(N__22030),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47873),
            .ce(),
            .sr(N__47389));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_10_5 .LUT_INIT=16'b0000000011011111;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_1_10_5  (
            .in0(N__18710),
            .in1(N__21806),
            .in2(N__20204),
            .in3(N__18722),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47873),
            .ce(),
            .sr(N__47389));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_10_6 .LUT_INIT=16'b1010101011111011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_1_10_6  (
            .in0(N__21833),
            .in1(N__18635),
            .in2(N__20261),
            .in3(N__19123),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47873),
            .ce(),
            .sr(N__47389));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_10_7 .LUT_INIT=16'b1010000011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_1_10_7  (
            .in0(N__21997),
            .in1(N__20259),
            .in2(N__20207),
            .in3(N__22248),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47873),
            .ce(),
            .sr(N__47389));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_11_7 .LUT_INIT=16'b1111010001010100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_1_11_7  (
            .in0(N__22242),
            .in1(N__20260),
            .in2(N__21761),
            .in3(N__20190),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47871),
            .ce(),
            .sr(N__47395));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_1_13_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_1_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_1_13_1  (
            .in0(N__21246),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21220),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_1_13_3 .C_ON=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_1_13_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_1_13_3  (
            .in0(N__47480),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pll_inst.red_c_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_14_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(N__19822),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_14_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_14_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_14_1  (
            .in0(_gnd_net_),
            .in1(N__18554),
            .in2(_gnd_net_),
            .in3(N__18545),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_14_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(N__18542),
            .in2(_gnd_net_),
            .in3(N__18533),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_14_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_14_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_14_3  (
            .in0(_gnd_net_),
            .in1(N__18530),
            .in2(_gnd_net_),
            .in3(N__18518),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_14_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(N__19067),
            .in2(_gnd_net_),
            .in3(N__18515),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_14_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_14_5  (
            .in0(_gnd_net_),
            .in1(N__38985),
            .in2(N__19031),
            .in3(N__18587),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_14_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_14_6  (
            .in0(_gnd_net_),
            .in1(N__18989),
            .in2(N__39055),
            .in3(N__18584),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_14_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(N__38989),
            .in2(N__18947),
            .in3(N__18581),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_15_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(N__18905),
            .in2(_gnd_net_),
            .in3(N__18578),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ),
            .ltout(),
            .carryin(bfn_1_15_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_15_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18860),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_15_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_15_2  (
            .in0(_gnd_net_),
            .in1(N__19367),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_15_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19325),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_15_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_15_4  (
            .in0(_gnd_net_),
            .in1(N__19283),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_15_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_15_5  (
            .in0(_gnd_net_),
            .in1(N__19244),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_15_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_15_6  (
            .in0(_gnd_net_),
            .in1(N__19220),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_15_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_15_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_15_7  (
            .in0(_gnd_net_),
            .in1(N__19196),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_16_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_16_0  (
            .in0(_gnd_net_),
            .in1(N__19172),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_16_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_16_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_16_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19145),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_16_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_16_2  (
            .in0(_gnd_net_),
            .in1(N__19568),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_16_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19466),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_16_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_16_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18605),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_1_16_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_1_16_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_1_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_1_16_6  (
            .in0(N__19802),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19424),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_1_17_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_1_17_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_1_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_1_17_3  (
            .in0(_gnd_net_),
            .in1(N__20093),
            .in2(_gnd_net_),
            .in3(N__18601),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_1_17_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_1_17_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_1_17_4 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_1_17_4  (
            .in0(N__18602),
            .in1(N__21202),
            .in2(N__18590),
            .in3(N__20081),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_1_17_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_1_17_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_1_17_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_1_17_5  (
            .in0(_gnd_net_),
            .in1(N__18700),
            .in2(_gnd_net_),
            .in3(N__20072),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_1_17_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_1_17_6 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_1_17_6  (
            .in0(N__18701),
            .in1(N__21203),
            .in2(N__18689),
            .in3(N__20060),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_17_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_17_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_17_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_17_7  (
            .in0(_gnd_net_),
            .in1(N__20476),
            .in2(_gnd_net_),
            .in3(N__20449),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_drv_RNO_0_LC_1_29_2.C_ON=1'b0;
    defparam rgb_drv_RNO_0_LC_1_29_2.SEQ_MODE=4'b0000;
    defparam rgb_drv_RNO_0_LC_1_29_2.LUT_INIT=16'b1010101001010101;
    LogicCell40 rgb_drv_RNO_0_LC_1_29_2 (
            .in0(N__47481),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34159),
            .lcout(N_38_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_drv_RNO_LC_1_30_2.C_ON=1'b0;
    defparam rgb_drv_RNO_LC_1_30_2.SEQ_MODE=4'b0000;
    defparam rgb_drv_RNO_LC_1_30_2.LUT_INIT=16'b0101010100000000;
    LogicCell40 rgb_drv_RNO_LC_1_30_2 (
            .in0(N__47482),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34163),
            .lcout(rgb_drv_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_2_7_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_2_7_6 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_2_7_6  (
            .in0(N__18674),
            .in1(N__19540),
            .in2(N__21379),
            .in3(N__18656),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_9_0 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_9_0  (
            .in0(N__22240),
            .in1(_gnd_net_),
            .in2(N__18737),
            .in3(N__20233),
            .lcout(\current_shift_inst.PI_CTRL.N_154 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_9_5 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_9_5  (
            .in0(N__21797),
            .in1(N__22239),
            .in2(_gnd_net_),
            .in3(N__18733),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_9_6 .LUT_INIT=16'b0101010100010000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_9_6  (
            .in0(N__21831),
            .in1(N__20234),
            .in2(N__18629),
            .in3(N__19124),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_10_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_10_0 .LUT_INIT=16'b1011101110101011;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_LC_2_10_0  (
            .in0(N__19928),
            .in1(N__18844),
            .in2(N__18826),
            .in3(N__18746),
            .lcout(\pwm_generator_inst.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_10_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_10_2 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_10_2  (
            .in0(N__20045),
            .in1(N__18843),
            .in2(N__18827),
            .in3(N__20290),
            .lcout(\pwm_generator_inst.N_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_10_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_10_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pwm_generator_inst.un1_duty_inputlto2_LC_2_10_3  (
            .in0(N__18796),
            .in1(N__18778),
            .in2(_gnd_net_),
            .in3(N__18760),
            .lcout(\pwm_generator_inst.un1_duty_inputlt3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_10_4 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_10_4  (
            .in0(N__21996),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21756),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_10_5 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_10_5  (
            .in0(N__22029),
            .in1(N__21696),
            .in2(N__18740),
            .in3(N__21730),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(\current_shift_inst.PI_CTRL.N_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_10_6 .LUT_INIT=16'b0011001100010011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_10_6  (
            .in0(N__21805),
            .in1(N__22241),
            .in2(N__18725),
            .in3(N__20235),
            .lcout(\current_shift_inst.PI_CTRL.N_149 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_2_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_2_11_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(N__22001),
            .in2(_gnd_net_),
            .in3(N__21729),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_2_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_2_11_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_2_11_3  (
            .in0(N__22031),
            .in1(N__21698),
            .in2(N__18713),
            .in3(N__21757),
            .lcout(\current_shift_inst.PI_CTRL.N_27 ),
            .ltout(\current_shift_inst.PI_CTRL.N_27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_11_4 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_11_4  (
            .in0(N__22215),
            .in1(N__19100),
            .in2(N__18704),
            .in3(N__20172),
            .lcout(\current_shift_inst.PI_CTRL.N_153 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_11_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(N__21801),
            .in2(_gnd_net_),
            .in3(N__21832),
            .lcout(\current_shift_inst.PI_CTRL.N_155 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_13_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_13_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(N__19094),
            .in2(N__19082),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ),
            .ltout(),
            .carryin(bfn_2_13_0_),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_13_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(N__19061),
            .in2(N__19046),
            .in3(N__19022),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_13_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_13_2  (
            .in0(_gnd_net_),
            .in1(N__19019),
            .in2(N__19004),
            .in3(N__18980),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_13_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__18977),
            .in2(N__18962),
            .in3(N__18938),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_13_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_13_4  (
            .in0(_gnd_net_),
            .in1(N__18935),
            .in2(N__18920),
            .in3(N__18896),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_13_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_13_5  (
            .in0(_gnd_net_),
            .in1(N__18893),
            .in2(N__18878),
            .in3(N__18848),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_13_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_13_6  (
            .in0(_gnd_net_),
            .in1(N__19394),
            .in2(N__19382),
            .in3(N__19358),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_13_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_13_7  (
            .in0(_gnd_net_),
            .in1(N__19355),
            .in2(N__19340),
            .in3(N__19313),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_14_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(N__19310),
            .in2(N__19298),
            .in3(N__19277),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ),
            .ltout(),
            .carryin(bfn_2_14_0_),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_14_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(N__19274),
            .in2(N__19259),
            .in3(N__19238),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_14_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(N__19235),
            .in2(N__19535),
            .in3(N__19214),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_14_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_14_3  (
            .in0(_gnd_net_),
            .in1(N__19211),
            .in2(N__19537),
            .in3(N__19190),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_14_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_14_4  (
            .in0(_gnd_net_),
            .in1(N__19187),
            .in2(N__19536),
            .in3(N__19163),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_14_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_14_5  (
            .in0(_gnd_net_),
            .in1(N__19160),
            .in2(N__19538),
            .in3(N__19133),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_14_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_14_6  (
            .in0(_gnd_net_),
            .in1(N__19525),
            .in2(N__19583),
            .in3(N__19559),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_14_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_14_7  (
            .in0(_gnd_net_),
            .in1(N__19556),
            .in2(N__19539),
            .in3(N__19454),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_15_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_15_0  (
            .in0(N__19451),
            .in1(N__19439),
            .in2(_gnd_net_),
            .in3(N__19427),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ),
            .ltout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_15_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_15_1 .LUT_INIT=16'b1010110001011100;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_15_1  (
            .in0(N__19784),
            .in1(N__19423),
            .in2(N__19409),
            .in3(N__19801),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_15_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_15_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_15_2  (
            .in0(N__20674),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20658),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_15_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_15_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(N__19405),
            .in2(_gnd_net_),
            .in3(N__20119),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_15_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_15_4 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_15_4  (
            .in0(N__19406),
            .in1(N__21169),
            .in2(N__19397),
            .in3(N__20105),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_2_15_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_2_15_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_2_15_6  (
            .in0(_gnd_net_),
            .in1(N__19738),
            .in2(_gnd_net_),
            .in3(N__19768),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_15_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_15_7 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_15_7  (
            .in0(N__19739),
            .in1(N__19754),
            .in2(N__19730),
            .in3(N__21168),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_2_16_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_2_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_2_16_0  (
            .in0(_gnd_net_),
            .in1(N__19712),
            .in2(_gnd_net_),
            .in3(N__19727),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_0 ),
            .ltout(),
            .carryin(bfn_2_16_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_2_16_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_2_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_2_16_1  (
            .in0(_gnd_net_),
            .in1(N__19691),
            .in2(_gnd_net_),
            .in3(N__19706),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_0 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_2_16_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_2_16_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_2_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_2_16_2  (
            .in0(_gnd_net_),
            .in1(N__19670),
            .in2(_gnd_net_),
            .in3(N__19685),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_1 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_2_16_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_2_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_2_16_3  (
            .in0(_gnd_net_),
            .in1(N__19649),
            .in2(_gnd_net_),
            .in3(N__19664),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_2 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_2_16_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_2_16_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_2_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_2_16_4  (
            .in0(_gnd_net_),
            .in1(N__19628),
            .in2(_gnd_net_),
            .in3(N__19643),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_3 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_2_16_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_2_16_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_2_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_2_16_5  (
            .in0(_gnd_net_),
            .in1(N__19607),
            .in2(_gnd_net_),
            .in3(N__19622),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_4 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_2_16_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_2_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_2_16_6  (
            .in0(_gnd_net_),
            .in1(N__19589),
            .in2(_gnd_net_),
            .in3(N__19601),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_5 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_2_16_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_2_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_2_16_7  (
            .in0(_gnd_net_),
            .in1(N__19880),
            .in2(_gnd_net_),
            .in3(N__19895),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_6 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_2_17_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_2_17_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_2_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_2_17_0  (
            .in0(_gnd_net_),
            .in1(N__19859),
            .in2(_gnd_net_),
            .in3(N__19874),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_8 ),
            .ltout(),
            .carryin(bfn_2_17_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_2_17_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_2_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_2_17_1  (
            .in0(_gnd_net_),
            .in1(N__19838),
            .in2(_gnd_net_),
            .in3(N__19853),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_8 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_2_17_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_2_17_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_2_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_2_17_2  (
            .in0(_gnd_net_),
            .in1(N__20445),
            .in2(_gnd_net_),
            .in3(N__19832),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_2_17_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_2_17_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_2_17_3  (
            .in0(N__21176),
            .in1(N__19829),
            .in2(_gnd_net_),
            .in3(N__19805),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_2_17_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_2_17_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_2_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_2_17_4  (
            .in0(_gnd_net_),
            .in1(N__19800),
            .in2(_gnd_net_),
            .in3(N__19775),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_2_17_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_2_17_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_2_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_2_17_5  (
            .in0(_gnd_net_),
            .in1(N__21253),
            .in2(_gnd_net_),
            .in3(N__19772),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_2_17_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_2_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_2_17_6  (
            .in0(_gnd_net_),
            .in1(N__19769),
            .in2(_gnd_net_),
            .in3(N__19742),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_2_17_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_2_17_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_2_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_2_17_7  (
            .in0(_gnd_net_),
            .in1(N__20120),
            .in2(_gnd_net_),
            .in3(N__20096),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_2_18_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_2_18_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_2_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_2_18_0  (
            .in0(_gnd_net_),
            .in1(N__20092),
            .in2(_gnd_net_),
            .in3(N__20075),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_2_18_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_2_18_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_2_18_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_2_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_2_18_1  (
            .in0(_gnd_net_),
            .in1(N__20071),
            .in2(_gnd_net_),
            .in3(N__20054),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_2_18_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_2_18_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_2_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_2_18_2  (
            .in0(_gnd_net_),
            .in1(N__20662),
            .in2(_gnd_net_),
            .in3(N__20051),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_2_18_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_2_18_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_2_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_2_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20048),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_3_9_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_3_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_3_9_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_3_9_1  (
            .in0(N__19922),
            .in1(N__19999),
            .in2(N__19963),
            .in3(N__20030),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_5_LC_3_9_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_5_LC_3_9_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_5_LC_3_9_7 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_5_LC_3_9_7  (
            .in0(N__21486),
            .in1(N__20756),
            .in2(N__21439),
            .in3(N__21554),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47872),
            .ce(),
            .sr(N__47371));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_10_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_10_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_10_0 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_10_0  (
            .in0(N__20026),
            .in1(N__20000),
            .in2(N__19964),
            .in3(N__20270),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_3_10_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_3_10_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_3_10_3 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_3_10_3  (
            .in0(N__19921),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20294),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_3_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_3_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_3_10_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_3_10_4  (
            .in0(N__20213),
            .in1(N__21959),
            .in2(N__21941),
            .in3(N__20807),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_3_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_3_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_3_10_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_3_10_5  (
            .in0(N__20903),
            .in1(N__20801),
            .in2(N__20264),
            .in3(N__20600),
            .lcout(\current_shift_inst.PI_CTRL.N_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_3_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_3_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_3_11_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_3_11_4  (
            .in0(_gnd_net_),
            .in1(N__22142),
            .in2(_gnd_net_),
            .in3(N__22160),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_3_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_3_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_3_11_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_3_11_7  (
            .in0(N__20771),
            .in1(N__20813),
            .in2(N__20795),
            .in3(N__20783),
            .lcout(\current_shift_inst.PI_CTRL.N_118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_12_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_12_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_12_0  (
            .in0(_gnd_net_),
            .in1(N__20312),
            .in2(N__20156),
            .in3(N__20878),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_3_12_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_12_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_12_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_12_1  (
            .in0(N__20856),
            .in1(N__20303),
            .in2(N__20147),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_12_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_12_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_12_2  (
            .in0(_gnd_net_),
            .in1(N__20135),
            .in2(N__20915),
            .in3(N__20836),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_12_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_12_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_12_3  (
            .in0(_gnd_net_),
            .in1(N__21656),
            .in2(N__20129),
            .in3(N__21111),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_12_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_12_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_12_4  (
            .in0(_gnd_net_),
            .in1(N__20399),
            .in2(N__20498),
            .in3(N__21090),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_12_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_12_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_12_5  (
            .in0(_gnd_net_),
            .in1(N__20378),
            .in2(N__20393),
            .in3(N__21069),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_12_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_12_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_12_6  (
            .in0(_gnd_net_),
            .in1(N__20486),
            .in2(N__20372),
            .in3(N__21048),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_12_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_12_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_12_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_12_7  (
            .in0(N__21027),
            .in1(N__20588),
            .in2(N__20363),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_13_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_13_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_13_0  (
            .in0(_gnd_net_),
            .in1(N__21614),
            .in2(N__20354),
            .in3(N__21006),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_3_13_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_13_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_13_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_13_1  (
            .in0(_gnd_net_),
            .in1(N__21665),
            .in2(N__20345),
            .in3(N__20934),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_3_13_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_3_13_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_3_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_3_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20336),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47860),
            .ce(),
            .sr(N__47396));
    defparam \pwm_generator_inst.threshold_0_LC_3_14_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_0_LC_3_14_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_0_LC_3_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_0_LC_3_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20417),
            .lcout(\pwm_generator_inst.thresholdZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47847),
            .ce(),
            .sr(N__47401));
    defparam \pwm_generator_inst.threshold_1_LC_3_14_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_1_LC_3_14_3 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_1_LC_3_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_1_LC_3_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20570),
            .lcout(\pwm_generator_inst.thresholdZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47847),
            .ce(),
            .sr(N__47401));
    defparam \pwm_generator_inst.threshold_4_LC_3_14_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_4_LC_3_14_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_4_LC_3_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_4_LC_3_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20579),
            .lcout(\pwm_generator_inst.thresholdZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47847),
            .ce(),
            .sr(N__47401));
    defparam \pwm_generator_inst.threshold_6_LC_3_14_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_6_LC_3_14_6 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_6_LC_3_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_6_LC_3_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20408),
            .lcout(\pwm_generator_inst.thresholdZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47847),
            .ce(),
            .sr(N__47401));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_3_15_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_3_15_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_3_15_2 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_3_15_2  (
            .in0(N__20477),
            .in1(N__20453),
            .in2(N__20429),
            .in3(N__21167),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_3_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_3_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_3_15_4 .LUT_INIT=16'b0011001100110010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_14_LC_3_15_4  (
            .in0(N__27162),
            .in1(N__27347),
            .in2(N__27431),
            .in3(N__24461),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47839),
            .ce(N__24365),
            .sr(N__47407));
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_3_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_3_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_3_15_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_10_LC_3_15_5  (
            .in0(N__27344),
            .in1(N__27163),
            .in2(N__27539),
            .in3(N__24469),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47839),
            .ce(N__24365),
            .sr(N__47407));
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_3_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_3_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_3_15_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_11_LC_3_15_6  (
            .in0(N__27161),
            .in1(N__27346),
            .in2(N__31256),
            .in3(N__24460),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47839),
            .ce(N__24365),
            .sr(N__47407));
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_3_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_3_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_3_15_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_12_LC_3_15_7  (
            .in0(N__27345),
            .in1(N__27164),
            .in2(N__27470),
            .in3(N__24470),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47839),
            .ce(N__24365),
            .sr(N__47407));
    defparam \pwm_generator_inst.threshold_ACC_0_LC_3_16_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_0_LC_3_16_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_0_LC_3_16_0 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_0_LC_3_16_0  (
            .in0(N__21582),
            .in1(N__20552),
            .in2(N__21434),
            .in3(N__21512),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47831),
            .ce(),
            .sr(N__47414));
    defparam \pwm_generator_inst.threshold_ACC_6_LC_3_16_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_6_LC_3_16_1 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_6_LC_3_16_1 .LUT_INIT=16'b1101110011011111;
    LogicCell40 \pwm_generator_inst.threshold_ACC_6_LC_3_16_1  (
            .in0(N__21515),
            .in1(N__20732),
            .in2(N__21437),
            .in3(N__21585),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47831),
            .ce(),
            .sr(N__47414));
    defparam \pwm_generator_inst.threshold_ACC_7_LC_3_16_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_7_LC_3_16_3 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_7_LC_3_16_3 .LUT_INIT=16'b1101110011011111;
    LogicCell40 \pwm_generator_inst.threshold_ACC_7_LC_3_16_3  (
            .in0(N__21516),
            .in1(N__20714),
            .in2(N__21438),
            .in3(N__21586),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47831),
            .ce(),
            .sr(N__47414));
    defparam \pwm_generator_inst.threshold_7_LC_3_16_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_7_LC_3_16_5 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_7_LC_3_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_7_LC_3_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20594),
            .lcout(\pwm_generator_inst.thresholdZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47831),
            .ce(),
            .sr(N__47414));
    defparam \pwm_generator_inst.threshold_ACC_4_LC_3_16_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_4_LC_3_16_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_4_LC_3_16_6 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_4_LC_3_16_6  (
            .in0(N__21584),
            .in1(N__20507),
            .in2(N__21435),
            .in3(N__21514),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47831),
            .ce(),
            .sr(N__47414));
    defparam \pwm_generator_inst.threshold_ACC_1_LC_3_16_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_1_LC_3_16_7 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_1_LC_3_16_7 .LUT_INIT=16'b1101110011011111;
    LogicCell40 \pwm_generator_inst.threshold_ACC_1_LC_3_16_7  (
            .in0(N__21513),
            .in1(N__20540),
            .in2(N__21436),
            .in3(N__21583),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47831),
            .ce(),
            .sr(N__47414));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_17_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_17_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_17_0  (
            .in0(_gnd_net_),
            .in1(N__20561),
            .in2(N__21208),
            .in3(N__21201),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_3_17_0_),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_17_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_17_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_17_1  (
            .in0(_gnd_net_),
            .in1(N__20546),
            .in2(_gnd_net_),
            .in3(N__20534),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_0 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_17_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_17_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_17_2  (
            .in0(_gnd_net_),
            .in1(N__20531),
            .in2(_gnd_net_),
            .in3(N__20522),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_1 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_17_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_17_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_17_3  (
            .in0(_gnd_net_),
            .in1(N__21119),
            .in2(_gnd_net_),
            .in3(N__20519),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_2 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_17_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_17_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_17_4  (
            .in0(_gnd_net_),
            .in1(N__20516),
            .in2(_gnd_net_),
            .in3(N__20501),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_3 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_17_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_17_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_17_5  (
            .in0(_gnd_net_),
            .in1(N__20765),
            .in2(_gnd_net_),
            .in3(N__20744),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_4 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_17_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_17_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_17_6  (
            .in0(_gnd_net_),
            .in1(N__20741),
            .in2(_gnd_net_),
            .in3(N__20726),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_5 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_17_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_17_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_17_7  (
            .in0(_gnd_net_),
            .in1(N__20723),
            .in2(_gnd_net_),
            .in3(N__20708),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_6 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_18_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_18_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_18_0  (
            .in0(_gnd_net_),
            .in1(N__20633),
            .in2(_gnd_net_),
            .in3(N__20705),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(bfn_3_18_0_),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_18_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_18_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_18_1 .LUT_INIT=16'b1001010101101010;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_18_1  (
            .in0(N__20702),
            .in1(N__20690),
            .in2(N__21209),
            .in3(N__20684),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_3_18_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_3_18_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_3_18_5 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_3_18_5  (
            .in0(N__20681),
            .in1(N__21204),
            .in2(N__20663),
            .in3(N__20639),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_3_30_5.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_3_30_5.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_3_30_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_3_30_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20627),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_4_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_4_10_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_4_10_1  (
            .in0(N__22280),
            .in1(N__22334),
            .in2(N__22316),
            .in3(N__20777),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_10_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_10_3  (
            .in0(_gnd_net_),
            .in1(N__21934),
            .in2(_gnd_net_),
            .in3(N__21970),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_10_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_10_4  (
            .in0(N__21955),
            .in1(N__22312),
            .in2(N__20816),
            .in3(N__20897),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_10_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_10_5  (
            .in0(N__22298),
            .in1(N__21971),
            .in2(N__22178),
            .in3(N__21890),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_10_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_10_6  (
            .in0(N__21920),
            .in1(N__22067),
            .in2(N__22052),
            .in3(N__21905),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_11_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_11_0  (
            .in0(N__22330),
            .in1(N__22138),
            .in2(N__22276),
            .in3(N__22156),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_11_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_11_2  (
            .in0(_gnd_net_),
            .in1(N__22174),
            .in2(_gnd_net_),
            .in3(N__21889),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_11_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_11_3  (
            .in0(N__22079),
            .in1(N__22345),
            .in2(N__20786),
            .in3(N__22360),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_4_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_4_11_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_4_11_4  (
            .in0(_gnd_net_),
            .in1(N__22096),
            .in2(_gnd_net_),
            .in3(N__22078),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_11_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_11_5  (
            .in0(N__22123),
            .in1(N__21904),
            .in2(N__22112),
            .in3(N__21919),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_11_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_11_6  (
            .in0(N__22361),
            .in1(N__22111),
            .in2(N__22349),
            .in3(N__22124),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_11_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_11_7  (
            .in0(N__22294),
            .in1(N__22066),
            .in2(N__22097),
            .in3(N__22045),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_4_12_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_4_12_1 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \pwm_generator_inst.counter_RNISQD2_0_LC_4_12_1  (
            .in0(N__20835),
            .in1(N__20877),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_4_12_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_4_12_2 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_1_LC_4_12_2  (
            .in0(N__21091),
            .in1(N__20857),
            .in2(N__20891),
            .in3(N__21112),
            .lcout(\pwm_generator_inst.un1_counterlt9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_4_12_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_4_12_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIVDL3_9_LC_4_12_4  (
            .in0(N__20936),
            .in1(N__21008),
            .in2(_gnd_net_),
            .in3(N__21028),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto9_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_4_12_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_4_12_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_5_LC_4_12_5  (
            .in0(N__21050),
            .in1(N__21071),
            .in2(N__20888),
            .in3(N__20885),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_0_LC_4_13_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_4_13_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_4_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_4_13_0  (
            .in0(N__20981),
            .in1(N__20879),
            .in2(_gnd_net_),
            .in3(N__20861),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_4_13_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__47848),
            .ce(),
            .sr(N__47390));
    defparam \pwm_generator_inst.counter_1_LC_4_13_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_4_13_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_4_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_4_13_1  (
            .in0(N__20966),
            .in1(N__20858),
            .in2(_gnd_net_),
            .in3(N__20840),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__47848),
            .ce(),
            .sr(N__47390));
    defparam \pwm_generator_inst.counter_2_LC_4_13_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_4_13_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_4_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_4_13_2  (
            .in0(N__20982),
            .in1(N__20837),
            .in2(_gnd_net_),
            .in3(N__20819),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__47848),
            .ce(),
            .sr(N__47390));
    defparam \pwm_generator_inst.counter_3_LC_4_13_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_4_13_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_4_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_4_13_3  (
            .in0(N__20967),
            .in1(N__21113),
            .in2(_gnd_net_),
            .in3(N__21095),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__47848),
            .ce(),
            .sr(N__47390));
    defparam \pwm_generator_inst.counter_4_LC_4_13_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_4_13_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_4_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_4_13_4  (
            .in0(N__20983),
            .in1(N__21092),
            .in2(_gnd_net_),
            .in3(N__21074),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__47848),
            .ce(),
            .sr(N__47390));
    defparam \pwm_generator_inst.counter_5_LC_4_13_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_4_13_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_4_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_4_13_5  (
            .in0(N__20968),
            .in1(N__21070),
            .in2(_gnd_net_),
            .in3(N__21053),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__47848),
            .ce(),
            .sr(N__47390));
    defparam \pwm_generator_inst.counter_6_LC_4_13_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_4_13_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_4_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_4_13_6  (
            .in0(N__20984),
            .in1(N__21049),
            .in2(_gnd_net_),
            .in3(N__21032),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__47848),
            .ce(),
            .sr(N__47390));
    defparam \pwm_generator_inst.counter_7_LC_4_13_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_4_13_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_4_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_4_13_7  (
            .in0(N__20969),
            .in1(N__21029),
            .in2(_gnd_net_),
            .in3(N__21011),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__47848),
            .ce(),
            .sr(N__47390));
    defparam \pwm_generator_inst.counter_8_LC_4_14_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_4_14_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_4_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_4_14_0  (
            .in0(N__20980),
            .in1(N__21007),
            .in2(_gnd_net_),
            .in3(N__20987),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_4_14_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__47840),
            .ce(),
            .sr(N__47397));
    defparam \pwm_generator_inst.counter_9_LC_4_14_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_4_14_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_4_14_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \pwm_generator_inst.counter_9_LC_4_14_1  (
            .in0(N__20935),
            .in1(N__20979),
            .in2(_gnd_net_),
            .in3(N__20939),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47840),
            .ce(),
            .sr(N__47397));
    defparam \pwm_generator_inst.threshold_2_LC_4_14_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_2_LC_4_14_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_2_LC_4_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_2_LC_4_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21635),
            .lcout(\pwm_generator_inst.thresholdZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47840),
            .ce(),
            .sr(N__47397));
    defparam \pwm_generator_inst.threshold_9_LC_4_15_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_9_LC_4_15_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_9_LC_4_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_9_LC_4_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21275),
            .lcout(\pwm_generator_inst.thresholdZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47832),
            .ce(),
            .sr(N__47402));
    defparam \pwm_generator_inst.threshold_3_LC_4_16_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_3_LC_4_16_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_3_LC_4_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_3_LC_4_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21620),
            .lcout(\pwm_generator_inst.thresholdZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47826),
            .ce(),
            .sr(N__47408));
    defparam \pwm_generator_inst.threshold_ACC_2_LC_4_16_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_2_LC_4_16_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_2_LC_4_16_2 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_2_LC_4_16_2  (
            .in0(N__21589),
            .in1(N__21464),
            .in2(N__21644),
            .in3(N__21527),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47826),
            .ce(),
            .sr(N__47408));
    defparam \pwm_generator_inst.threshold_ACC_3_LC_4_16_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_3_LC_4_16_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_3_LC_4_16_3 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_3_LC_4_16_3  (
            .in0(N__21528),
            .in1(N__21590),
            .in2(N__21470),
            .in3(N__21626),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47826),
            .ce(),
            .sr(N__47408));
    defparam \pwm_generator_inst.threshold_8_LC_4_16_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_8_LC_4_16_6 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_8_LC_4_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_8_LC_4_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21596),
            .lcout(\pwm_generator_inst.thresholdZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47826),
            .ce(),
            .sr(N__47408));
    defparam \pwm_generator_inst.threshold_ACC_8_LC_4_17_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_8_LC_4_17_0 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_8_LC_4_17_0 .LUT_INIT=16'b1100110111111101;
    LogicCell40 \pwm_generator_inst.threshold_ACC_8_LC_4_17_0  (
            .in0(N__21587),
            .in1(N__21602),
            .in2(N__21469),
            .in3(N__21529),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47820),
            .ce(),
            .sr(N__47415));
    defparam \pwm_generator_inst.threshold_ACC_9_LC_4_17_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_9_LC_4_17_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_9_LC_4_17_2 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_9_LC_4_17_2  (
            .in0(N__21588),
            .in1(N__21530),
            .in2(N__21468),
            .in3(N__21281),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47820),
            .ce(),
            .sr(N__47415));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_4_17_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_4_17_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_4_17_7 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_4_17_7  (
            .in0(N__21266),
            .in1(N__21257),
            .in2(N__21230),
            .in3(N__21197),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_4_3.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_4_3.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_4_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D1_LC_5_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21875),
            .lcout(il_max_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47875),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_9_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_9_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_9_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_9_0  (
            .in0(_gnd_net_),
            .in1(N__28358),
            .in2(N__23579),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(bfn_5_9_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .clk(N__47868),
            .ce(),
            .sr(N__47352));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_9_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_9_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_9_1  (
            .in0(_gnd_net_),
            .in1(N__28337),
            .in2(N__30569),
            .in3(N__21848),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .clk(N__47868),
            .ce(),
            .sr(N__47352));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_9_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_9_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_9_2  (
            .in0(_gnd_net_),
            .in1(N__26176),
            .in2(N__30803),
            .in3(N__21836),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .clk(N__47868),
            .ce(),
            .sr(N__47352));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_9_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_9_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_9_3  (
            .in0(_gnd_net_),
            .in1(N__22478),
            .in2(N__25714),
            .in3(N__21809),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .clk(N__47868),
            .ce(),
            .sr(N__47352));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_9_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_9_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_9_4  (
            .in0(_gnd_net_),
            .in1(N__25754),
            .in2(N__28604),
            .in3(N__21764),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__47868),
            .ce(),
            .sr(N__47352));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_9_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_9_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_9_5  (
            .in0(_gnd_net_),
            .in1(N__25795),
            .in2(N__28589),
            .in3(N__21734),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__47868),
            .ce(),
            .sr(N__47352));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_9_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_9_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_9_6  (
            .in0(_gnd_net_),
            .in1(N__28426),
            .in2(N__22406),
            .in3(N__21701),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__47868),
            .ce(),
            .sr(N__47352));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_9_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_9_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_9_7  (
            .in0(_gnd_net_),
            .in1(N__28346),
            .in2(N__22769),
            .in3(N__21668),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__47868),
            .ce(),
            .sr(N__47352));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(N__22499),
            .in2(N__30782),
            .in3(N__22004),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(bfn_5_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__47865),
            .ce(),
            .sr(N__47363));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_10_1  (
            .in0(_gnd_net_),
            .in1(N__25948),
            .in2(N__22490),
            .in3(N__21974),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__47865),
            .ce(),
            .sr(N__47363));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_10_2  (
            .in0(_gnd_net_),
            .in1(N__22967),
            .in2(N__26015),
            .in3(N__21962),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__47865),
            .ce(),
            .sr(N__47363));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_10_3  (
            .in0(_gnd_net_),
            .in1(N__22466),
            .in2(N__25510),
            .in3(N__21944),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__47865),
            .ce(),
            .sr(N__47363));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_10_4  (
            .in0(_gnd_net_),
            .in1(N__22925),
            .in2(N__28490),
            .in3(N__21923),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__47865),
            .ce(),
            .sr(N__47363));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_10_5  (
            .in0(_gnd_net_),
            .in1(N__40546),
            .in2(N__22951),
            .in3(N__21908),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__47865),
            .ce(),
            .sr(N__47363));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_10_6  (
            .in0(_gnd_net_),
            .in1(N__22929),
            .in2(N__25565),
            .in3(N__21893),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__47865),
            .ce(),
            .sr(N__47363));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_10_7  (
            .in0(_gnd_net_),
            .in1(N__24047),
            .in2(N__22952),
            .in3(N__21878),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__47865),
            .ce(),
            .sr(N__47363));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_11_0  (
            .in0(_gnd_net_),
            .in1(N__22892),
            .in2(N__25381),
            .in3(N__22163),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(bfn_5_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__47861),
            .ce(),
            .sr(N__47372));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(N__25855),
            .in2(N__22933),
            .in3(N__22145),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__47861),
            .ce(),
            .sr(N__47372));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_11_2  (
            .in0(_gnd_net_),
            .in1(N__22896),
            .in2(N__25907),
            .in3(N__22127),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__47861),
            .ce(),
            .sr(N__47372));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(N__27599),
            .in2(N__22934),
            .in3(N__22115),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__47861),
            .ce(),
            .sr(N__47372));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_11_4  (
            .in0(_gnd_net_),
            .in1(N__22900),
            .in2(N__26237),
            .in3(N__22100),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__47861),
            .ce(),
            .sr(N__47372));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_11_5  (
            .in0(_gnd_net_),
            .in1(N__30697),
            .in2(N__22935),
            .in3(N__22082),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__47861),
            .ce(),
            .sr(N__47372));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_11_6  (
            .in0(_gnd_net_),
            .in1(N__22904),
            .in2(N__26072),
            .in3(N__22070),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__47861),
            .ce(),
            .sr(N__47372));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(N__26359),
            .in2(N__22936),
            .in3(N__22055),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__47861),
            .ce(),
            .sr(N__47372));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_12_0  (
            .in0(_gnd_net_),
            .in1(N__22937),
            .in2(N__30500),
            .in3(N__22034),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(bfn_5_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__47849),
            .ce(),
            .sr(N__47378));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(N__26300),
            .in2(N__22953),
            .in3(N__22352),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__47849),
            .ce(),
            .sr(N__47378));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(N__22941),
            .in2(N__26126),
            .in3(N__22337),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__47849),
            .ce(),
            .sr(N__47378));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(N__29272),
            .in2(N__22954),
            .in3(N__22319),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__47849),
            .ce(),
            .sr(N__47378));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(N__22945),
            .in2(N__24098),
            .in3(N__22301),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__47849),
            .ce(),
            .sr(N__47378));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_12_5  (
            .in0(_gnd_net_),
            .in1(N__24135),
            .in2(N__22955),
            .in3(N__22283),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__47849),
            .ce(),
            .sr(N__47378));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_12_6  (
            .in0(_gnd_net_),
            .in1(N__22949),
            .in2(N__40613),
            .in3(N__22259),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__47849),
            .ce(),
            .sr(N__47378));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_12_7  (
            .in0(N__22950),
            .in1(N__28305),
            .in2(_gnd_net_),
            .in3(N__22256),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47849),
            .ce(),
            .sr(N__47378));
    defparam SB_DFF_inst_PH2_MAX_D2_LC_7_6_6.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_7_6_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_7_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D2_LC_7_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22190),
            .lcout(il_max_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47869),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_7_7_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_7_7_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_7_7_2  (
            .in0(N__26364),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDA7M_0_15_LC_7_7_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDA7M_0_15_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDA7M_0_15_LC_7_7_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDA7M_0_15_LC_7_7_3  (
            .in0(N__25890),
            .in1(N__25840),
            .in2(N__24041),
            .in3(N__26226),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_29_LC_7_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_29_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_29_LC_7_7_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_29_LC_7_7_4  (
            .in0(N__26363),
            .in1(N__25380),
            .in2(N__26014),
            .in3(N__24136),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_29_LC_7_7_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_29_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_29_LC_7_7_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICA8M_29_LC_7_7_7  (
            .in0(N__25379),
            .in1(N__26006),
            .in2(N__24140),
            .in3(N__26365),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC4P2_19_LC_7_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC4P2_19_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC4P2_19_LC_7_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIGC4P2_19_LC_7_8_0  (
            .in0(N__22433),
            .in1(N__22814),
            .in2(N__25406),
            .in3(N__22391),
            .lcout(\current_shift_inst.PI_CTRL.N_74_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNID9B11_22_LC_7_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID9B11_22_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID9B11_22_LC_7_8_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNID9B11_22_LC_7_8_2  (
            .in0(N__26054),
            .in1(N__25509),
            .in2(_gnd_net_),
            .in3(N__22382),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_12_LC_7_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_12_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_12_LC_7_8_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_12_LC_7_8_3  (
            .in0(N__25421),
            .in1(N__22376),
            .in2(N__22370),
            .in3(N__22412),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_4_LC_7_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_4_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_4_LC_7_8_4 .LUT_INIT=16'b1111000000100000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIC35V7_4_LC_7_8_4  (
            .in0(N__22427),
            .in1(N__25750),
            .in2(N__22367),
            .in3(N__22451),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_75_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIE7HME_11_LC_7_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIE7HME_11_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIE7HME_11_LC_7_8_5 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIE7HME_11_LC_7_8_5  (
            .in0(N__25655),
            .in1(N__22439),
            .in2(N__22364),
            .in3(N__22831),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_7_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_7_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_7_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26005),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDAC11_11_LC_7_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDAC11_11_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDAC11_11_LC_7_8_7 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDAC11_11_LC_7_8_7  (
            .in0(N__22846),
            .in1(_gnd_net_),
            .in2(N__25511),
            .in3(N__28317),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFE9M_19_LC_7_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFE9M_19_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFE9M_19_LC_7_9_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFE9M_19_LC_7_9_1  (
            .in0(N__30475),
            .in1(N__30679),
            .in2(N__27596),
            .in3(N__26102),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_28_LC_7_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_28_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_28_LC_7_9_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIMMAM_28_LC_7_9_2  (
            .in0(N__26101),
            .in1(N__24096),
            .in2(N__29271),
            .in3(N__26279),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQB1L1_0_LC_7_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQB1L1_0_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQB1L1_0_LC_7_9_3 .LUT_INIT=16'b0101010101010111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIQB1L1_0_LC_7_9_3  (
            .in0(N__25713),
            .in1(N__30568),
            .in2(N__26180),
            .in3(N__23571),
            .lcout(\current_shift_inst.PI_CTRL.N_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDA7M_15_LC_7_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDA7M_15_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDA7M_15_LC_7_9_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDA7M_15_LC_7_9_4  (
            .in0(N__25889),
            .in1(N__25842),
            .in2(N__24040),
            .in3(N__26215),
            .lcout(\current_shift_inst.PI_CTRL.N_74_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_7_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_7_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_7_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29263),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBB5B_28_LC_7_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBB5B_28_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBB5B_28_LC_7_9_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIBB5B_28_LC_7_9_6  (
            .in0(_gnd_net_),
            .in1(N__24097),
            .in2(_gnd_net_),
            .in3(N__26278),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI01LC1_30_LC_7_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI01LC1_30_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI01LC1_30_LC_7_9_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI01LC1_30_LC_7_9_7  (
            .in0(N__40601),
            .in1(N__29264),
            .in2(N__22421),
            .in3(N__22418),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_7_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_7_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_7_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_7_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30869),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47850),
            .ce(),
            .sr(N__47341));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_7_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_7_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_7_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31094),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47850),
            .ce(),
            .sr(N__47341));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_7_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_7_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_7_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_7_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31061),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47850),
            .ce(),
            .sr(N__47341));
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_7_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_7_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_7_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_3_LC_7_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30947),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47850),
            .ce(),
            .sr(N__47341));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_7_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_7_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_7_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_7_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31133),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47850),
            .ce(),
            .sr(N__47341));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_7_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_7_11_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(N__22761),
            .in2(_gnd_net_),
            .in3(N__25785),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_7_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_7_11_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_7_11_2  (
            .in0(N__22762),
            .in1(N__30768),
            .in2(N__28419),
            .in3(N__25935),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_7_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_7_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25934),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_7_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_7_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_7_11_7 .LUT_INIT=16'b0011101100001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_7_11_7  (
            .in0(N__28269),
            .in1(N__23882),
            .in2(N__28152),
            .in3(N__27977),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47841),
            .ce(),
            .sr(N__47353));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_7_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_7_12_0 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_7_12_0  (
            .in0(N__25936),
            .in1(N__22457),
            .in2(N__30781),
            .in3(N__28415),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_7_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_7_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_7_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23572),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_7_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_7_12_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_7_12_3  (
            .in0(N__33678),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28839),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_7_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_7_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_7_12_6  (
            .in0(N__28974),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33677),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_1_c_inv_LC_7_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_1_c_inv_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_1_c_inv_LC_7_13_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_1_c_inv_LC_7_13_0  (
            .in0(N__23343),
            .in1(N__23441),
            .in2(N__22553),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_2_c_inv_LC_7_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_2_c_inv_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_2_c_inv_LC_7_13_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_2_c_inv_LC_7_13_1  (
            .in0(N__23092),
            .in1(N__23387),
            .in2(N__22544),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_3_c_inv_LC_7_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_3_c_inv_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_3_c_inv_LC_7_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_3_c_inv_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(N__23453),
            .in2(N__22535),
            .in3(N__23074),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_4_c_inv_LC_7_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_4_c_inv_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_4_c_inv_LC_7_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_4_c_inv_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(N__23375),
            .in2(N__22526),
            .in3(N__23059),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_5_c_inv_LC_7_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_5_c_inv_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_5_c_inv_LC_7_13_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_5_c_inv_LC_7_13_4  (
            .in0(N__23044),
            .in1(N__23477),
            .in2(N__22517),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_6_c_inv_LC_7_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_6_c_inv_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_6_c_inv_LC_7_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_6_c_inv_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(N__23399),
            .in2(N__22508),
            .in3(N__23029),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_7_c_inv_LC_7_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_7_c_inv_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_7_c_inv_LC_7_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_7_c_inv_LC_7_13_6  (
            .in0(_gnd_net_),
            .in1(N__24377),
            .in2(N__22670),
            .in3(N__23014),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_8_c_inv_LC_7_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_8_c_inv_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_8_c_inv_LC_7_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_8_c_inv_LC_7_13_7  (
            .in0(_gnd_net_),
            .in1(N__23465),
            .in2(N__22661),
            .in3(N__22999),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_9_c_inv_LC_7_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_9_c_inv_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_9_c_inv_LC_7_14_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_9_c_inv_LC_7_14_0  (
            .in0(N__22981),
            .in1(N__24245),
            .in2(N__22652),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_7_14_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_10_c_inv_LC_7_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_10_c_inv_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_10_c_inv_LC_7_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_10_c_inv_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(N__22643),
            .in2(N__22631),
            .in3(N__23227),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_11_c_inv_LC_7_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_11_c_inv_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_11_c_inv_LC_7_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_11_c_inv_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(N__22622),
            .in2(N__22610),
            .in3(N__23212),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_12_c_inv_LC_7_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_12_c_inv_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_12_c_inv_LC_7_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_12_c_inv_LC_7_14_3  (
            .in0(_gnd_net_),
            .in1(N__22601),
            .in2(N__22589),
            .in3(N__23197),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_13_c_inv_LC_7_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_13_c_inv_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_13_c_inv_LC_7_14_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_13_c_inv_LC_7_14_4  (
            .in0(N__23182),
            .in1(N__22580),
            .in2(N__24236),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_14_c_inv_LC_7_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_14_c_inv_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_14_c_inv_LC_7_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_14_c_inv_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(N__22574),
            .in2(N__22562),
            .in3(N__23167),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_15_c_inv_LC_7_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_15_c_inv_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_15_c_inv_LC_7_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_15_c_inv_LC_7_14_6  (
            .in0(_gnd_net_),
            .in1(N__24179),
            .in2(N__22721),
            .in3(N__23152),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_16_c_inv_LC_7_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_16_c_inv_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_16_c_inv_LC_7_14_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_16_c_inv_LC_7_14_7  (
            .in0(N__23137),
            .in1(N__24188),
            .in2(N__22709),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_17_c_inv_LC_7_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_17_c_inv_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_17_c_inv_LC_7_15_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_17_c_inv_LC_7_15_0  (
            .in0(N__23122),
            .in1(N__24200),
            .in2(N__22700),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_18_c_inv_LC_7_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_18_c_inv_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_18_c_inv_LC_7_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_18_c_inv_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(N__24212),
            .in2(N__22691),
            .in3(N__23107),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_inv_LC_7_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_inv_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_inv_LC_7_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_inv_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(N__24224),
            .in2(N__22682),
            .in3(N__23359),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_LUT4_0_LC_7_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_LUT4_0_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_LUT4_0_LC_7_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_LUT4_0_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22673),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNI5B6O_0_LC_7_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNI5B6O_0_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNI5B6O_0_LC_7_15_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNI5B6O_0_LC_7_15_5  (
            .in0(N__36284),
            .in1(N__36252),
            .in2(_gnd_net_),
            .in3(N__23300),
            .lcout(\phase_controller_inst1.stoper_hc.running_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.running_LC_7_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_LC_7_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.running_LC_7_16_1 .LUT_INIT=16'b1010101000101110;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_LC_7_16_1  (
            .in0(N__23264),
            .in1(N__23249),
            .in2(N__36300),
            .in3(N__23321),
            .lcout(\phase_controller_inst1.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47809),
            .ce(),
            .sr(N__47391));
    defparam \phase_controller_inst2.start_timer_hc_RNO_1_LC_7_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_RNO_1_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_hc_RNO_1_LC_7_16_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_RNO_1_LC_7_16_2  (
            .in0(_gnd_net_),
            .in1(N__32419),
            .in2(_gnd_net_),
            .in3(N__32067),
            .lcout(),
            .ltout(\phase_controller_inst2.start_timer_hc_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_hc_LC_7_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_LC_7_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_hc_LC_7_16_3 .LUT_INIT=16'b1111000111110000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_LC_7_16_3  (
            .in0(N__34827),
            .in1(N__22730),
            .in2(N__22733),
            .in3(N__27738),
            .lcout(\phase_controller_inst2.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47809),
            .ce(),
            .sr(N__47391));
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_7_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_7_16_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_RNO_0_LC_7_16_4  (
            .in0(_gnd_net_),
            .in1(N__32138),
            .in2(_gnd_net_),
            .in3(N__32112),
            .lcout(\phase_controller_inst2.start_timer_hc_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_2_LC_7_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_2_LC_7_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_2_LC_7_16_5 .LUT_INIT=16'b1111001000100010;
    LogicCell40 \phase_controller_inst2.state_2_LC_7_16_5  (
            .in0(N__32139),
            .in1(N__32113),
            .in2(N__32074),
            .in3(N__32420),
            .lcout(\phase_controller_inst2.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47809),
            .ce(),
            .sr(N__47391));
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_7_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_7_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_7_16_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_LC_7_16_6  (
            .in0(N__36253),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47809),
            .ce(),
            .sr(N__47391));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_7_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_7_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_7_18_0 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_7_18_0  (
            .in0(N__22793),
            .in1(N__27015),
            .in2(N__22808),
            .in3(N__24801),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47798),
            .ce(),
            .sr(N__47403));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNINJB21_LC_7_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNINJB21_LC_7_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNINJB21_LC_7_18_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNINJB21_LC_7_18_1  (
            .in0(_gnd_net_),
            .in1(N__22792),
            .in2(_gnd_net_),
            .in3(N__22804),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNINJBZ0Z21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_7_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_7_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_7_18_2 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_7_18_2  (
            .in0(N__34598),
            .in1(N__34625),
            .in2(N__35742),
            .in3(N__42102),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47798),
            .ce(),
            .sr(N__47403));
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_7_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_7_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_7_19_1 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_LC_7_19_1  (
            .in0(N__27698),
            .in1(N__32111),
            .in2(N__27750),
            .in3(N__27653),
            .lcout(\phase_controller_inst2.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47793),
            .ce(),
            .sr(N__47409));
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_7_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_7_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_7_19_2 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_7_19_2  (
            .in0(N__27666),
            .in1(N__27696),
            .in2(_gnd_net_),
            .in3(N__27739),
            .lcout(\phase_controller_inst2.stoper_hc.un2_start_0 ),
            .ltout(\phase_controller_inst2.stoper_hc.un2_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.running_LC_7_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_LC_7_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.running_LC_7_19_3 .LUT_INIT=16'b1100110001011100;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_LC_7_19_3  (
            .in0(N__27699),
            .in1(N__27667),
            .in2(N__22724),
            .in3(N__27761),
            .lcout(\phase_controller_inst2.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47793),
            .ce(),
            .sr(N__47409));
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_7_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_7_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_7_19_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_LC_7_19_5  (
            .in0(N__27743),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47793),
            .ce(),
            .sr(N__47409));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNIV5S7_LC_7_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNIV5S7_LC_7_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNIV5S7_LC_7_19_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNIV5S7_LC_7_19_6  (
            .in0(_gnd_net_),
            .in1(N__27697),
            .in2(_gnd_net_),
            .in3(N__27782),
            .lcout(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_7_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_7_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_7_19_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_7_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22796),
            .in3(N__22791),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_7_20_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_7_20_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_7_20_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_7_20_5  (
            .in0(_gnd_net_),
            .in1(N__27705),
            .in2(_gnd_net_),
            .in3(N__27749),
            .lcout(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_5_5.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_5_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_5_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH1_MAX_D1_LC_8_5_5 (
            .in0(N__22778),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_max_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47870),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_8_7_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_8_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_8_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25841),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGQQ01_11_LC_8_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGQQ01_11_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGQQ01_11_LC_8_8_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIGQQ01_11_LC_8_8_0  (
            .in0(N__22752),
            .in1(N__33774),
            .in2(N__31132),
            .in3(N__28712),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_8_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_8_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22751),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_8_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_8_8_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_8_8_2 .LUT_INIT=16'b0000110111011101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_8_8_2  (
            .in0(N__28316),
            .in1(N__28143),
            .in2(N__27979),
            .in3(N__23675),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47862),
            .ce(),
            .sr(N__47330));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_8_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_8_8_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_8_8_3 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_8_8_3  (
            .in0(N__23846),
            .in1(N__28314),
            .in2(N__28165),
            .in3(N__27935),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47862),
            .ce(),
            .sr(N__47330));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_8_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_8_8_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_8_8_5 .LUT_INIT=16'b0111010100110000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_8_8_5  (
            .in0(N__28145),
            .in1(N__23807),
            .in2(N__27980),
            .in3(N__28315),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47862),
            .ce(),
            .sr(N__47330));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_8_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_8_8_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_8_8_6 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_8_8_6  (
            .in0(N__28313),
            .in1(N__28144),
            .in2(N__27978),
            .in3(N__23786),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47862),
            .ce(),
            .sr(N__47330));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIJD8U_9_LC_8_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIJD8U_9_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIJD8U_9_LC_8_9_0 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIJD8U_9_LC_8_9_0  (
            .in0(N__25775),
            .in1(N__31057),
            .in2(N__33776),
            .in3(N__28742),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_8_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_8_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25774),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_8_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_8_9_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_8_9_2 .LUT_INIT=16'b0101111100010011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_8_9_2  (
            .in0(N__28002),
            .in1(N__28304),
            .in2(N__23726),
            .in3(N__28100),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47851),
            .ce(),
            .sr(N__47333));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_8_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_8_9_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_8_9_3 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_8_9_3  (
            .in0(N__28300),
            .in1(N__28003),
            .in2(N__28148),
            .in3(N__23774),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47851),
            .ce(),
            .sr(N__47333));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_8_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_8_9_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_8_9_4 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_8_9_4  (
            .in0(N__28000),
            .in1(N__28302),
            .in2(N__23756),
            .in3(N__28098),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47851),
            .ce(),
            .sr(N__47333));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_8_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_8_9_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_8_9_5 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_8_9_5  (
            .in0(N__28301),
            .in1(N__28004),
            .in2(N__28149),
            .in3(N__23981),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47851),
            .ce(),
            .sr(N__47333));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_8_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_8_9_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_8_9_6 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_8_9_6  (
            .in0(N__28001),
            .in1(N__28303),
            .in2(N__23969),
            .in3(N__28099),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47851),
            .ce(),
            .sr(N__47333));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBA9M_19_LC_8_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBA9M_19_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBA9M_19_LC_8_9_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIBA9M_19_LC_8_9_7  (
            .in0(N__30476),
            .in1(N__30680),
            .in2(N__27597),
            .in3(N__26053),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_11_LC_8_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_11_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_11_LC_8_10_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_11_LC_8_10_0  (
            .in0(N__22847),
            .in1(N__25490),
            .in2(N__22835),
            .in3(N__25654),
            .lcout(\current_shift_inst.PI_CTRL.N_103 ),
            .ltout(\current_shift_inst.PI_CTRL.N_103_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_8_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_8_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_8_10_1 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_8_10_1  (
            .in0(N__28296),
            .in1(N__27952),
            .in2(N__22817),
            .in3(N__23606),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47842),
            .ce(),
            .sr(N__47335));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_8_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_8_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25489),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_8_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_8_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_8_10_5 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_8_10_5  (
            .in0(N__28297),
            .in1(N__27953),
            .in2(N__28160),
            .in3(N__23936),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47842),
            .ce(),
            .sr(N__47335));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_8_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_8_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_8_10_6 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_8_10_6  (
            .in0(N__27951),
            .in1(N__28299),
            .in2(N__23927),
            .in3(N__28129),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47842),
            .ce(),
            .sr(N__47335));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_8_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_8_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_8_10_7 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_8_10_7  (
            .in0(N__28298),
            .in1(N__27954),
            .in2(N__28161),
            .in3(N__23903),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47842),
            .ce(),
            .sr(N__47335));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_8_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_8_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_8_11_0 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_8_11_0  (
            .in0(N__28265),
            .in1(N__27956),
            .in2(N__28147),
            .in3(N__23945),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47833),
            .ce(),
            .sr(N__47342));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_8_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_8_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_8_11_1 .LUT_INIT=16'b0000110010101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_8_11_1  (
            .in0(N__27955),
            .in1(N__28266),
            .in2(N__28150),
            .in3(N__24158),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47833),
            .ce(),
            .sr(N__47342));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_8_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_8_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_8_11_2 .LUT_INIT=16'b0011101100001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_8_11_2  (
            .in0(N__28264),
            .in1(N__23825),
            .in2(N__28146),
            .in3(N__27960),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47833),
            .ce(),
            .sr(N__47342));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_8_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_8_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_8_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31028),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47833),
            .ce(),
            .sr(N__47342));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_8_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_8_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_8_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33773),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47833),
            .ce(),
            .sr(N__47342));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_8_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_8_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_8_11_5 .LUT_INIT=16'b0101000111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_8_11_5  (
            .in0(N__23702),
            .in1(N__28267),
            .in2(N__28151),
            .in3(N__27961),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47833),
            .ce(),
            .sr(N__47342));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_8_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_8_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_8_11_7 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_8_11_7  (
            .in0(N__28101),
            .in1(N__28268),
            .in2(N__27996),
            .in3(N__23648),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47833),
            .ce(),
            .sr(N__47342));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_8_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_8_12_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_8_12_1  (
            .in0(N__28408),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_8_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_8_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_8_12_3 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_8_12_3  (
            .in0(N__28261),
            .in1(N__27983),
            .in2(N__28163),
            .in3(N__23870),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47827),
            .ce(),
            .sr(N__47354));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_8_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_8_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_8_12_4 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_8_12_4  (
            .in0(N__27981),
            .in1(N__28263),
            .in2(N__24170),
            .in3(N__28139),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47827),
            .ce(),
            .sr(N__47354));
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_8_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_8_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_8_12_5 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_31_LC_8_12_5  (
            .in0(N__28262),
            .in1(N__27984),
            .in2(N__28164),
            .in3(N__24146),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47827),
            .ce(),
            .sr(N__47354));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_8_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_8_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_8_12_7 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_8_12_7  (
            .in0(N__28260),
            .in1(N__27982),
            .in2(N__28162),
            .in3(N__23624),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47827),
            .ce(),
            .sr(N__47354));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_8_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_8_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(N__23309),
            .in2(N__23348),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_13_1  (
            .in0(N__24352),
            .in1(N__23093),
            .in2(_gnd_net_),
            .in3(N__23081),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__47821),
            .ce(),
            .sr(N__47364));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_13_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_13_2  (
            .in0(N__24323),
            .in1(N__23273),
            .in2(N__23078),
            .in3(N__23063),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__47821),
            .ce(),
            .sr(N__47364));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_13_3  (
            .in0(N__24353),
            .in1(N__23060),
            .in2(_gnd_net_),
            .in3(N__23048),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__47821),
            .ce(),
            .sr(N__47364));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_13_4  (
            .in0(N__24324),
            .in1(N__23045),
            .in2(_gnd_net_),
            .in3(N__23033),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__47821),
            .ce(),
            .sr(N__47364));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_13_5  (
            .in0(N__24354),
            .in1(N__23030),
            .in2(_gnd_net_),
            .in3(N__23018),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__47821),
            .ce(),
            .sr(N__47364));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_13_6  (
            .in0(N__24325),
            .in1(N__23015),
            .in2(_gnd_net_),
            .in3(N__23003),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__47821),
            .ce(),
            .sr(N__47364));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_13_7  (
            .in0(N__24355),
            .in1(N__23000),
            .in2(_gnd_net_),
            .in3(N__22985),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__47821),
            .ce(),
            .sr(N__47364));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_14_0  (
            .in0(N__24364),
            .in1(N__22982),
            .in2(_gnd_net_),
            .in3(N__22970),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__47816),
            .ce(),
            .sr(N__47373));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_14_1  (
            .in0(N__24326),
            .in1(N__23228),
            .in2(_gnd_net_),
            .in3(N__23216),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__47816),
            .ce(),
            .sr(N__47373));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_14_2  (
            .in0(N__24361),
            .in1(N__23213),
            .in2(_gnd_net_),
            .in3(N__23201),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__47816),
            .ce(),
            .sr(N__47373));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_14_3  (
            .in0(N__24327),
            .in1(N__23198),
            .in2(_gnd_net_),
            .in3(N__23186),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__47816),
            .ce(),
            .sr(N__47373));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_14_4  (
            .in0(N__24362),
            .in1(N__23183),
            .in2(_gnd_net_),
            .in3(N__23171),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__47816),
            .ce(),
            .sr(N__47373));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_14_5  (
            .in0(N__24328),
            .in1(N__23168),
            .in2(_gnd_net_),
            .in3(N__23156),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__47816),
            .ce(),
            .sr(N__47373));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_14_6  (
            .in0(N__24363),
            .in1(N__23153),
            .in2(_gnd_net_),
            .in3(N__23141),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__47816),
            .ce(),
            .sr(N__47373));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_14_7  (
            .in0(N__24329),
            .in1(N__23138),
            .in2(_gnd_net_),
            .in3(N__23126),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__47816),
            .ce(),
            .sr(N__47373));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_15_0  (
            .in0(N__24330),
            .in1(N__23123),
            .in2(_gnd_net_),
            .in3(N__23111),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_8_15_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__47810),
            .ce(),
            .sr(N__47379));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_15_1  (
            .in0(N__24360),
            .in1(N__23108),
            .in2(_gnd_net_),
            .in3(N__23096),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__47810),
            .ce(),
            .sr(N__47379));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_15_2  (
            .in0(N__24331),
            .in1(N__23360),
            .in2(_gnd_net_),
            .in3(N__23363),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47810),
            .ce(),
            .sr(N__47379));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_15_5 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_15_5  (
            .in0(N__23248),
            .in1(N__23288),
            .in2(N__23347),
            .in3(N__24332),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47810),
            .ce(),
            .sr(N__47379));
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_8_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_8_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_8_16_0 .LUT_INIT=16'b1111111111001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_3_LC_8_16_0  (
            .in0(N__24870),
            .in1(N__26550),
            .in2(N__24953),
            .in3(N__24406),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47803),
            .ce(N__27021),
            .sr(N__47387));
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_8_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_8_16_1 .LUT_INIT=16'b0000000010111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_8_16_1  (
            .in0(N__23263),
            .in1(N__36241),
            .in2(N__36293),
            .in3(N__23320),
            .lcout(\phase_controller_inst1.stoper_hc.un1_start_latched2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_8_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_8_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_8_16_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_8_16_3  (
            .in0(_gnd_net_),
            .in1(N__23246),
            .in2(_gnd_net_),
            .in3(N__23287),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNI5B6O_LC_8_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNI5B6O_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNI5B6O_LC_8_16_4 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNI5B6O_LC_8_16_4  (
            .in0(N__36240),
            .in1(N__36280),
            .in2(_gnd_net_),
            .in3(N__23299),
            .lcout(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNIQVTI1_LC_8_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNIQVTI1_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNIQVTI1_LC_8_16_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNIQVTI1_LC_8_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23276),
            .in3(N__23247),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNIQVTIZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_8_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_8_16_6 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_8_16_6  (
            .in0(N__36239),
            .in1(N__23262),
            .in2(_gnd_net_),
            .in3(N__36279),
            .lcout(\phase_controller_inst1.stoper_hc.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_8_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_8_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_8_17_0 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_6_LC_8_17_0  (
            .in0(N__24941),
            .in1(N__24871),
            .in2(N__24581),
            .in3(N__27297),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47799),
            .ce(N__27020),
            .sr(N__47392));
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_8_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_8_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_8_17_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_7_LC_8_17_1  (
            .in0(N__27293),
            .in1(N__26860),
            .in2(_gnd_net_),
            .in3(N__24943),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47799),
            .ce(N__27020),
            .sr(N__47392));
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_8_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_8_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_8_17_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_8_LC_8_17_3  (
            .in0(N__27294),
            .in1(N__26831),
            .in2(_gnd_net_),
            .in3(N__24944),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47799),
            .ce(N__27020),
            .sr(N__47392));
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_8_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_8_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_8_17_4 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_16_LC_8_17_4  (
            .in0(N__27149),
            .in1(N__27292),
            .in2(_gnd_net_),
            .in3(N__33940),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47799),
            .ce(N__27020),
            .sr(N__47392));
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_8_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_8_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_8_17_5 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_5_LC_8_17_5  (
            .in0(N__27295),
            .in1(N__24863),
            .in2(N__26798),
            .in3(N__24942),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47799),
            .ce(N__27020),
            .sr(N__47392));
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_8_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_8_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_8_17_6 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_18_LC_8_17_6  (
            .in0(N__26646),
            .in1(N__27150),
            .in2(_gnd_net_),
            .in3(N__27296),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47799),
            .ce(N__27020),
            .sr(N__47392));
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_8_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_8_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_8_17_7 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_1_LC_8_17_7  (
            .in0(N__24518),
            .in1(N__24535),
            .in2(N__24875),
            .in3(N__24388),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47799),
            .ce(N__27020),
            .sr(N__47392));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_8_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_8_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_8_18_0 .LUT_INIT=16'b0000000000100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_LC_8_18_0  (
            .in0(N__24580),
            .in1(N__24869),
            .in2(N__24951),
            .in3(N__27350),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47794),
            .ce(N__24356),
            .sr(N__47398));
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_8_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_8_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_8_18_1 .LUT_INIT=16'b0000001100000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_2_LC_8_18_1  (
            .in0(N__24867),
            .in1(N__24497),
            .in2(N__27359),
            .in3(N__24938),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47794),
            .ce(N__24356),
            .sr(N__47398));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_8_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_8_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_8_18_2 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_LC_8_18_2  (
            .in0(N__24866),
            .in1(N__26702),
            .in2(N__24950),
            .in3(N__27349),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47794),
            .ce(N__24356),
            .sr(N__47398));
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_8_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_8_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_8_18_3 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_5_LC_8_18_3  (
            .in0(N__27354),
            .in1(N__24940),
            .in2(N__26797),
            .in3(N__24865),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47794),
            .ce(N__24356),
            .sr(N__47398));
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_8_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_8_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_8_18_4 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_8_LC_8_18_4  (
            .in0(_gnd_net_),
            .in1(N__27348),
            .in2(N__24952),
            .in3(N__26827),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47794),
            .ce(N__24356),
            .sr(N__47398));
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_8_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_8_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_8_18_5 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_3_LC_8_18_5  (
            .in0(N__24868),
            .in1(N__24939),
            .in2(N__24407),
            .in3(N__26554),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47794),
            .ce(N__24356),
            .sr(N__47398));
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_8_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_8_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_8_18_6 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_1_LC_8_18_6  (
            .in0(N__24864),
            .in1(N__24389),
            .in2(N__24536),
            .in3(N__24517),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47794),
            .ce(N__24356),
            .sr(N__47398));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_8_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_8_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_8_18_7 .LUT_INIT=16'b0001000111011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_8_18_7  (
            .in0(N__40484),
            .in1(N__44077),
            .in2(_gnd_net_),
            .in3(N__40835),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_8_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_8_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_8_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_8_19_0  (
            .in0(_gnd_net_),
            .in1(N__23429),
            .in2(N__24805),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_19_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_8_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_8_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_8_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_8_19_1  (
            .in0(N__26960),
            .in1(N__24764),
            .in2(_gnd_net_),
            .in3(N__23423),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__47788),
            .ce(),
            .sr(N__47404));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_8_19_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_8_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_8_19_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_8_19_2  (
            .in0(N__26964),
            .in1(N__24743),
            .in2(N__23420),
            .in3(N__23408),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__47788),
            .ce(),
            .sr(N__47404));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_8_19_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_8_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_8_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_8_19_3  (
            .in0(N__26961),
            .in1(N__24706),
            .in2(_gnd_net_),
            .in3(N__23405),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__47788),
            .ce(),
            .sr(N__47404));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_8_19_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_8_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_8_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_8_19_4  (
            .in0(N__26965),
            .in1(N__24665),
            .in2(_gnd_net_),
            .in3(N__23402),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__47788),
            .ce(),
            .sr(N__47404));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_8_19_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_8_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_8_19_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_8_19_5  (
            .in0(N__26962),
            .in1(N__24644),
            .in2(_gnd_net_),
            .in3(N__23504),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__47788),
            .ce(),
            .sr(N__47404));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_8_19_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_8_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_8_19_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_8_19_6  (
            .in0(N__26966),
            .in1(N__24602),
            .in2(_gnd_net_),
            .in3(N__23501),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__47788),
            .ce(),
            .sr(N__47404));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_8_19_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_8_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_8_19_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_8_19_7  (
            .in0(N__26963),
            .in1(N__25159),
            .in2(_gnd_net_),
            .in3(N__23498),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__47788),
            .ce(),
            .sr(N__47404));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_8_20_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_8_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_8_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_8_20_0  (
            .in0(N__27009),
            .in1(N__25127),
            .in2(_gnd_net_),
            .in3(N__23495),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_8_20_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__47784),
            .ce(),
            .sr(N__47410));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_8_20_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_8_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_8_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_8_20_1  (
            .in0(N__26953),
            .in1(N__25100),
            .in2(_gnd_net_),
            .in3(N__23492),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__47784),
            .ce(),
            .sr(N__47410));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_8_20_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_8_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_8_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_8_20_2  (
            .in0(N__27006),
            .in1(N__25067),
            .in2(_gnd_net_),
            .in3(N__23489),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__47784),
            .ce(),
            .sr(N__47410));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_8_20_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_8_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_8_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_8_20_3  (
            .in0(N__26954),
            .in1(N__25034),
            .in2(_gnd_net_),
            .in3(N__23486),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__47784),
            .ce(),
            .sr(N__47410));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_8_20_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_8_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_8_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_8_20_4  (
            .in0(N__27007),
            .in1(N__25007),
            .in2(_gnd_net_),
            .in3(N__23483),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__47784),
            .ce(),
            .sr(N__47410));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_8_20_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_8_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_8_20_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_8_20_5  (
            .in0(N__26955),
            .in1(N__24974),
            .in2(_gnd_net_),
            .in3(N__23480),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__47784),
            .ce(),
            .sr(N__47410));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_8_20_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_8_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_8_20_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_8_20_6  (
            .in0(N__27008),
            .in1(N__25325),
            .in2(_gnd_net_),
            .in3(N__23519),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__47784),
            .ce(),
            .sr(N__47410));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_8_20_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_8_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_8_20_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_8_20_7  (
            .in0(N__26956),
            .in1(N__25298),
            .in2(_gnd_net_),
            .in3(N__23516),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__47784),
            .ce(),
            .sr(N__47410));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_8_21_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_8_21_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_8_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_8_21_0  (
            .in0(N__26957),
            .in1(N__25277),
            .in2(_gnd_net_),
            .in3(N__23513),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_8_21_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__47779),
            .ce(),
            .sr(N__47416));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_8_21_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_8_21_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_8_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_8_21_1  (
            .in0(N__26959),
            .in1(N__25244),
            .in2(_gnd_net_),
            .in3(N__23510),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__47779),
            .ce(),
            .sr(N__47416));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_8_21_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_8_21_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_8_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_8_21_2  (
            .in0(N__26958),
            .in1(N__25223),
            .in2(_gnd_net_),
            .in3(N__23507),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47779),
            .ce(),
            .sr(N__47416));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_9_7_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_9_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26225),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_9_7_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_9_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_9_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25687),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_9_7_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_9_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_9_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25378),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_9_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_9_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25546),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_9_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_9_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_9_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25888),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_9_7_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_9_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_9_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26121),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_9_7_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_9_7_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_9_7_7  (
            .in0(_gnd_net_),
            .in1(N__33377),
            .in2(_gnd_net_),
            .in3(N__33851),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_434_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_9_8_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_9_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(N__30514),
            .in2(N__30518),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_9_8_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_9_8_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_9_8_1 .LUT_INIT=16'b0010100010000010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_0_LC_9_8_1  (
            .in0(N__27975),
            .in1(N__25615),
            .in2(N__25592),
            .in3(N__23540),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ),
            .clk(N__47852),
            .ce(),
            .sr(N__47327));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_9_8_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_9_8_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_9_8_2 .LUT_INIT=16'b0010100010000010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_9_8_2  (
            .in0(N__27965),
            .in1(N__30527),
            .in2(N__28370),
            .in3(N__23537),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ),
            .clk(N__47852),
            .ce(),
            .sr(N__47327));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_9_8_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_9_8_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_9_8_3 .LUT_INIT=16'b0010100010000010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_9_8_3  (
            .in0(N__27976),
            .in1(N__26138),
            .in2(N__25574),
            .in3(N__23534),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ),
            .clk(N__47852),
            .ce(),
            .sr(N__47327));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_9_8_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_9_8_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_9_8_4 .LUT_INIT=16'b0111110111010111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_9_8_4  (
            .in0(N__27966),
            .in1(N__23531),
            .in2(N__25394),
            .in3(N__23525),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ),
            .clk(N__47852),
            .ce(),
            .sr(N__47327));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_9_8_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_9_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_9_8_5  (
            .in0(_gnd_net_),
            .in1(N__25178),
            .in2(N__25457),
            .in3(N__23522),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_9_8_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_9_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_9_8_6  (
            .in0(_gnd_net_),
            .in1(N__23744),
            .in2(N__23738),
            .in3(N__23717),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_9_8_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_9_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(N__23714),
            .in2(N__28382),
            .in3(N__23693),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_9_9_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_9_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__23690),
            .in2(N__23684),
            .in3(N__23666),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_9_9_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_9_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__30728),
            .in2(N__25583),
            .in3(N__23663),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_9_9_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_9_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__23660),
            .in2(N__25916),
            .in3(N__23639),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_9_9_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_9_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__23636),
            .in2(N__25970),
            .in3(N__23615),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_9_9_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_9_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__23612),
            .in2(N__25466),
            .in3(N__23600),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_9_9_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_9_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(N__25517),
            .in2(N__28442),
            .in3(N__23597),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_9_9_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_9_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__40502),
            .in2(N__25961),
            .in3(N__23861),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_9_9_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_9_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_9_9_7  (
            .in0(_gnd_net_),
            .in1(N__23858),
            .in2(N__25526),
            .in3(N__23849),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_9_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_9_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(N__24002),
            .in2(N__24059),
            .in3(N__23837),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(bfn_9_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_9_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_9_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__23834),
            .in2(N__25334),
            .in3(N__23819),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_9_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_9_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(N__23816),
            .in2(N__25817),
            .in3(N__23798),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_9_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_9_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(N__23795),
            .in2(N__25865),
            .in3(N__23777),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_9_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_9_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(N__28505),
            .in2(N__26246),
            .in3(N__23768),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_9_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_9_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(N__23765),
            .in2(N__26189),
            .in3(N__23747),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_9_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_9_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(N__30653),
            .in2(N__25805),
            .in3(N__23972),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_9_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_9_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(N__23993),
            .in2(N__26027),
            .in3(N__23960),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_9_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_9_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(N__23957),
            .in2(N__26327),
            .in3(N__23939),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_9_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_9_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_9_11_1  (
            .in0(_gnd_net_),
            .in1(N__30449),
            .in2(N__26315),
            .in3(N__23930),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_9_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_9_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(N__26258),
            .in2(N__25628),
            .in3(N__23918),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_9_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_9_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(N__26078),
            .in2(N__23915),
            .in3(N__23897),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_9_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_9_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(N__23894),
            .in2(N__29231),
            .in3(N__23873),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_9_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_9_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_9_11_5  (
            .in0(_gnd_net_),
            .in1(N__24065),
            .in2(N__33503),
            .in3(N__23864),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_9_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_9_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_9_11_6  (
            .in0(_gnd_net_),
            .in1(N__33501),
            .in2(N__24107),
            .in3(N__24161),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_9_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_9_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_9_11_7  (
            .in0(_gnd_net_),
            .in1(N__33502),
            .in2(N__40565),
            .in3(N__24152),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_9_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_9_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_9_12_0  (
            .in0(N__28233),
            .in1(N__33727),
            .in2(_gnd_net_),
            .in3(N__24149),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_9_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_9_12_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_9_12_1  (
            .in0(N__24126),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_9_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_9_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24084),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_9_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_9_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_9_12_4  (
            .in0(N__29013),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33725),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_9_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_9_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24045),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5I_LC_9_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5I_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5I_LC_9_12_6 .LUT_INIT=16'b0011111111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5I_LC_9_12_6  (
            .in0(N__24046),
            .in1(N__33726),
            .in2(N__28897),
            .in3(N__28871),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_9_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_9_12_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_9_12_7  (
            .in0(_gnd_net_),
            .in1(N__26061),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_9_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_9_13_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_9_13_0  (
            .in0(N__33743),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29108),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_9_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_9_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(N__28896),
            .in2(_gnd_net_),
            .in3(N__33742),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_9_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_9_13_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__36301),
            .in2(_gnd_net_),
            .in3(N__36254),
            .lcout(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_9_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_9_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_9_14_0 .LUT_INIT=16'b0000000011111110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_9_LC_9_14_0  (
            .in0(N__24449),
            .in1(N__27122),
            .in2(N__35816),
            .in3(N__24482),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47811),
            .ce(N__24336),
            .sr(N__47365));
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_9_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_9_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_9_14_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_13_LC_9_14_1  (
            .in0(N__27339),
            .in1(N__27114),
            .in2(N__27505),
            .in3(N__24450),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47811),
            .ce(N__24336),
            .sr(N__47365));
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_9_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_9_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_9_14_2 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_19_LC_9_14_2  (
            .in0(N__27111),
            .in1(N__26617),
            .in2(_gnd_net_),
            .in3(N__27342),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47811),
            .ce(N__24336),
            .sr(N__47365));
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_9_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_9_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_9_14_3 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_18_LC_9_14_3  (
            .in0(N__27337),
            .in1(N__26647),
            .in2(_gnd_net_),
            .in3(N__27115),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47811),
            .ce(N__24336),
            .sr(N__47365));
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_9_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_9_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_9_14_4 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_17_LC_9_14_4  (
            .in0(N__27110),
            .in1(N__27340),
            .in2(_gnd_net_),
            .in3(N__26675),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47811),
            .ce(N__24336),
            .sr(N__47365));
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_9_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_9_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_9_14_5 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_16_LC_9_14_5  (
            .in0(N__27336),
            .in1(N__27113),
            .in2(_gnd_net_),
            .in3(N__33939),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47811),
            .ce(N__24336),
            .sr(N__47365));
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_9_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_9_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_9_14_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_15_LC_9_14_6  (
            .in0(N__27112),
            .in1(N__27341),
            .in2(N__27836),
            .in3(N__27196),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47811),
            .ce(N__24336),
            .sr(N__47365));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_9_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_9_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_9_14_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_LC_9_14_7  (
            .in0(N__27338),
            .in1(N__26864),
            .in2(_gnd_net_),
            .in3(N__24945),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47811),
            .ce(N__24336),
            .sr(N__47365));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62CED1_19_LC_9_15_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62CED1_19_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62CED1_19_LC_9_15_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62CED1_19_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__26429),
            .in2(_gnd_net_),
            .in3(N__26749),
            .lcout(elapsed_time_ns_1_RNI62CED1_0_19),
            .ltout(elapsed_time_ns_1_RNI62CED1_0_19_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_9_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_9_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_9_15_2 .LUT_INIT=16'b0011001100110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_19_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__27355),
            .in2(N__24254),
            .in3(N__27118),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47804),
            .ce(N__27023),
            .sr(N__47374));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_10_LC_9_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_10_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_10_LC_9_15_3 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_a2_10_LC_9_15_3  (
            .in0(N__27832),
            .in1(N__27426),
            .in2(_gnd_net_),
            .in3(N__27188),
            .lcout(\phase_controller_inst1.stoper_hc.N_315 ),
            .ltout(\phase_controller_inst1.stoper_hc.N_315_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_9_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_9_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_9_15_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_11_LC_9_15_4  (
            .in0(N__31246),
            .in1(N__27356),
            .in2(N__24251),
            .in3(N__27119),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47804),
            .ce(N__27023),
            .sr(N__47374));
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_9_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_9_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_9_15_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_12_LC_9_15_6  (
            .in0(N__24459),
            .in1(N__27357),
            .in2(N__27469),
            .in3(N__27117),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47804),
            .ce(N__27023),
            .sr(N__47374));
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_9_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_9_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_9_15_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_13_LC_9_15_7  (
            .in0(N__27116),
            .in1(N__27358),
            .in2(N__24467),
            .in3(N__27509),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47804),
            .ce(N__27023),
            .sr(N__47374));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILKVDQ_18_LC_9_16_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILKVDQ_18_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILKVDQ_18_LC_9_16_0 .LUT_INIT=16'b1111101011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILKVDQ_18_LC_9_16_0  (
            .in0(N__35927),
            .in1(N__26648),
            .in2(N__31958),
            .in3(N__36974),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI51CED1_18_LC_9_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI51CED1_18_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI51CED1_18_LC_9_16_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI51CED1_18_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24248),
            .in3(N__26752),
            .lcout(elapsed_time_ns_1_RNI51CED1_0_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ4OD11_31_LC_9_16_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ4OD11_31_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ4OD11_31_LC_9_16_3 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ4OD11_31_LC_9_16_3  (
            .in0(N__27251),
            .in1(N__37147),
            .in2(N__36996),
            .in3(N__31791),
            .lcout(elapsed_time_ns_1_RNIQ4OD11_0_31),
            .ltout(elapsed_time_ns_1_RNIQ4OD11_0_31_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_1_9_LC_9_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_1_9_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_1_9_LC_9_16_4 .LUT_INIT=16'b1111001111110010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_i_1_9_LC_9_16_4  (
            .in0(N__27365),
            .in1(N__27105),
            .in2(N__24485),
            .in3(N__26591),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_1Z0Z_9 ),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_1Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_9_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_9_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_9_16_5 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_9_LC_9_16_5  (
            .in0(N__35815),
            .in1(N__27121),
            .in2(N__24473),
            .in3(N__24458),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47800),
            .ce(N__27022),
            .sr(N__47380));
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_9_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_9_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_9_16_6 .LUT_INIT=16'b0000000011111110;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_14_LC_9_16_6  (
            .in0(N__27427),
            .in1(N__27106),
            .in2(N__24468),
            .in3(N__27255),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47800),
            .ce(N__27022),
            .sr(N__47380));
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_9_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_9_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_9_16_7 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_10_LC_9_16_7  (
            .in0(N__27529),
            .in1(N__27120),
            .in2(N__27299),
            .in3(N__24457),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47800),
            .ce(N__27022),
            .sr(N__47380));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_3_LC_9_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_3_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_3_LC_9_17_0 .LUT_INIT=16'b1010101011101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_3_LC_9_17_0  (
            .in0(N__27266),
            .in1(N__24557),
            .in2(N__26576),
            .in3(N__27148),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_0_2_LC_9_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_0_2_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_0_2_LC_9_17_1 .LUT_INIT=16'b0100111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_0_2_LC_9_17_1  (
            .in0(N__26537),
            .in1(N__24555),
            .in2(N__37256),
            .in3(N__26574),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_o2_1_LC_9_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_o2_1_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_o2_1_LC_9_17_2 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_0_o2_1_LC_9_17_2  (
            .in0(_gnd_net_),
            .in1(N__26536),
            .in2(_gnd_net_),
            .in3(N__37252),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.N_283_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_a5_1_LC_9_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_a5_1_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_a5_1_LC_9_17_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_0_a5_1_LC_9_17_3  (
            .in0(N__27147),
            .in1(N__24556),
            .in2(N__24392),
            .in3(N__26575),
            .lcout(\phase_controller_inst1.stoper_hc.N_307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2IMJQ_6_LC_9_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2IMJQ_6_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2IMJQ_6_LC_9_17_4 .LUT_INIT=16'b1111101011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2IMJQ_6_LC_9_17_4  (
            .in0(N__35926),
            .in1(N__24576),
            .in2(N__31871),
            .in3(N__36970),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIU2KD1_6_LC_9_17_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIU2KD1_6_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIU2KD1_6_LC_9_17_5 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIU2KD1_6_LC_9_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24584),
            .in3(N__26751),
            .lcout(elapsed_time_ns_1_RNIIU2KD1_0_6),
            .ltout(elapsed_time_ns_1_RNIIU2KD1_0_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0_2_LC_9_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0_2_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0_2_LC_9_17_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0_2_LC_9_17_6  (
            .in0(N__27376),
            .in1(N__26819),
            .in2(N__24560),
            .in3(N__26847),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2 ),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_6_LC_9_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_6_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_6_LC_9_17_7 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_6_LC_9_17_7  (
            .in0(N__27146),
            .in1(_gnd_net_),
            .in2(N__24542),
            .in3(N__27819),
            .lcout(\phase_controller_inst1.stoper_hc.N_327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0_6_LC_9_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0_6_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0_6_LC_9_18_1 .LUT_INIT=16'b0000101000001110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0_6_LC_9_18_1  (
            .in0(N__27192),
            .in1(N__27383),
            .in2(N__27160),
            .in3(N__27818),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0Z0Z_6 ),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_1_LC_9_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_1_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_1_LC_9_18_2 .LUT_INIT=16'b1111111100110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_1_LC_9_18_2  (
            .in0(_gnd_net_),
            .in1(N__24515),
            .in2(N__24539),
            .in3(N__27300),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITCMJQ_1_LC_9_18_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITCMJQ_1_LC_9_18_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITCMJQ_1_LC_9_18_3 .LUT_INIT=16'b1100111111101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITCMJQ_1_LC_9_18_3  (
            .in0(N__24516),
            .in1(N__35928),
            .in2(N__31574),
            .in3(N__37001),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDP2KD1_1_LC_9_18_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDP2KD1_1_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDP2KD1_1_LC_9_18_4 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDP2KD1_1_LC_9_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24521),
            .in3(N__26756),
            .lcout(elapsed_time_ns_1_RNIDP2KD1_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_9_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_9_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_9_18_6 .LUT_INIT=16'b0000000000110010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_2_LC_9_18_6  (
            .in0(N__24861),
            .in1(N__24496),
            .in2(N__24949),
            .in3(N__27304),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47789),
            .ce(N__27014),
            .sr(N__47393));
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_9_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_9_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_9_18_7 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_4_LC_9_18_7  (
            .in0(N__26698),
            .in1(N__24925),
            .in2(N__27343),
            .in3(N__24862),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47789),
            .ce(N__27014),
            .sr(N__47393));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_1_c_inv_LC_9_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_1_c_inv_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_1_c_inv_LC_9_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_1_c_inv_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__24818),
            .in2(N__24779),
            .in3(N__24806),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_2_c_inv_LC_9_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_2_c_inv_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_2_c_inv_LC_9_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_2_c_inv_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__24770),
            .in2(N__24752),
            .in3(N__24763),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_3_c_inv_LC_9_19_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_3_c_inv_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_3_c_inv_LC_9_19_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_3_c_inv_LC_9_19_2  (
            .in0(N__24742),
            .in1(N__24731),
            .in2(N__24719),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_4_c_inv_LC_9_19_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_4_c_inv_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_4_c_inv_LC_9_19_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_4_c_inv_LC_9_19_3  (
            .in0(N__24710),
            .in1(N__24692),
            .in2(N__24686),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_5_c_inv_LC_9_19_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_5_c_inv_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_5_c_inv_LC_9_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_5_c_inv_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(N__24674),
            .in2(N__24653),
            .in3(N__24664),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_6_c_inv_LC_9_19_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_6_c_inv_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_6_c_inv_LC_9_19_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_6_c_inv_LC_9_19_5  (
            .in0(N__24643),
            .in1(N__24620),
            .in2(N__24632),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_7_c_inv_LC_9_19_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_7_c_inv_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_7_c_inv_LC_9_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_7_c_inv_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(N__24590),
            .in2(N__24614),
            .in3(N__24601),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_8_c_inv_LC_9_19_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_8_c_inv_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_8_c_inv_LC_9_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_8_c_inv_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(N__25145),
            .in2(N__25172),
            .in3(N__25160),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_9_c_inv_LC_9_20_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_9_c_inv_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_9_c_inv_LC_9_20_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_9_c_inv_LC_9_20_0  (
            .in0(_gnd_net_),
            .in1(N__25115),
            .in2(N__25139),
            .in3(N__25126),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_9_20_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_10_c_inv_LC_9_20_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_10_c_inv_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_10_c_inv_LC_9_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_10_c_inv_LC_9_20_1  (
            .in0(_gnd_net_),
            .in1(N__25109),
            .in2(N__25088),
            .in3(N__25099),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_11_c_inv_LC_9_20_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_11_c_inv_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_11_c_inv_LC_9_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_11_c_inv_LC_9_20_2  (
            .in0(_gnd_net_),
            .in1(N__25079),
            .in2(N__25055),
            .in3(N__25066),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_12_c_inv_LC_9_20_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_12_c_inv_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_12_c_inv_LC_9_20_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_12_c_inv_LC_9_20_3  (
            .in0(_gnd_net_),
            .in1(N__25022),
            .in2(N__25046),
            .in3(N__25033),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_13_c_inv_LC_9_20_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_13_c_inv_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_13_c_inv_LC_9_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_13_c_inv_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(N__25016),
            .in2(N__24995),
            .in3(N__25006),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_14_c_inv_LC_9_20_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_14_c_inv_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_14_c_inv_LC_9_20_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_14_c_inv_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(N__24983),
            .in2(N__24962),
            .in3(N__24973),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_15_c_inv_LC_9_20_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_15_c_inv_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_15_c_inv_LC_9_20_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_15_c_inv_LC_9_20_6  (
            .in0(N__25324),
            .in1(N__25313),
            .in2(N__27035),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_16_c_inv_LC_9_20_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_16_c_inv_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_16_c_inv_LC_9_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_16_c_inv_LC_9_20_7  (
            .in0(_gnd_net_),
            .in1(N__25307),
            .in2(N__25286),
            .in3(N__25297),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_17_c_inv_LC_9_21_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_17_c_inv_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_17_c_inv_LC_9_21_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_17_c_inv_LC_9_21_0  (
            .in0(_gnd_net_),
            .in1(N__26462),
            .in2(N__25265),
            .in3(N__25276),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_9_21_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_18_c_inv_LC_9_21_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_18_c_inv_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_18_c_inv_LC_9_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_18_c_inv_LC_9_21_1  (
            .in0(_gnd_net_),
            .in1(N__25256),
            .in2(N__25232),
            .in3(N__25243),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_inv_LC_9_21_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_inv_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_inv_LC_9_21_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_inv_LC_9_21_2  (
            .in0(N__25222),
            .in1(N__25199),
            .in2(N__25211),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_LUT4_0_LC_9_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_LUT4_0_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_LUT4_0_LC_9_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_LUT4_0_LC_9_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25193),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.S1_LC_9_23_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.S1_LC_9_23_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S1_LC_9_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S1_LC_9_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32418),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47767),
            .ce(),
            .sr(N__47418));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIF87U_8_LC_10_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIF87U_8_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIF87U_8_LC_10_8_0 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIF87U_8_LC_10_8_0  (
            .in0(N__25736),
            .in1(N__31090),
            .in2(N__33775),
            .in3(N__28760),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_10_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_10_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_10_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25735),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_10_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_10_8_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_10_8_2 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_10_8_2  (
            .in0(N__28308),
            .in1(N__28158),
            .in2(N__27999),
            .in3(N__25445),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47834),
            .ce(),
            .sr(N__47317));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_10_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_10_8_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_10_8_3 .LUT_INIT=16'b0100111101000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_10_8_3  (
            .in0(N__28156),
            .in1(N__28309),
            .in2(N__25439),
            .in3(N__27974),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47834),
            .ce(),
            .sr(N__47317));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_10_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_10_8_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_10_8_4 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_10_8_4  (
            .in0(N__27967),
            .in1(N__25430),
            .in2(N__28319),
            .in3(N__28159),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47834),
            .ce(),
            .sr(N__47317));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI428M_12_LC_10_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI428M_12_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI428M_12_LC_10_8_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI428M_12_LC_10_8_5  (
            .in0(N__25548),
            .in1(N__40519),
            .in2(N__28479),
            .in3(N__28306),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_10_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_10_8_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_10_8_6 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_10_8_6  (
            .in0(N__28307),
            .in1(N__28157),
            .in2(N__27998),
            .in3(N__25412),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47834),
            .ce(),
            .sr(N__47317));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI318M_30_LC_10_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI318M_30_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI318M_30_LC_10_8_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI318M_30_LC_10_8_7  (
            .in0(N__25547),
            .in1(N__40520),
            .in2(N__28478),
            .in3(N__40605),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIB36U_7_LC_10_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIB36U_7_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIB36U_7_LC_10_9_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIB36U_7_LC_10_9_0  (
            .in0(N__25697),
            .in1(N__33695),
            .in2(N__30830),
            .in3(N__28769),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6I_LC_10_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6I_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6I_LC_10_9_1 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6I_LC_10_9_1  (
            .in0(N__25382),
            .in1(N__30644),
            .in2(N__33757),
            .in3(N__28859),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_10_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_10_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_10_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26298),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_10_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_10_9_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_10_9_3  (
            .in0(N__33692),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28636),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIVJ2U_4_LC_10_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIVJ2U_4_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIVJ2U_4_LC_10_9_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIVJ2U_4_LC_10_9_4  (
            .in0(N__25616),
            .in1(N__33693),
            .in2(N__30923),
            .in3(N__28538),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKP_LC_10_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKP_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKP_LC_10_9_5 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKP_LC_10_9_5  (
            .in0(N__30767),
            .in1(N__28696),
            .in2(N__33756),
            .in3(N__28679),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI7U4U_6_LC_10_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI7U4U_6_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI7U4U_6_LC_10_9_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI7U4U_6_LC_10_9_6  (
            .in0(N__26165),
            .in1(N__33694),
            .in2(N__30868),
            .in3(N__28514),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84I_LC_10_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84I_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84I_LC_10_10_0 .LUT_INIT=16'b0101101011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84I_LC_10_10_0  (
            .in0(N__28937),
            .in1(N__25558),
            .in2(N__28913),
            .in3(N__33712),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22I_LC_10_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22I_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22I_LC_10_10_1 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22I_LC_10_10_1  (
            .in0(N__28483),
            .in1(N__28991),
            .in2(N__33759),
            .in3(N__29015),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_10_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_10_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_10_10_2  (
            .in0(N__29036),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33703),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ),
            .ltout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0I_LC_10_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0I_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0I_LC_10_10_3 .LUT_INIT=16'b0101111111110101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0I_LC_10_10_3  (
            .in0(N__33708),
            .in1(N__25505),
            .in2(N__25469),
            .in3(N__29024),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVH_LC_10_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVH_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVH_LC_10_10_4 .LUT_INIT=16'b0101101011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVH_LC_10_10_4  (
            .in0(N__28635),
            .in1(N__26013),
            .in2(N__28616),
            .in3(N__33707),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53I_LC_10_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53I_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53I_LC_10_10_5 .LUT_INIT=16'b0011110011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53I_LC_10_10_5  (
            .in0(N__40536),
            .in1(N__28979),
            .in2(N__28952),
            .in3(N__33741),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_inv_LC_10_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_inv_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_inv_LC_10_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_inv_LC_10_10_6  (
            .in0(_gnd_net_),
            .in1(N__28697),
            .in2(_gnd_net_),
            .in3(N__33702),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MP_LC_10_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MP_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MP_LC_10_10_7 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MP_LC_10_10_7  (
            .in0(N__25952),
            .in1(N__28663),
            .in2(N__33758),
            .in3(N__28646),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31J_LC_10_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31J_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31J_LC_10_11_0 .LUT_INIT=16'b0011111111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31J_LC_10_11_0  (
            .in0(N__25906),
            .in1(N__33718),
            .in2(N__28808),
            .in3(N__28778),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_inv_LC_10_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_inv_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_inv_LC_10_11_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_inv_LC_10_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33760),
            .in3(N__28667),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00J_LC_10_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00J_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00J_LC_10_11_2 .LUT_INIT=16'b0011111111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00J_LC_10_11_2  (
            .in0(N__25856),
            .in1(N__33717),
            .in2(N__28847),
            .in3(N__28817),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45J_LC_10_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45J_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45J_LC_10_11_3 .LUT_INIT=16'b0101111110101111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45J_LC_10_11_3  (
            .in0(N__31361),
            .in1(N__30698),
            .in2(N__33761),
            .in3(N__29132),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_10_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_10_11_4 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_10_11_4  (
            .in0(N__25796),
            .in1(N__25746),
            .in2(N__25715),
            .in3(N__25664),
            .lcout(\current_shift_inst.PI_CTRL.N_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_10_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_10_11_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_10_11_5  (
            .in0(N__33716),
            .in1(N__29165),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ),
            .ltout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62J_LC_10_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62J_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62J_LC_10_11_6 .LUT_INIT=16'b0101111111110101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62J_LC_10_11_6  (
            .in0(N__33755),
            .in1(N__27598),
            .in2(N__26249),
            .in3(N__29153),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14J_LC_10_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14J_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14J_LC_10_11_7 .LUT_INIT=16'b0110111101101111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14J_LC_10_11_7  (
            .in0(N__31289),
            .in1(N__29144),
            .in2(N__33762),
            .in3(N__26236),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_10_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_10_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_10_12_0  (
            .in0(N__28933),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33669),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_10_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_10_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_10_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26175),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_10_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_10_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_10_12_2  (
            .in0(N__29057),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33670),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ),
            .ltout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJ_LC_10_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJ_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJ_LC_10_12_3 .LUT_INIT=16'b0101111111110101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJ_LC_10_12_3  (
            .in0(N__33676),
            .in1(N__26125),
            .in2(N__26081),
            .in3(N__29045),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76J_LC_10_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76J_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76J_LC_10_12_4 .LUT_INIT=16'b0101101011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76J_LC_10_12_4  (
            .in0(N__31313),
            .in1(N__26071),
            .in2(N__29120),
            .in3(N__33671),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP2ND11_21_LC_10_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP2ND11_21_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP2ND11_21_LC_10_12_5 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP2ND11_21_LC_10_12_5  (
            .in0(N__26506),
            .in1(N__37154),
            .in2(N__31703),
            .in3(N__36981),
            .lcout(elapsed_time_ns_1_RNIP2ND11_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7J_LC_10_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7J_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7J_LC_10_12_6 .LUT_INIT=16'b0101101011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7J_LC_10_12_6  (
            .in0(N__29106),
            .in1(N__26366),
            .in2(N__29087),
            .in3(N__33672),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8J_LC_10_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8J_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8J_LC_10_12_7 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8J_LC_10_12_7  (
            .in0(N__30499),
            .in1(N__31388),
            .in2(N__33745),
            .in3(N__29075),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIURK5B_31_LC_10_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIURK5B_31_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIURK5B_31_LC_10_13_0 .LUT_INIT=16'b0101010101000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIURK5B_31_LC_10_13_0  (
            .in0(N__31793),
            .in1(N__31526),
            .in2(N__31844),
            .in3(N__31817),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc5 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHGVDQ_14_LC_10_13_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHGVDQ_14_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHGVDQ_14_LC_10_13_1 .LUT_INIT=16'b1111101011111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHGVDQ_14_LC_10_13_1  (
            .in0(N__31898),
            .in1(N__27404),
            .in2(N__26306),
            .in3(N__36897),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1TBED1_14_LC_10_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1TBED1_14_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1TBED1_14_LC_10_13_2 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1TBED1_14_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26303),
            .in3(N__26735),
            .lcout(elapsed_time_ns_1_RNI1TBED1_0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV8ND11_27_LC_10_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV8ND11_27_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV8ND11_27_LC_10_13_3 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV8ND11_27_LC_10_13_3  (
            .in0(N__37102),
            .in1(N__26393),
            .in2(N__29402),
            .in3(N__36895),
            .lcout(elapsed_time_ns_1_RNIV8ND11_0_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9J_LC_10_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9J_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9J_LC_10_13_4 .LUT_INIT=16'b0111101101111011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9J_LC_10_13_4  (
            .in0(N__29066),
            .in1(N__33744),
            .in2(N__31337),
            .in3(N__26299),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU7ND11_26_LC_10_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU7ND11_26_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU7ND11_26_LC_10_13_5 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU7ND11_26_LC_10_13_5  (
            .in0(N__37103),
            .in1(N__26378),
            .in2(N__29426),
            .in3(N__36896),
            .lcout(elapsed_time_ns_1_RNIU7ND11_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL13KD1_9_LC_10_13_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL13KD1_9_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL13KD1_9_LC_10_13_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL13KD1_9_LC_10_13_6  (
            .in0(_gnd_net_),
            .in1(N__26734),
            .in2(_gnd_net_),
            .in3(N__35780),
            .lcout(elapsed_time_ns_1_RNIL13KD1_0_9),
            .ltout(elapsed_time_ns_1_RNIL13KD1_0_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_9_LC_10_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_9_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_9_LC_10_13_7 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_9_LC_10_13_7  (
            .in0(_gnd_net_),
            .in1(N__27831),
            .in2(N__26423),
            .in3(N__27403),
            .lcout(\phase_controller_inst1.stoper_hc.N_328 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1BND11_29_LC_10_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1BND11_29_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1BND11_29_LC_10_14_0 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1BND11_29_LC_10_14_0  (
            .in0(N__37075),
            .in1(N__26420),
            .in2(N__29348),
            .in3(N__36864),
            .lcout(elapsed_time_ns_1_RNI1BND11_0_29),
            .ltout(elapsed_time_ns_1_RNI1BND11_0_29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0_15_LC_10_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0_15_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0_15_LC_10_14_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0_15_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26414),
            .in3(N__29212),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGCC0J_31_LC_10_14_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGCC0J_31_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGCC0J_31_LC_10_14_2 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGCC0J_31_LC_10_14_2  (
            .in0(N__47479),
            .in1(N__29171),
            .in2(N__31792),
            .in3(N__29195),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ2MD11_13_LC_10_14_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ2MD11_13_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ2MD11_13_LC_10_14_3 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ2MD11_13_LC_10_14_3  (
            .in0(N__36867),
            .in1(N__37078),
            .in2(N__31445),
            .in3(N__27503),
            .lcout(elapsed_time_ns_1_RNIQ2MD11_0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0AND11_28_LC_10_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0AND11_28_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0AND11_28_LC_10_14_4 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0AND11_28_LC_10_14_4  (
            .in0(N__37077),
            .in1(N__26402),
            .in2(N__29375),
            .in3(N__36866),
            .lcout(elapsed_time_ns_1_RNI0AND11_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS5ND11_24_LC_10_14_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS5ND11_24_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS5ND11_24_LC_10_14_5 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS5ND11_24_LC_10_14_5  (
            .in0(N__36868),
            .in1(N__26492),
            .in2(N__37153),
            .in3(N__29468),
            .lcout(elapsed_time_ns_1_RNIS5ND11_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIT6ND11_25_LC_10_14_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIT6ND11_25_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIT6ND11_25_LC_10_14_6 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIT6ND11_25_LC_10_14_6  (
            .in0(N__37076),
            .in1(N__36865),
            .in2(N__26411),
            .in3(N__29450),
            .lcout(elapsed_time_ns_1_RNIT6ND11_0_25),
            .ltout(elapsed_time_ns_1_RNIT6ND11_0_25_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6_15_LC_10_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6_15_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6_15_LC_10_14_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6_15_LC_10_14_7  (
            .in0(N__26401),
            .in1(N__26392),
            .in2(N__26381),
            .in3(N__26377),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7_15_LC_10_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7_15_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7_15_LC_10_15_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7_15_LC_10_15_0  (
            .in0(N__26437),
            .in1(N__26449),
            .in2(N__26510),
            .in3(N__26491),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_15_LC_10_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_15_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_15_LC_10_15_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_o5_15_LC_10_15_1  (
            .in0(N__26480),
            .in1(N__36815),
            .in2(N__26474),
            .in3(N__26471),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_10_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_10_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_10_15_2 .LUT_INIT=16'b0011001100110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_17_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(N__27298),
            .in2(N__26465),
            .in3(N__26673),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47795),
            .ce(N__27013),
            .sr(N__47358));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ3ND11_22_LC_10_15_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ3ND11_22_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ3ND11_22_LC_10_15_3 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ3ND11_22_LC_10_15_3  (
            .in0(N__26450),
            .in1(N__37106),
            .in2(N__31721),
            .in3(N__36898),
            .lcout(elapsed_time_ns_1_RNIQ3ND11_0_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKJVDQ_17_LC_10_15_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKJVDQ_17_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKJVDQ_17_LC_10_15_5 .LUT_INIT=16'b1111111011110010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKJVDQ_17_LC_10_15_5  (
            .in0(N__26674),
            .in1(N__36899),
            .in2(N__35922),
            .in3(N__31973),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI40CED1_17_LC_10_15_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI40CED1_17_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI40CED1_17_LC_10_15_6 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI40CED1_17_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26441),
            .in3(N__26748),
            .lcout(elapsed_time_ns_1_RNI40CED1_0_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIR4ND11_23_LC_10_15_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIR4ND11_23_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIR4ND11_23_LC_10_15_7 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIR4ND11_23_LC_10_15_7  (
            .in0(N__37105),
            .in1(N__26438),
            .in2(N__36994),
            .in3(N__29486),
            .lcout(elapsed_time_ns_1_RNIR4ND11_0_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMLVDQ_19_LC_10_16_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMLVDQ_19_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMLVDQ_19_LC_10_16_0 .LUT_INIT=16'b1111111010111010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMLVDQ_19_LC_10_16_0  (
            .in0(N__35918),
            .in1(N__36969),
            .in2(N__26618),
            .in3(N__31926),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQURR91_3_LC_10_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQURR91_3_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQURR91_3_LC_10_16_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQURR91_3_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(N__35917),
            .in2(_gnd_net_),
            .in3(N__26516),
            .lcout(elapsed_time_ns_1_RNIQURR91_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992_24_LC_10_16_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992_24_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992_24_LC_10_16_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992_24_LC_10_16_2  (
            .in0(N__26561),
            .in1(N__27545),
            .in2(N__29446),
            .in3(N__29464),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3VBED1_16_LC_10_16_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3VBED1_16_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3VBED1_16_LC_10_16_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3VBED1_16_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(N__33878),
            .in2(_gnd_net_),
            .in3(N__26750),
            .lcout(elapsed_time_ns_1_RNI3VBED1_0_16),
            .ltout(elapsed_time_ns_1_RNI3VBED1_0_16_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_9_LC_10_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_9_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_9_LC_10_16_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_9_LC_10_16_4  (
            .in0(N__26671),
            .in1(N__26638),
            .in2(N__26705),
            .in3(N__26612),
            .lcout(\phase_controller_inst1.stoper_hc.N_278 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA3DJ11_4_LC_10_16_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA3DJ11_4_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA3DJ11_4_LC_10_16_5 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA3DJ11_4_LC_10_16_5  (
            .in0(N__37146),
            .in1(N__31592),
            .in2(N__36995),
            .in3(N__26691),
            .lcout(elapsed_time_ns_1_RNIA3DJ11_0_4),
            .ltout(elapsed_time_ns_1_RNIA3DJ11_0_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3_2_LC_10_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3_2_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3_2_LC_10_16_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3_2_LC_10_16_6  (
            .in0(N__26672),
            .in1(N__26787),
            .in2(N__26651),
            .in3(N__33929),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_2_LC_10_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_2_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_2_LC_10_16_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_2_LC_10_16_7  (
            .in0(N__26639),
            .in1(N__26613),
            .in2(N__26594),
            .in3(N__26590),
            .lcout(\phase_controller_inst1.stoper_hc.N_337 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9PDO_26_LC_10_17_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9PDO_26_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9PDO_26_LC_10_17_0 .LUT_INIT=16'b1111111011111110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9PDO_26_LC_10_17_0  (
            .in0(N__29416),
            .in1(N__29389),
            .in2(N__29368),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP1MD11_12_LC_10_17_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP1MD11_12_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP1MD11_12_LC_10_17_1 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP1MD11_12_LC_10_17_1  (
            .in0(N__36961),
            .in1(N__37145),
            .in2(N__31499),
            .in3(N__27448),
            .lcout(elapsed_time_ns_1_RNIP1MD11_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS27MU_3_LC_10_17_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS27MU_3_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS27MU_3_LC_10_17_2 .LUT_INIT=16'b1110111011111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS27MU_3_LC_10_17_2  (
            .in0(N__31547),
            .in1(N__31985),
            .in2(N__26555),
            .in3(N__36962),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTI01_20_LC_10_17_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTI01_20_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTI01_20_LC_10_17_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTI01_20_LC_10_17_3  (
            .in0(N__29338),
            .in1(N__29482),
            .in2(N__37018),
            .in3(N__29653),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVLD11_10_LC_10_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVLD11_10_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVLD11_10_LC_10_17_4 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVLD11_10_LC_10_17_4  (
            .in0(N__27525),
            .in1(N__31484),
            .in2(N__36982),
            .in3(N__37144),
            .lcout(elapsed_time_ns_1_RNINVLD11_0_10),
            .ltout(elapsed_time_ns_1_RNINVLD11_0_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2_2_LC_10_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2_2_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2_2_LC_10_17_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2_2_LC_10_17_5  (
            .in0(N__31245),
            .in1(N__27504),
            .in2(N__27473),
            .in3(N__27447),
            .lcout(\phase_controller_inst1.stoper_hc.N_319 ),
            .ltout(\phase_controller_inst1.stoper_hc.N_319_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0_6_LC_10_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0_6_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0_6_LC_10_17_6 .LUT_INIT=16'b0101000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0_6_LC_10_17_6  (
            .in0(N__35820),
            .in1(_gnd_net_),
            .in2(N__27434),
            .in3(N__27416),
            .lcout(\phase_controller_inst1.stoper_hc.N_275 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a5_1_0_9_LC_10_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a5_1_0_9_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a5_1_0_9_LC_10_17_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a5_1_0_9_LC_10_17_7  (
            .in0(N__27817),
            .in1(N__35821),
            .in2(_gnd_net_),
            .in3(N__27377),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_a5_1_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_10_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_10_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_10_18_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_15_LC_10_18_0  (
            .in0(N__27820),
            .in1(N__27305),
            .in2(N__27197),
            .in3(N__27142),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47781),
            .ce(N__27016),
            .sr(N__47381));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNID6DJ11_7_LC_10_18_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNID6DJ11_7_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNID6DJ11_7_LC_10_18_1 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNID6DJ11_7_LC_10_18_1  (
            .in0(N__37143),
            .in1(N__31166),
            .in2(N__37000),
            .in3(N__26853),
            .lcout(elapsed_time_ns_1_RNID6DJ11_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE7DJ11_8_LC_10_18_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE7DJ11_8_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE7DJ11_8_LC_10_18_3 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE7DJ11_8_LC_10_18_3  (
            .in0(N__37142),
            .in1(N__31187),
            .in2(N__36999),
            .in3(N__26826),
            .lcout(elapsed_time_ns_1_RNIE7DJ11_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB4DJ11_5_LC_10_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB4DJ11_5_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB4DJ11_5_LC_10_18_5 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB4DJ11_5_LC_10_18_5  (
            .in0(N__37141),
            .in1(N__36984),
            .in2(N__31613),
            .in3(N__26786),
            .lcout(elapsed_time_ns_1_RNIB4DJ11_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS4MD11_15_LC_10_18_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS4MD11_15_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS4MD11_15_LC_10_18_7 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS4MD11_15_LC_10_18_7  (
            .in0(N__31211),
            .in1(N__27821),
            .in2(N__37155),
            .in3(N__36983),
            .lcout(elapsed_time_ns_1_RNIS4MD11_0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNI8HMG_LC_10_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNI8HMG_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNI8HMG_LC_10_19_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNI8HMG_LC_10_19_0  (
            .in0(N__27706),
            .in1(N__27751),
            .in2(_gnd_net_),
            .in3(N__27781),
            .lcout(\phase_controller_inst2.stoper_hc.running_1_sqmuxa ),
            .ltout(\phase_controller_inst2.stoper_hc.running_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_10_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_10_19_1 .LUT_INIT=16'b0000111100000111;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_10_19_1  (
            .in0(N__27752),
            .in1(N__27707),
            .in2(N__27674),
            .in3(N__27671),
            .lcout(\phase_controller_inst2.stoper_hc.un1_start_latched2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.S2_LC_10_24_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.S2_LC_10_24_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S2_LC_10_24_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S2_LC_10_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34043),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47761),
            .ce(),
            .sr(N__47417));
    defparam SB_DFF_inst_PH1_MAX_D2_LC_11_5_5.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_11_5_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_11_5_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D2_LC_11_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27629),
            .lcout(il_max_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47854),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D1_LC_11_6_0.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_11_6_0.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_11_6_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH2_MIN_D1_LC_11_6_0 (
            .in0(N__27620),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_min_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47843),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D2_LC_11_6_6.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_11_6_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_11_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MIN_D2_LC_11_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27605),
            .lcout(il_min_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47843),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_11_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_11_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(N__28800),
            .in2(_gnd_net_),
            .in3(N__33763),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_11_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_11_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27595),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_11_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_11_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28465),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI5R941_10_LC_11_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI5R941_10_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI5R941_10_LC_11_8_4 .LUT_INIT=16'b1111000000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI5R941_10_LC_11_8_4  (
            .in0(N__28427),
            .in1(N__31024),
            .in2(N__28727),
            .in3(N__33765),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI3P3U_5_LC_11_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI3P3U_5_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI3P3U_5_LC_11_8_7 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI3P3U_5_LC_11_8_7  (
            .in0(N__33764),
            .in1(N__30558),
            .in2(N__28529),
            .in3(N__30892),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_11_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_11_9_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_11_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_0_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36161),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47822),
            .ce(),
            .sr(N__47318));
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_11_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_11_9_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_11_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_0_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28574),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47822),
            .ce(),
            .sr(N__47318));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_11_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_11_9_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_11_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30829),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47822),
            .ce(),
            .sr(N__47318));
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_11_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_11_9_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_11_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_1_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30983),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47822),
            .ce(),
            .sr(N__47318));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_11_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_11_9_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_11_9_5 .LUT_INIT=16'b0101000111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_11_9_5  (
            .in0(N__28328),
            .in1(N__28318),
            .in2(N__28166),
            .in3(N__27997),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47822),
            .ce(),
            .sr(N__47318));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_11_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_11_9_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_11_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30922),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47822),
            .ce(),
            .sr(N__47318));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_11_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_11_9_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_11_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30893),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47822),
            .ce(),
            .sr(N__47318));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_11_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_11_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__28562),
            .in2(_gnd_net_),
            .in3(N__28573),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_11_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_11_10_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_11_10_1  (
            .in0(N__30979),
            .in1(N__28556),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_11_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_11_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(N__28550),
            .in2(_gnd_net_),
            .in3(N__30961),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_11_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_11_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__28544),
            .in2(_gnd_net_),
            .in3(N__30937),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_11_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_11_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(N__30995),
            .in2(_gnd_net_),
            .in3(N__28532),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_11_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_11_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(N__30716),
            .in2(_gnd_net_),
            .in3(N__28517),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_11_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_11_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(N__30704),
            .in2(_gnd_net_),
            .in3(N__28508),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_11_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_11_10_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(N__30788),
            .in2(_gnd_net_),
            .in3(N__28763),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_11_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_11_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__31067),
            .in2(_gnd_net_),
            .in3(N__28745),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_8 ),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_11_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_11_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(N__31034),
            .in2(_gnd_net_),
            .in3(N__28730),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_11_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_11_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(N__31001),
            .in2(_gnd_net_),
            .in3(N__28715),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_11_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_11_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(N__30710),
            .in2(_gnd_net_),
            .in3(N__28700),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_LUT4_0_LC_11_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_LUT4_0_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_LUT4_0_LC_11_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_LUT4_0_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(N__28695),
            .in2(_gnd_net_),
            .in3(N__28670),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_LUT4_0_LC_11_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_LUT4_0_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_LUT4_0_LC_11_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_LUT4_0_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(N__28662),
            .in2(_gnd_net_),
            .in3(N__28640),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_11_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_11_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_11_11_6  (
            .in0(_gnd_net_),
            .in1(N__28637),
            .in2(_gnd_net_),
            .in3(N__28607),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_11_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_11_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(N__29035),
            .in2(_gnd_net_),
            .in3(N__29018),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_11_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_11_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(N__29014),
            .in2(_gnd_net_),
            .in3(N__28982),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_11_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_11_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_11_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(N__28975),
            .in2(_gnd_net_),
            .in3(N__28940),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_11_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_11_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(N__28929),
            .in2(_gnd_net_),
            .in3(N__28901),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_11_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_11_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(N__28898),
            .in2(_gnd_net_),
            .in3(N__28862),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_11_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_11_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(N__30640),
            .in2(_gnd_net_),
            .in3(N__28850),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_11_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_11_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(N__28840),
            .in2(_gnd_net_),
            .in3(N__28811),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_11_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_11_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(N__28801),
            .in2(_gnd_net_),
            .in3(N__28772),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_11_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_11_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_11_12_7  (
            .in0(_gnd_net_),
            .in1(N__29164),
            .in2(_gnd_net_),
            .in3(N__29147),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_11_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_11_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__31281),
            .in2(_gnd_net_),
            .in3(N__29135),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO ),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_11_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_11_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(N__31353),
            .in2(_gnd_net_),
            .in3(N__29123),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_11_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_11_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(N__31305),
            .in2(_gnd_net_),
            .in3(N__29111),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_11_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_11_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(N__29107),
            .in2(_gnd_net_),
            .in3(N__29078),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_11_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_11_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31384),
            .in3(N__29069),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_11_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_11_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(N__31329),
            .in2(_gnd_net_),
            .in3(N__29060),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_11_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_11_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(N__29056),
            .in2(_gnd_net_),
            .in3(N__29039),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54K_LC_11_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54K_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54K_LC_11_13_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54K_LC_11_13_7  (
            .in0(N__29273),
            .in1(N__33602),
            .in2(_gnd_net_),
            .in3(N__29234),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5I_31_LC_11_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5I_31_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5I_31_LC_11_14_0 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5I_31_LC_11_14_0  (
            .in0(N__32003),
            .in1(N__47476),
            .in2(N__31622),
            .in3(N__31505),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK670F_31_LC_11_14_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK670F_31_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK670F_31_LC_11_14_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK670F_31_LC_11_14_1  (
            .in0(N__32002),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31732),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_382_i ),
            .ltout(\delay_measurement_inst.delay_hc_timer.N_382_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP3OD11_30_LC_11_14_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP3OD11_30_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP3OD11_30_LC_11_14_2 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP3OD11_30_LC_11_14_2  (
            .in0(N__29213),
            .in1(N__29660),
            .in2(N__29216),
            .in3(N__37131),
            .lcout(elapsed_time_ns_1_RNIP3OD11_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91_7_LC_11_14_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91_7_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91_7_LC_11_14_3 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91_7_LC_11_14_3  (
            .in0(N__35845),
            .in1(N__31183),
            .in2(_gnd_net_),
            .in3(N__31162),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2_15_LC_11_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2_15_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2_15_LC_11_14_4 .LUT_INIT=16'b1110111011101100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2_15_LC_11_14_4  (
            .in0(N__31894),
            .in1(N__31210),
            .in2(N__29201),
            .in3(N__31423),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6_15_LC_11_14_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6_15_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6_15_LC_11_14_5 .LUT_INIT=16'b1111111110110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6_15_LC_11_14_5  (
            .in0(N__31904),
            .in1(N__31681),
            .in2(N__29198),
            .in3(N__29188),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719_21_LC_11_14_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719_21_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719_21_LC_11_14_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719_21_LC_11_14_6  (
            .in0(N__31682),
            .in1(N__47475),
            .in2(N__29189),
            .in3(N__32001),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9_24_LC_11_14_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9_24_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9_24_LC_11_14_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9_24_LC_11_14_7  (
            .in0(N__31519),
            .in1(N__29184),
            .in2(_gnd_net_),
            .in3(N__31403),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_11_15_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_11_15_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_11_15_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__29636),
            .in2(N__29608),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__47790),
            .ce(N__37177),
            .sr(N__47349));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_11_15_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_11_15_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_11_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__37225),
            .in2(N__29576),
            .in3(N__29297),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__47790),
            .ce(N__37177),
            .sr(N__47349));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_11_15_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_11_15_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_11_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(N__29609),
            .in2(N__29545),
            .in3(N__29294),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__47790),
            .ce(N__37177),
            .sr(N__47349));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_11_15_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_11_15_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_11_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__29575),
            .in2(N__29518),
            .in3(N__29291),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc5lto6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__47790),
            .ce(N__37177),
            .sr(N__47349));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_11_15_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_11_15_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_11_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__29884),
            .in2(N__29546),
            .in3(N__29288),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__47790),
            .ce(N__37177),
            .sr(N__47349));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_11_15_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_11_15_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_11_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(N__29857),
            .in2(N__29519),
            .in3(N__29285),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__47790),
            .ce(N__37177),
            .sr(N__47349));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_11_15_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_11_15_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_11_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(N__29827),
            .in2(N__29888),
            .in3(N__29282),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc5lto9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__47790),
            .ce(N__37177),
            .sr(N__47349));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_11_15_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_11_15_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_11_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(N__29858),
            .in2(N__29800),
            .in3(N__29279),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__47790),
            .ce(N__37177),
            .sr(N__47349));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_11_16_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_11_16_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_11_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_11_16_0  (
            .in0(_gnd_net_),
            .in1(N__29767),
            .in2(N__29834),
            .in3(N__29276),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_11_16_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__47785),
            .ce(N__37176),
            .sr(N__47359));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_11_16_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_11_16_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_11_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(N__29801),
            .in2(N__29743),
            .in3(N__29324),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__47785),
            .ce(N__37176),
            .sr(N__47359));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_11_16_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_11_16_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_11_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(N__29768),
            .in2(N__29716),
            .in3(N__29321),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__47785),
            .ce(N__37176),
            .sr(N__47359));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_11_16_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_11_16_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_11_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_11_16_3  (
            .in0(_gnd_net_),
            .in1(N__29686),
            .in2(N__29744),
            .in3(N__29318),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc5lto14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__47785),
            .ce(N__37176),
            .sr(N__47359));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_11_16_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_11_16_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_11_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(N__30106),
            .in2(N__29717),
            .in3(N__29315),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc5lto15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__47785),
            .ce(N__37176),
            .sr(N__47359));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_11_16_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_11_16_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_11_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(N__30079),
            .in2(N__29690),
            .in3(N__29312),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__47785),
            .ce(N__37176),
            .sr(N__47359));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_11_16_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_11_16_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_11_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__30052),
            .in2(N__30110),
            .in3(N__29309),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__47785),
            .ce(N__37176),
            .sr(N__47359));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_11_16_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_11_16_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_11_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_11_16_7  (
            .in0(_gnd_net_),
            .in1(N__30080),
            .in2(N__30022),
            .in3(N__29306),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__47785),
            .ce(N__37176),
            .sr(N__47359));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_11_17_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_11_17_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_11_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_11_17_0  (
            .in0(_gnd_net_),
            .in1(N__29986),
            .in2(N__30056),
            .in3(N__29303),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__47782),
            .ce(N__37175),
            .sr(N__47366));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_11_17_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_11_17_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_11_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(N__29959),
            .in2(N__30023),
            .in3(N__29300),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__47782),
            .ce(N__37175),
            .sr(N__47366));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_11_17_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_11_17_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_11_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(N__29938),
            .in2(N__29990),
            .in3(N__29492),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__47782),
            .ce(N__37175),
            .sr(N__47366));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_11_17_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_11_17_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_11_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(N__29960),
            .in2(N__29918),
            .in3(N__29489),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__47782),
            .ce(N__37175),
            .sr(N__47366));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_11_17_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_11_17_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_11_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(N__29939),
            .in2(N__30436),
            .in3(N__29471),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__47782),
            .ce(N__37175),
            .sr(N__47366));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_11_17_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_11_17_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_11_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(N__29917),
            .in2(N__30409),
            .in3(N__29453),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__47782),
            .ce(N__37175),
            .sr(N__47366));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_11_17_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_11_17_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_11_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(N__30379),
            .in2(N__30437),
            .in3(N__29429),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__47782),
            .ce(N__37175),
            .sr(N__47366));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_11_17_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_11_17_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_11_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(N__30355),
            .in2(N__30410),
            .in3(N__29405),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__47782),
            .ce(N__37175),
            .sr(N__47366));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_11_18_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_11_18_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_11_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(N__30325),
            .in2(N__30383),
            .in3(N__29378),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__47777),
            .ce(N__37174),
            .sr(N__47375));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_11_18_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_11_18_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_11_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(N__30356),
            .in2(N__30298),
            .in3(N__29351),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__47777),
            .ce(N__37174),
            .sr(N__47375));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_11_18_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_11_18_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_11_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(N__30272),
            .in2(N__30329),
            .in3(N__29327),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__47777),
            .ce(N__37174),
            .sr(N__47375));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_11_18_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_11_18_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_11_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(N__30251),
            .in2(N__30299),
            .in3(N__29642),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__47777),
            .ce(N__37174),
            .sr(N__47375));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_11_18_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_11_18_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_11_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29639),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47777),
            .ce(N__37174),
            .sr(N__47375));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_11_18_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_11_18_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_11_18_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_11_18_7  (
            .in0(_gnd_net_),
            .in1(N__29635),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47777),
            .ce(N__37174),
            .sr(N__47375));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_11_19_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_11_19_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_11_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_11_19_0  (
            .in0(N__30233),
            .in1(N__29631),
            .in2(_gnd_net_),
            .in3(N__29615),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_11_19_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__47772),
            .ce(N__32312),
            .sr(N__47382));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_11_19_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_11_19_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_11_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_11_19_1  (
            .in0(N__30229),
            .in1(N__37218),
            .in2(_gnd_net_),
            .in3(N__29612),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__47772),
            .ce(N__32312),
            .sr(N__47382));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_11_19_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_11_19_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_11_19_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_11_19_2  (
            .in0(N__30234),
            .in1(N__29601),
            .in2(_gnd_net_),
            .in3(N__29579),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__47772),
            .ce(N__32312),
            .sr(N__47382));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_11_19_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_11_19_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_11_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_11_19_3  (
            .in0(N__30230),
            .in1(N__29565),
            .in2(_gnd_net_),
            .in3(N__29549),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__47772),
            .ce(N__32312),
            .sr(N__47382));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_11_19_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_11_19_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_11_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_11_19_4  (
            .in0(N__30235),
            .in1(N__29538),
            .in2(_gnd_net_),
            .in3(N__29522),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__47772),
            .ce(N__32312),
            .sr(N__47382));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_11_19_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_11_19_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_11_19_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_11_19_5  (
            .in0(N__30231),
            .in1(N__29506),
            .in2(_gnd_net_),
            .in3(N__29891),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__47772),
            .ce(N__32312),
            .sr(N__47382));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_11_19_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_11_19_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_11_19_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_11_19_6  (
            .in0(N__30236),
            .in1(N__29877),
            .in2(_gnd_net_),
            .in3(N__29861),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__47772),
            .ce(N__32312),
            .sr(N__47382));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_11_19_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_11_19_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_11_19_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_11_19_7  (
            .in0(N__30232),
            .in1(N__29851),
            .in2(_gnd_net_),
            .in3(N__29837),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__47772),
            .ce(N__32312),
            .sr(N__47382));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_11_20_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_11_20_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_11_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_11_20_0  (
            .in0(N__30220),
            .in1(N__29826),
            .in2(_gnd_net_),
            .in3(N__29804),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_11_20_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__47769),
            .ce(N__32307),
            .sr(N__47388));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_11_20_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_11_20_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_11_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_11_20_1  (
            .in0(N__30224),
            .in1(N__29793),
            .in2(_gnd_net_),
            .in3(N__29771),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__47769),
            .ce(N__32307),
            .sr(N__47388));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_11_20_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_11_20_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_11_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_11_20_2  (
            .in0(N__30217),
            .in1(N__29761),
            .in2(_gnd_net_),
            .in3(N__29747),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__47769),
            .ce(N__32307),
            .sr(N__47388));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_11_20_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_11_20_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_11_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_11_20_3  (
            .in0(N__30221),
            .in1(N__29736),
            .in2(_gnd_net_),
            .in3(N__29720),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__47769),
            .ce(N__32307),
            .sr(N__47388));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_11_20_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_11_20_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_11_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_11_20_4  (
            .in0(N__30218),
            .in1(N__29709),
            .in2(_gnd_net_),
            .in3(N__29693),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__47769),
            .ce(N__32307),
            .sr(N__47388));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_11_20_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_11_20_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_11_20_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_11_20_5  (
            .in0(N__30222),
            .in1(N__29679),
            .in2(_gnd_net_),
            .in3(N__29663),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__47769),
            .ce(N__32307),
            .sr(N__47388));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_11_20_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_11_20_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_11_20_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_11_20_6  (
            .in0(N__30219),
            .in1(N__30099),
            .in2(_gnd_net_),
            .in3(N__30083),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__47769),
            .ce(N__32307),
            .sr(N__47388));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_11_20_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_11_20_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_11_20_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_11_20_7  (
            .in0(N__30223),
            .in1(N__30073),
            .in2(_gnd_net_),
            .in3(N__30059),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__47769),
            .ce(N__32307),
            .sr(N__47388));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_11_21_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_11_21_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_11_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_11_21_0  (
            .in0(N__30213),
            .in1(N__30045),
            .in2(_gnd_net_),
            .in3(N__30026),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_11_21_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__47764),
            .ce(N__32311),
            .sr(N__47394));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_11_21_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_11_21_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_11_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_11_21_1  (
            .in0(N__30225),
            .in1(N__30009),
            .in2(_gnd_net_),
            .in3(N__29993),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__47764),
            .ce(N__32311),
            .sr(N__47394));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_11_21_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_11_21_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_11_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_11_21_2  (
            .in0(N__30214),
            .in1(N__29979),
            .in2(_gnd_net_),
            .in3(N__29963),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__47764),
            .ce(N__32311),
            .sr(N__47394));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_11_21_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_11_21_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_11_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_11_21_3  (
            .in0(N__30226),
            .in1(N__29958),
            .in2(_gnd_net_),
            .in3(N__29942),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__47764),
            .ce(N__32311),
            .sr(N__47394));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_11_21_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_11_21_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_11_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_11_21_4  (
            .in0(N__30215),
            .in1(N__29937),
            .in2(_gnd_net_),
            .in3(N__29921),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__47764),
            .ce(N__32311),
            .sr(N__47394));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_11_21_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_11_21_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_11_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_11_21_5  (
            .in0(N__30227),
            .in1(N__29913),
            .in2(_gnd_net_),
            .in3(N__29894),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__47764),
            .ce(N__32311),
            .sr(N__47394));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_11_21_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_11_21_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_11_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_11_21_6  (
            .in0(N__30216),
            .in1(N__30429),
            .in2(_gnd_net_),
            .in3(N__30413),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__47764),
            .ce(N__32311),
            .sr(N__47394));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_11_21_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_11_21_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_11_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_11_21_7  (
            .in0(N__30228),
            .in1(N__30402),
            .in2(_gnd_net_),
            .in3(N__30386),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__47764),
            .ce(N__32311),
            .sr(N__47394));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_11_22_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_11_22_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_11_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_11_22_0  (
            .in0(N__30189),
            .in1(N__30378),
            .in2(_gnd_net_),
            .in3(N__30359),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_11_22_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__47762),
            .ce(N__32294),
            .sr(N__47399));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_11_22_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_11_22_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_11_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_11_22_1  (
            .in0(N__30193),
            .in1(N__30348),
            .in2(_gnd_net_),
            .in3(N__30332),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__47762),
            .ce(N__32294),
            .sr(N__47399));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_11_22_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_11_22_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_11_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_11_22_2  (
            .in0(N__30190),
            .in1(N__30318),
            .in2(_gnd_net_),
            .in3(N__30302),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__47762),
            .ce(N__32294),
            .sr(N__47399));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_11_22_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_11_22_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_11_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_11_22_3  (
            .in0(N__30194),
            .in1(N__30291),
            .in2(_gnd_net_),
            .in3(N__30275),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__47762),
            .ce(N__32294),
            .sr(N__47399));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_11_22_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_11_22_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_11_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_11_22_4  (
            .in0(N__30191),
            .in1(N__30271),
            .in2(_gnd_net_),
            .in3(N__30257),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__47762),
            .ce(N__32294),
            .sr(N__47399));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_11_22_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_11_22_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_11_22_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_11_22_5  (
            .in0(N__30250),
            .in1(N__30192),
            .in2(_gnd_net_),
            .in3(N__30254),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47762),
            .ce(N__32294),
            .sr(N__47399));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_11_23_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_11_23_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_11_23_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_11_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32217),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_11_24_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_11_24_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_11_24_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_11_24_7  (
            .in0(_gnd_net_),
            .in1(N__32216),
            .in2(_gnd_net_),
            .in3(N__32246),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_432_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D2_LC_12_4_1.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_12_4_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_12_4_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D2_LC_12_4_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30587),
            .lcout(il_min_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47853),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D1_LC_12_4_3.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_12_4_3.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_12_4_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D1_LC_12_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30599),
            .lcout(il_min_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47853),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_hc_LC_12_6_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_12_6_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_hc_LC_12_6_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_12_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32267),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30580),
            .ce(),
            .sr(N__47299));
    defparam \delay_measurement_inst.stop_timer_hc_LC_12_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_12_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_hc_LC_12_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_12_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32268),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30581),
            .ce(),
            .sr(N__47304));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_12_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_12_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_12_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30557),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_0_12_LC_12_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_0_12_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_0_12_LC_12_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_0_12_LC_12_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33766),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_i_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_12_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_12_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_12_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30495),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_12_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_12_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_12_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33376),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_12_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_12_9_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_12_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_2_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30965),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47817),
            .ce(),
            .sr(N__47314));
    defparam \phase_controller_inst1.stoper_tr.running_LC_12_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_LC_12_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.running_LC_12_9_7 .LUT_INIT=16'b1010101000101110;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_LC_12_9_7  (
            .in0(N__42900),
            .in1(N__42845),
            .in2(N__42980),
            .in3(N__43043),
            .lcout(\phase_controller_inst1.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47817),
            .ce(),
            .sr(N__47314));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_12_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_12_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30814),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_12_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_12_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30746),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30885),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31119),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30849),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_12_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_12_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30696),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_12_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_12_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_12_10_6  (
            .in0(N__30639),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33679),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_12_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_12_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30907),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(N__30989),
            .in2(_gnd_net_),
            .in3(N__36157),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ),
            .ltout(),
            .carryin(bfn_12_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_12_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_12_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_12_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_1_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(N__35942),
            .in2(_gnd_net_),
            .in3(N__30968),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .clk(N__47805),
            .ce(),
            .sr(N__47323));
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_12_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_12_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_12_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_LC_12_11_2  (
            .in0(_gnd_net_),
            .in1(N__31265),
            .in2(_gnd_net_),
            .in3(N__30950),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .clk(N__47805),
            .ce(),
            .sr(N__47323));
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_12_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_12_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_12_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_3_LC_12_11_3  (
            .in0(_gnd_net_),
            .in1(N__31397),
            .in2(_gnd_net_),
            .in3(N__30926),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .clk(N__47805),
            .ce(),
            .sr(N__47323));
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_12_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_12_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_12_11_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_4_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33956),
            .in3(N__30896),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .clk(N__47805),
            .ce(),
            .sr(N__47323));
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_12_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_12_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_12_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_5_LC_12_11_5  (
            .in0(_gnd_net_),
            .in1(N__34523),
            .in2(_gnd_net_),
            .in3(N__30872),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .clk(N__47805),
            .ce(),
            .sr(N__47323));
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_12_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_12_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_12_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_6_LC_12_11_6  (
            .in0(_gnd_net_),
            .in1(N__33788),
            .in2(_gnd_net_),
            .in3(N__30833),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .clk(N__47805),
            .ce(),
            .sr(N__47323));
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_12_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_12_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_12_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_7_LC_12_11_7  (
            .in0(_gnd_net_),
            .in1(N__34571),
            .in2(_gnd_net_),
            .in3(N__31145),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .clk(N__47805),
            .ce(),
            .sr(N__47323));
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_12_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_12_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_12_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_8_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__33293),
            .in2(_gnd_net_),
            .in3(N__31142),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_8 ),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .clk(N__47801),
            .ce(),
            .sr(N__47328));
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_12_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_12_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_12_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_9_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__33476),
            .in2(_gnd_net_),
            .in3(N__31139),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .clk(N__47801),
            .ce(),
            .sr(N__47328));
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_12_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_12_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_12_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_10_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__32324),
            .in2(_gnd_net_),
            .in3(N__31136),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .clk(N__47801),
            .ce(),
            .sr(N__47328));
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_12_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_12_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_12_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_11_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(N__33863),
            .in2(_gnd_net_),
            .in3(N__31100),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .clk(N__47801),
            .ce(),
            .sr(N__47328));
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_12_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_12_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_12_12_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_12_LC_12_12_4  (
            .in0(_gnd_net_),
            .in1(N__36671),
            .in2(_gnd_net_),
            .in3(N__31097),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47801),
            .ce(),
            .sr(N__47328));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_12_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_12_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31078),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_12_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_12_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_12_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31045),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31012),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36512),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_12_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_12_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_12_13_2  (
            .in0(N__31383),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33600),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_12_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_12_13_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_12_13_3  (
            .in0(N__33598),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31357),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_12_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_12_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_12_13_4  (
            .in0(N__31333),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33601),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_12_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_12_13_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_12_13_5  (
            .in0(N__33599),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31309),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_12_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_12_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_12_13_6  (
            .in0(N__31285),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33597),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36125),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO0MD11_11_LC_12_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO0MD11_11_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO0MD11_11_LC_12_14_0 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO0MD11_11_LC_12_14_0  (
            .in0(N__31235),
            .in1(N__36934),
            .in2(N__31469),
            .in3(N__37104),
            .lcout(elapsed_time_ns_1_RNIO0MD11_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542_15_LC_12_14_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542_15_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542_15_LC_12_14_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542_15_LC_12_14_1  (
            .in0(N__31209),
            .in1(N__31182),
            .in2(N__31427),
            .in3(N__31161),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU4A94_9_LC_12_14_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU4A94_9_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU4A94_9_LC_12_14_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU4A94_9_LC_12_14_2  (
            .in0(N__35844),
            .in1(N__31580),
            .in2(N__31631),
            .in3(N__31628),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKR_2_LC_12_14_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKR_2_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKR_2_LC_12_14_3 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKR_2_LC_12_14_3  (
            .in0(N__31539),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37201),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKRZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847_31_LC_12_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847_31_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847_31_LC_12_14_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847_31_LC_12_14_4  (
            .in0(N__47474),
            .in1(N__31786),
            .in2(_gnd_net_),
            .in3(N__31813),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_12_14_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_12_14_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(N__31603),
            .in2(_gnd_net_),
            .in3(N__31591),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352_1_LC_12_14_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352_1_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352_1_LC_12_14_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352_1_LC_12_14_6  (
            .in0(N__37202),
            .in1(N__31573),
            .in2(N__31550),
            .in3(N__31540),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4_31_LC_12_14_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4_31_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4_31_LC_12_14_7 .LUT_INIT=16'b1101110000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4_31_LC_12_14_7  (
            .in0(N__31787),
            .in1(N__47473),
            .in2(N__31508),
            .in3(N__31837),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_12_15_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_12_15_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_12_15_0  (
            .in0(N__31495),
            .in1(N__31480),
            .in2(N__31462),
            .in3(N__31438),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3PJ05_15_LC_12_15_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3PJ05_15_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3PJ05_15_LC_12_15_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3PJ05_15_LC_12_15_1  (
            .in0(N__47477),
            .in1(N__31833),
            .in2(N__31675),
            .in3(N__31409),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_a3_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJV461_16_LC_12_15_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJV461_16_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJV461_16_LC_12_15_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJV461_16_LC_12_15_2  (
            .in0(N__31887),
            .in1(N__31861),
            .in2(N__33898),
            .in3(N__31951),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_17_LC_12_15_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_17_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_17_LC_12_15_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_17_LC_12_15_3  (
            .in0(N__31972),
            .in1(N__31934),
            .in2(N__32012),
            .in3(N__32009),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58F_31_LC_12_15_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58F_31_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58F_31_LC_12_15_4 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58F_31_LC_12_15_4  (
            .in0(N__31733),
            .in1(_gnd_net_),
            .in2(N__31988),
            .in3(N__47478),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58FZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_12_15_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_12_15_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_12_15_5  (
            .in0(N__31971),
            .in1(N__31950),
            .in2(N__31933),
            .in3(N__33891),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642_6_LC_12_15_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642_6_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642_6_LC_12_15_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642_6_LC_12_15_6  (
            .in0(N__31886),
            .in1(N__31860),
            .in2(N__31847),
            .in3(N__35843),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09_31_LC_12_15_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09_31_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09_31_LC_12_15_7 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09_31_LC_12_15_7  (
            .in0(N__31812),
            .in1(_gnd_net_),
            .in2(N__31796),
            .in3(N__31771),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_12_16_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_12_16_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__31714),
            .in2(_gnd_net_),
            .in3(N__31693),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_12_16_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_12_16_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_12_16_2 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_12_16_2  (
            .in0(N__33847),
            .in1(N__33360),
            .in2(_gnd_net_),
            .in3(N__33821),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47780),
            .ce(),
            .sr(N__47350));
    defparam \phase_controller_inst2.T01_LC_12_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.T01_LC_12_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.T01_LC_12_16_5 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \phase_controller_inst2.T01_LC_12_16_5  (
            .in0(N__31642),
            .in1(N__32398),
            .in2(_gnd_net_),
            .in3(N__32148),
            .lcout(T01_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47780),
            .ce(),
            .sr(N__47350));
    defparam \phase_controller_inst2.T12_LC_12_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.T12_LC_12_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.T12_LC_12_16_7 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \phase_controller_inst2.T12_LC_12_16_7  (
            .in0(N__32167),
            .in1(N__34029),
            .in2(_gnd_net_),
            .in3(N__32149),
            .lcout(T12_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47780),
            .ce(),
            .sr(N__47350));
    defparam \phase_controller_inst2.state_1_LC_12_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_1_LC_12_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_1_LC_12_17_2 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \phase_controller_inst2.state_1_LC_12_17_2  (
            .in0(N__33996),
            .in1(N__32156),
            .in2(N__32123),
            .in3(N__34027),
            .lcout(\phase_controller_inst2.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47776),
            .ce(),
            .sr(N__47360));
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_12_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_12_17_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(N__34696),
            .in2(_gnd_net_),
            .in3(N__34656),
            .lcout(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_0_LC_12_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_0_LC_12_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_0_LC_12_17_4 .LUT_INIT=16'b1100000011101010;
    LogicCell40 \phase_controller_inst2.state_0_LC_12_17_4  (
            .in0(N__32362),
            .in1(N__34028),
            .in2(N__34001),
            .in3(N__34769),
            .lcout(\phase_controller_inst2.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47776),
            .ce(),
            .sr(N__47360));
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNI9M3O_LC_12_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNI9M3O_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNI9M3O_LC_12_17_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_RNI9M3O_LC_12_17_5  (
            .in0(_gnd_net_),
            .in1(N__34768),
            .in2(_gnd_net_),
            .in3(N__32361),
            .lcout(\phase_controller_inst2.time_passed_RNI9M3O ),
            .ltout(\phase_controller_inst2.time_passed_RNI9M3O_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_3_LC_12_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_3_LC_12_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_3_LC_12_17_6 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \phase_controller_inst2.state_3_LC_12_17_6  (
            .in0(N__32399),
            .in1(N__32084),
            .in2(N__32048),
            .in3(N__37585),
            .lcout(\phase_controller_inst2.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47776),
            .ce(),
            .sr(N__47360));
    defparam \phase_controller_inst2.start_timer_tr_LC_12_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_LC_12_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_tr_LC_12_18_1 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \phase_controller_inst2.start_timer_tr_LC_12_18_1  (
            .in0(N__34812),
            .in1(N__32045),
            .in2(N__34677),
            .in3(N__33962),
            .lcout(\phase_controller_inst2.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47771),
            .ce(),
            .sr(N__47367));
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_12_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_12_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_12_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_LC_12_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34660),
            .lcout(\phase_controller_inst2.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47771),
            .ce(),
            .sr(N__47367));
    defparam \phase_controller_inst2.T23_LC_12_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.T23_LC_12_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.T23_LC_12_19_0 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \phase_controller_inst2.T23_LC_12_19_0  (
            .in0(N__32023),
            .in1(N__34036),
            .in2(_gnd_net_),
            .in3(N__32368),
            .lcout(T23_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47768),
            .ce(),
            .sr(N__47376));
    defparam \phase_controller_inst2.T45_LC_12_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.T45_LC_12_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.T45_LC_12_19_2 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \phase_controller_inst2.T45_LC_12_19_2  (
            .in0(N__32408),
            .in1(N__32335),
            .in2(_gnd_net_),
            .in3(N__32369),
            .lcout(T45_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47768),
            .ce(),
            .sr(N__47376));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_12_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_12_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_12_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36407),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_4_LC_12_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_12_20_2 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_12_20_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.state_4_LC_12_20_2  (
            .in0(_gnd_net_),
            .in1(N__34147),
            .in2(_gnd_net_),
            .in3(N__34802),
            .lcout(phase_controller_inst1_state_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47763),
            .ce(),
            .sr(N__47383));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_12_23_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_12_23_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_12_23_3 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_12_23_3  (
            .in0(N__32218),
            .in1(N__32275),
            .in2(_gnd_net_),
            .in3(N__32244),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_433_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_12_24_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_12_24_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_12_24_1 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_12_24_1  (
            .in0(N__32219),
            .in1(N__32276),
            .in2(_gnd_net_),
            .in3(N__32245),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47758),
            .ce(),
            .sr(N__47405));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_13_5_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_13_5_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_13_5_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_13_5_0  (
            .in0(N__32600),
            .in1(N__34059),
            .in2(_gnd_net_),
            .in3(N__32195),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_13_5_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__47855),
            .ce(N__33335),
            .sr(N__47285));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_13_5_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_13_5_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_13_5_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_13_5_1  (
            .in0(N__32596),
            .in1(N__34338),
            .in2(_gnd_net_),
            .in3(N__32192),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__47855),
            .ce(N__33335),
            .sr(N__47285));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_13_5_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_13_5_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_13_5_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_13_5_2  (
            .in0(N__32601),
            .in1(N__32835),
            .in2(_gnd_net_),
            .in3(N__32189),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__47855),
            .ce(N__33335),
            .sr(N__47285));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_13_5_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_13_5_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_13_5_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_13_5_3  (
            .in0(N__32597),
            .in1(N__32809),
            .in2(_gnd_net_),
            .in3(N__32186),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__47855),
            .ce(N__33335),
            .sr(N__47285));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_13_5_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_13_5_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_13_5_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_13_5_4  (
            .in0(N__32602),
            .in1(N__32784),
            .in2(_gnd_net_),
            .in3(N__32447),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__47855),
            .ce(N__33335),
            .sr(N__47285));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_13_5_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_13_5_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_13_5_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_13_5_5  (
            .in0(N__32598),
            .in1(N__32760),
            .in2(_gnd_net_),
            .in3(N__32444),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__47855),
            .ce(N__33335),
            .sr(N__47285));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_13_5_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_13_5_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_13_5_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_13_5_6  (
            .in0(N__32603),
            .in1(N__32731),
            .in2(_gnd_net_),
            .in3(N__32441),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__47855),
            .ce(N__33335),
            .sr(N__47285));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_13_5_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_13_5_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_13_5_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_13_5_7  (
            .in0(N__32599),
            .in1(N__32701),
            .in2(_gnd_net_),
            .in3(N__32438),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__47855),
            .ce(N__33335),
            .sr(N__47285));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_13_6_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_13_6_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_13_6_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_13_6_0  (
            .in0(N__32591),
            .in1(N__32673),
            .in2(_gnd_net_),
            .in3(N__32435),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_13_6_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__47844),
            .ce(N__33338),
            .sr(N__47293));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_13_6_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_13_6_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_13_6_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_13_6_1  (
            .in0(N__32595),
            .in1(N__32643),
            .in2(_gnd_net_),
            .in3(N__32432),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__47844),
            .ce(N__33338),
            .sr(N__47293));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_13_6_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_13_6_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_13_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_13_6_2  (
            .in0(N__32588),
            .in1(N__33061),
            .in2(_gnd_net_),
            .in3(N__32429),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__47844),
            .ce(N__33338),
            .sr(N__47293));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_13_6_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_13_6_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_13_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_13_6_3  (
            .in0(N__32592),
            .in1(N__33037),
            .in2(_gnd_net_),
            .in3(N__32426),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__47844),
            .ce(N__33338),
            .sr(N__47293));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_13_6_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_13_6_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_13_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_13_6_4  (
            .in0(N__32589),
            .in1(N__33012),
            .in2(_gnd_net_),
            .in3(N__32423),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__47844),
            .ce(N__33338),
            .sr(N__47293));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_13_6_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_13_6_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_13_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_13_6_5  (
            .in0(N__32593),
            .in1(N__32985),
            .in2(_gnd_net_),
            .in3(N__32474),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__47844),
            .ce(N__33338),
            .sr(N__47293));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_13_6_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_13_6_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_13_6_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_13_6_6  (
            .in0(N__32590),
            .in1(N__32959),
            .in2(_gnd_net_),
            .in3(N__32471),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__47844),
            .ce(N__33338),
            .sr(N__47293));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_13_6_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_13_6_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_13_6_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_13_6_7  (
            .in0(N__32594),
            .in1(N__32931),
            .in2(_gnd_net_),
            .in3(N__32468),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__47844),
            .ce(N__33338),
            .sr(N__47293));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_13_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_13_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_13_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_13_7_0  (
            .in0(N__32560),
            .in1(N__32901),
            .in2(_gnd_net_),
            .in3(N__32465),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_13_7_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__47835),
            .ce(N__33337),
            .sr(N__47300));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_13_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_13_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_13_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_13_7_1  (
            .in0(N__32564),
            .in1(N__32871),
            .in2(_gnd_net_),
            .in3(N__32462),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__47835),
            .ce(N__33337),
            .sr(N__47300));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_13_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_13_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_13_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_13_7_2  (
            .in0(N__32561),
            .in1(N__33279),
            .in2(_gnd_net_),
            .in3(N__32459),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__47835),
            .ce(N__33337),
            .sr(N__47300));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_13_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_13_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_13_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_13_7_3  (
            .in0(N__32565),
            .in1(N__33258),
            .in2(_gnd_net_),
            .in3(N__32456),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__47835),
            .ce(N__33337),
            .sr(N__47300));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_13_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_13_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_13_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_13_7_4  (
            .in0(N__32562),
            .in1(N__33231),
            .in2(_gnd_net_),
            .in3(N__32453),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__47835),
            .ce(N__33337),
            .sr(N__47300));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_13_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_13_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_13_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_13_7_5  (
            .in0(N__32566),
            .in1(N__33204),
            .in2(_gnd_net_),
            .in3(N__32450),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__47835),
            .ce(N__33337),
            .sr(N__47300));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_13_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_13_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_13_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_13_7_6  (
            .in0(N__32563),
            .in1(N__33178),
            .in2(_gnd_net_),
            .in3(N__32624),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__47835),
            .ce(N__33337),
            .sr(N__47300));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_13_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_13_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_13_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_13_7_7  (
            .in0(N__32567),
            .in1(N__33150),
            .in2(_gnd_net_),
            .in3(N__32621),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__47835),
            .ce(N__33337),
            .sr(N__47300));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_13_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_13_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_13_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_13_8_0  (
            .in0(N__32556),
            .in1(N__33117),
            .in2(_gnd_net_),
            .in3(N__32618),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_13_8_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__47828),
            .ce(N__33336),
            .sr(N__47305));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_13_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_13_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_13_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_13_8_1  (
            .in0(N__32568),
            .in1(N__33093),
            .in2(_gnd_net_),
            .in3(N__32615),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__47828),
            .ce(N__33336),
            .sr(N__47305));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_13_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_13_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_13_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_13_8_2  (
            .in0(N__32557),
            .in1(N__33462),
            .in2(_gnd_net_),
            .in3(N__32612),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__47828),
            .ce(N__33336),
            .sr(N__47305));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_13_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_13_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_13_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_13_8_3  (
            .in0(N__32569),
            .in1(N__33399),
            .in2(_gnd_net_),
            .in3(N__32609),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__47828),
            .ce(N__33336),
            .sr(N__47305));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_13_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_13_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_13_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_13_8_4  (
            .in0(N__32558),
            .in1(N__33442),
            .in2(_gnd_net_),
            .in3(N__32606),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__47828),
            .ce(N__33336),
            .sr(N__47305));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_13_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_13_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_13_8_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_13_8_5  (
            .in0(N__33424),
            .in1(N__32559),
            .in2(_gnd_net_),
            .in3(N__32477),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47828),
            .ce(N__33336),
            .sr(N__47305));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_13_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_13_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_13_9_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_13_9_0  (
            .in0(_gnd_net_),
            .in1(N__34064),
            .in2(N__32846),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_13_9_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__47823),
            .ce(N__34300),
            .sr(N__47311));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_13_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_13_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_13_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_13_9_1  (
            .in0(_gnd_net_),
            .in1(N__32815),
            .in2(N__34352),
            .in3(N__32849),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__47823),
            .ce(N__34300),
            .sr(N__47311));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_13_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_13_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_13_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_13_9_2  (
            .in0(_gnd_net_),
            .in1(N__32845),
            .in2(N__32791),
            .in3(N__32819),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__47823),
            .ce(N__34300),
            .sr(N__47311));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_13_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_13_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_13_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_13_9_3  (
            .in0(_gnd_net_),
            .in1(N__32816),
            .in2(N__32765),
            .in3(N__32795),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__47823),
            .ce(N__34300),
            .sr(N__47311));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_13_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_13_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_13_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_13_9_4  (
            .in0(_gnd_net_),
            .in1(N__32737),
            .in2(N__32792),
            .in3(N__32768),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__47823),
            .ce(N__34300),
            .sr(N__47311));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_13_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_13_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_13_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_13_9_5  (
            .in0(_gnd_net_),
            .in1(N__32764),
            .in2(N__32713),
            .in3(N__32741),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__47823),
            .ce(N__34300),
            .sr(N__47311));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_13_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_13_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_13_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_13_9_6  (
            .in0(_gnd_net_),
            .in1(N__32738),
            .in2(N__32680),
            .in3(N__32717),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__47823),
            .ce(N__34300),
            .sr(N__47311));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_13_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_13_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_13_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_13_9_7  (
            .in0(_gnd_net_),
            .in1(N__32644),
            .in2(N__32714),
            .in3(N__32687),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__47823),
            .ce(N__34300),
            .sr(N__47311));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_13_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_13_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_13_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(N__33067),
            .in2(N__32684),
            .in3(N__32654),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_13_10_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__47818),
            .ce(N__34302),
            .sr(N__47315));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_13_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_13_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_13_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_13_10_1  (
            .in0(_gnd_net_),
            .in1(N__33043),
            .in2(N__32651),
            .in3(N__33071),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__47818),
            .ce(N__34302),
            .sr(N__47315));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_13_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_13_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_13_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_13_10_2  (
            .in0(_gnd_net_),
            .in1(N__33068),
            .in2(N__33019),
            .in3(N__33047),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__47818),
            .ce(N__34302),
            .sr(N__47315));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_13_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_13_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_13_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_13_10_3  (
            .in0(_gnd_net_),
            .in1(N__33044),
            .in2(N__32992),
            .in3(N__33023),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__47818),
            .ce(N__34302),
            .sr(N__47315));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_13_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_13_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_13_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_13_10_4  (
            .in0(_gnd_net_),
            .in1(N__32965),
            .in2(N__33020),
            .in3(N__32996),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__47818),
            .ce(N__34302),
            .sr(N__47315));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_13_10_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_13_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_13_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_13_10_5  (
            .in0(_gnd_net_),
            .in1(N__32938),
            .in2(N__32993),
            .in3(N__32969),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__47818),
            .ce(N__34302),
            .sr(N__47315));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_13_10_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_13_10_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_13_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_13_10_6  (
            .in0(_gnd_net_),
            .in1(N__32966),
            .in2(N__32908),
            .in3(N__32945),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__47818),
            .ce(N__34302),
            .sr(N__47315));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_13_10_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_13_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_13_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_13_10_7  (
            .in0(_gnd_net_),
            .in1(N__32872),
            .in2(N__32942),
            .in3(N__32915),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__47818),
            .ce(N__34302),
            .sr(N__47315));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_13_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_13_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_13_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(N__33280),
            .in2(N__32912),
            .in3(N__32882),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_13_11_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__47812),
            .ce(N__34303),
            .sr(N__47319));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_13_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_13_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_13_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_13_11_1  (
            .in0(_gnd_net_),
            .in1(N__33259),
            .in2(N__32879),
            .in3(N__32852),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__47812),
            .ce(N__34303),
            .sr(N__47319));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_13_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_13_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_13_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_13_11_2  (
            .in0(_gnd_net_),
            .in1(N__33281),
            .in2(N__33238),
            .in3(N__33263),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__47812),
            .ce(N__34303),
            .sr(N__47319));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_13_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_13_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_13_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_13_11_3  (
            .in0(_gnd_net_),
            .in1(N__33260),
            .in2(N__33211),
            .in3(N__33242),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__47812),
            .ce(N__34303),
            .sr(N__47319));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_13_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_13_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_13_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_13_11_4  (
            .in0(_gnd_net_),
            .in1(N__33184),
            .in2(N__33239),
            .in3(N__33215),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__47812),
            .ce(N__34303),
            .sr(N__47319));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_13_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_13_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_13_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_13_11_5  (
            .in0(_gnd_net_),
            .in1(N__33157),
            .in2(N__33212),
            .in3(N__33188),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__47812),
            .ce(N__34303),
            .sr(N__47319));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_13_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_13_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_13_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_13_11_6  (
            .in0(_gnd_net_),
            .in1(N__33185),
            .in2(N__33130),
            .in3(N__33164),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__47812),
            .ce(N__34303),
            .sr(N__47319));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_13_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_13_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_13_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_13_11_7  (
            .in0(_gnd_net_),
            .in1(N__33094),
            .in2(N__33161),
            .in3(N__33134),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__47812),
            .ce(N__34303),
            .sr(N__47319));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_13_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_13_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_13_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_13_12_0  (
            .in0(_gnd_net_),
            .in1(N__33463),
            .in2(N__33131),
            .in3(N__33101),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_13_12_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__47806),
            .ce(N__34304),
            .sr(N__47324));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_13_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_13_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_13_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__33406),
            .in2(N__33098),
            .in3(N__33074),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__47806),
            .ce(N__34304),
            .sr(N__47324));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_13_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_13_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_13_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(N__33464),
            .in2(N__33446),
            .in3(N__33428),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__47806),
            .ce(N__34304),
            .sr(N__47324));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_13_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_13_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_13_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(N__33425),
            .in2(N__33410),
            .in3(N__33383),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__47806),
            .ce(N__34304),
            .sr(N__47324));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_13_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_13_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_13_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33380),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47806),
            .ce(N__34304),
            .sr(N__47324));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_13_13_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_13_13_1 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_13_13_1  (
            .in0(N__33366),
            .in1(N__33840),
            .in2(_gnd_net_),
            .in3(N__33815),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_435_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_13_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_13_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36437),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_13_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_13_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_13_13_4 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_13_13_4  (
            .in0(N__34719),
            .in1(N__34734),
            .in2(_gnd_net_),
            .in3(N__34678),
            .lcout(\phase_controller_inst2.stoper_tr.un2_start_0 ),
            .ltout(\phase_controller_inst2.stoper_tr.un2_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNI2FGQ1_LC_13_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNI2FGQ1_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNI2FGQ1_LC_13_13_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNI2FGQ1_LC_13_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33287),
            .in3(N__34612),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNI2FGQZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNIP8O21_0_LC_13_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNIP8O21_0_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNIP8O21_0_LC_13_13_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNIP8O21_0_LC_13_13_6  (
            .in0(N__34720),
            .in1(N__34679),
            .in2(_gnd_net_),
            .in3(N__35546),
            .lcout(\phase_controller_inst2.stoper_tr.running_1_sqmuxa ),
            .ltout(\phase_controller_inst2.stoper_tr.running_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_13_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_13_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_13_13_7 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_13_13_7  (
            .in0(N__34735),
            .in1(N__34680),
            .in2(N__33284),
            .in3(N__34721),
            .lcout(\phase_controller_inst2.stoper_tr.un1_start_latched2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_tr_LC_13_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_13_14_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_tr_LC_13_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_13_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33820),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33797),
            .ce(),
            .sr(N__47331));
    defparam \delay_measurement_inst.start_timer_tr_LC_13_14_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_13_14_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_tr_LC_13_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_13_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33819),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33797),
            .ce(),
            .sr(N__47331));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_13_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_13_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_13_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36467),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_13_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_13_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_13_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33691),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_i_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_13_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_13_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_13_15_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_13_15_7  (
            .in0(N__44586),
            .in1(N__48084),
            .in2(N__45070),
            .in3(N__41111),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_13_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_13_16_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_13_16_0  (
            .in0(N__44626),
            .in1(N__45237),
            .in2(N__45488),
            .in3(N__43882),
            .lcout(\current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_13_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_13_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36422),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_13_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_13_16_2 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_13_16_2  (
            .in0(N__44628),
            .in1(N__45234),
            .in2(N__46361),
            .in3(N__43613),
            .lcout(\current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_13_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_13_16_3 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_13_16_3  (
            .in0(N__45233),
            .in1(N__44627),
            .in2(N__41216),
            .in3(N__46424),
            .lcout(\current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_13_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_13_16_4 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_13_16_4  (
            .in0(N__44625),
            .in1(N__45236),
            .in2(N__45917),
            .in3(N__40774),
            .lcout(\current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_13_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_13_16_5 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_13_16_5  (
            .in0(N__45235),
            .in1(N__44629),
            .in2(N__46241),
            .in3(N__43552),
            .lcout(\current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_13_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_13_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_inv_LC_13_16_6  (
            .in0(N__38798),
            .in1(N__38557),
            .in2(_gnd_net_),
            .in3(N__34091),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_31 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_13_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_13_16_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_13_16_7  (
            .in0(N__40637),
            .in1(_gnd_net_),
            .in2(N__33866),
            .in3(N__38799),
            .lcout(\current_shift_inst.un38_control_input_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_13_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_13_17_0 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_13_17_0  (
            .in0(N__46873),
            .in1(N__44622),
            .in2(N__41002),
            .in3(N__45241),
            .lcout(\current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_13_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_13_17_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_13_17_1  (
            .in0(N__44623),
            .in1(N__48242),
            .in2(N__45278),
            .in3(N__45323),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_13_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_13_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36664),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_13_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_13_17_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_13_17_5  (
            .in0(N__44025),
            .in1(N__46872),
            .in2(_gnd_net_),
            .in3(N__40995),
            .lcout(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_13_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_13_17_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_13_17_6  (
            .in0(N__44014),
            .in1(N__46234),
            .in2(_gnd_net_),
            .in3(N__43553),
            .lcout(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_13_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_13_17_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_13_17_7  (
            .in0(N__44621),
            .in1(N__45915),
            .in2(N__45279),
            .in3(N__40778),
            .lcout(\current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_13_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_13_18_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_13_18_0  (
            .in0(N__44624),
            .in1(N__46874),
            .in2(N__45280),
            .in3(N__41003),
            .lcout(\current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_13_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_13_18_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_13_18_2  (
            .in0(N__43996),
            .in1(N__46946),
            .in2(_gnd_net_),
            .in3(N__41156),
            .lcout(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_13_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_13_18_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.start_timer_tr_RNO_0_LC_13_18_5  (
            .in0(N__34026),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34000),
            .lcout(\phase_controller_inst2.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_13_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_13_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_13_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36497),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJIVDQ_16_LC_13_18_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJIVDQ_16_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJIVDQ_16_LC_13_18_7 .LUT_INIT=16'b1111111011011100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJIVDQ_16_LC_13_18_7  (
            .in0(N__36980),
            .in1(N__35930),
            .in2(N__33941),
            .in3(N__33902),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_13_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_13_19_0 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_13_19_0  (
            .in0(N__44657),
            .in1(N__48002),
            .in2(N__41288),
            .in3(N__45147),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_RNO_1_11_LC_13_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_RNO_1_11_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_RNO_1_11_LC_13_19_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.control_input_RNO_1_11_LC_13_19_3  (
            .in0(N__45146),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44658),
            .lcout(\current_shift_inst.un38_control_input_axb_31_s0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_13_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_13_19_4 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_13_19_4  (
            .in0(N__44655),
            .in1(N__46750),
            .in2(N__40970),
            .in3(N__45148),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_13_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_13_19_5 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_13_19_5  (
            .in0(N__46751),
            .in1(N__40969),
            .in2(N__45232),
            .in3(N__44656),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_13_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_13_19_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_13_19_6  (
            .in0(N__43997),
            .in1(N__46749),
            .in2(_gnd_net_),
            .in3(N__40965),
            .lcout(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_13_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_13_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_13_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_13_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47021),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47773),
            .ce(N__47509),
            .sr(N__47368));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_13_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_13_20_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_13_20_0  (
            .in0(N__44659),
            .in1(N__48167),
            .in2(N__45293),
            .in3(N__44201),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_13_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_13_20_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_13_20_2  (
            .in0(N__44660),
            .in1(N__48001),
            .in2(N__45292),
            .in3(N__41284),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_13_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_13_20_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_13_20_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.state_ns_i_a3_1_LC_13_20_7  (
            .in0(_gnd_net_),
            .in1(N__34146),
            .in2(_gnd_net_),
            .in3(N__34801),
            .lcout(state_ns_i_a3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_13_23_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_13_23_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_13_23_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_13_23_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_24_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_24_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_24_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47020),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47760),
            .ce(N__47508),
            .sr(N__47400));
    defparam \phase_controller_inst1.S2_LC_13_25_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_13_25_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_13_25_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_13_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38438),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47759),
            .ce(),
            .sr(N__47406));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_14_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_14_6_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_14_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_14_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34063),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47856),
            .ce(N__34299),
            .sr(N__47286));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI56UV7_1_LC_14_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI56UV7_1_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI56UV7_1_LC_14_7_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI56UV7_1_LC_14_7_0  (
            .in0(N__34404),
            .in1(N__34474),
            .in2(N__34448),
            .in3(N__34181),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_359_1 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_359_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILL1NA_6_LC_14_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILL1NA_6_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILL1NA_6_LC_14_7_1 .LUT_INIT=16'b1000000010000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILL1NA_6_LC_14_7_1  (
            .in0(N__47470),
            .in1(N__34230),
            .in2(N__34184),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_358 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_14_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_14_7_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_14_7_2  (
            .in0(N__34318),
            .in1(N__41896),
            .in2(N__34367),
            .in3(N__37392),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_345 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_345_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_14_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_14_7_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_14_7_3 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_14_7_3  (
            .in0(N__35386),
            .in1(N__37720),
            .in2(N__34175),
            .in3(N__35200),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_348 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_14_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_14_7_5 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_14_7_5  (
            .in0(N__39574),
            .in1(N__41820),
            .in2(N__40079),
            .in3(N__34319),
            .lcout(elapsed_time_ns_1_RNIAE2591_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_16_LC_14_7_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_16_LC_14_7_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_16_LC_14_7_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_16_LC_14_7_7  (
            .in0(N__34475),
            .in1(N__34446),
            .in2(N__34253),
            .in3(N__34405),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_381 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_14_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_14_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_14_8_0  (
            .in0(N__40127),
            .in1(N__34271),
            .in2(N__37903),
            .in3(N__35193),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_14_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_14_8_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_14_8_1  (
            .in0(N__34207),
            .in1(N__37687),
            .in2(N__35107),
            .in3(N__41877),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_367 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_14_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_14_8_2 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_14_8_2  (
            .in0(N__35103),
            .in1(N__34208),
            .in2(N__37393),
            .in3(N__34317),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_16_LC_14_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_16_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_16_LC_14_8_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_16_LC_14_8_3  (
            .in0(N__34169),
            .in1(N__41878),
            .in2(N__34172),
            .in3(N__34366),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_380 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGE841_17_LC_14_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGE841_17_LC_14_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGE841_17_LC_14_8_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGE841_17_LC_14_8_4  (
            .in0(N__37686),
            .in1(N__40131),
            .in2(N__37902),
            .in3(N__35192),
            .lcout(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_14_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_14_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_14_8_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_14_8_5  (
            .in0(_gnd_net_),
            .in1(N__35119),
            .in2(_gnd_net_),
            .in3(N__37657),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_341 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_14_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_14_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_14_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_14_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34351),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47836),
            .ce(N__34301),
            .sr(N__47301));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO7LR2_9_LC_14_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO7LR2_9_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO7LR2_9_LC_14_9_1 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO7LR2_9_LC_14_9_1  (
            .in0(N__40132),
            .in1(N__34457),
            .in2(_gnd_net_),
            .in3(N__34280),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_349_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3GEH5_15_LC_14_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3GEH5_15_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3GEH5_15_LC_14_9_2 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3GEH5_15_LC_14_9_2  (
            .in0(N__40096),
            .in1(N__34270),
            .in2(N__34259),
            .in3(N__37889),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_363_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_14_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_14_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_14_9_3 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_14_9_3  (
            .in0(N__38167),
            .in1(N__34406),
            .in2(N__34256),
            .in3(N__34473),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_16_LC_14_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_16_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_16_LC_14_9_4 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_16_LC_14_9_4  (
            .in0(N__34447),
            .in1(N__34252),
            .in2(N__34238),
            .in3(N__47471),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_14_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_14_9_5 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_14_9_5  (
            .in0(N__47472),
            .in1(N__34232),
            .in2(N__34235),
            .in3(N__38170),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_14_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_14_9_6 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_14_9_6  (
            .in0(N__34231),
            .in1(N__34217),
            .in2(N__35153),
            .in3(N__38168),
            .lcout(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ),
            .ltout(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_14_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_14_9_7 .LUT_INIT=16'b1111111111001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_14_9_7  (
            .in0(N__38245),
            .in1(N__34201),
            .in2(N__34187),
            .in3(N__41555),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_14_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_14_10_1 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_14_10_1  (
            .in0(N__35222),
            .in1(N__34424),
            .in2(N__41754),
            .in3(N__40038),
            .lcout(elapsed_time_ns_1_RNI1HIF91_0_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_14_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_14_10_2 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_14_10_2  (
            .in0(N__40039),
            .in1(N__34484),
            .in2(N__41769),
            .in3(N__37963),
            .lcout(elapsed_time_ns_1_RNIQ9IF91_0_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_14_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_14_10_3 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_14_10_3  (
            .in0(N__41700),
            .in1(N__35447),
            .in2(N__40068),
            .in3(N__34498),
            .lcout(elapsed_time_ns_1_RNI0GIF91_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIME943_20_LC_14_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIME943_20_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIME943_20_LC_14_10_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIME943_20_LC_14_10_4  (
            .in0(N__35239),
            .in1(N__34373),
            .in2(N__34499),
            .in3(N__34483),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_14_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_14_10_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_14_10_5  (
            .in0(N__35356),
            .in1(N__35398),
            .in2(N__35335),
            .in3(N__35278),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_347 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_347_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_7_LC_14_10_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_7_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_7_LC_14_10_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_7_LC_14_10_6  (
            .in0(N__40095),
            .in1(N__35382),
            .in2(N__34451),
            .in3(N__37716),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_365 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_14_10_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_14_10_7 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_14_10_7  (
            .in0(N__34535),
            .in1(N__34385),
            .in2(N__41753),
            .in3(N__40037),
            .lcout(elapsed_time_ns_1_RNIUDIF91_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_14_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_14_11_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_14_11_2  (
            .in0(N__35257),
            .in1(N__35425),
            .in2(N__34423),
            .in3(N__35164),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_14_11_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_14_11_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_14_11_3  (
            .in0(N__38014),
            .in1(N__38032),
            .in2(N__34562),
            .in3(N__34384),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_14_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_14_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_14_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36452),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_14_11_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_14_11_5 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_14_11_5  (
            .in0(N__41721),
            .in1(N__34561),
            .in2(N__34547),
            .in3(N__40052),
            .lcout(elapsed_time_ns_1_RNITCIF91_0_23),
            .ltout(elapsed_time_ns_1_RNITCIF91_0_23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_15_LC_14_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_15_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_15_LC_14_11_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_15_LC_14_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34538),
            .in3(N__34534),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_14_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_14_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_14_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36482),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_14_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_14_12_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_0_LC_14_12_1  (
            .in0(_gnd_net_),
            .in1(N__34509),
            .in2(_gnd_net_),
            .in3(N__36189),
            .lcout(),
            .ltout(\phase_controller_inst1.N_55_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_LC_14_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_14_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_14_12_2 .LUT_INIT=16'b1010101110101010;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_14_12_2  (
            .in0(N__37484),
            .in1(N__34828),
            .in2(N__34514),
            .in3(N__36220),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47813),
            .ce(),
            .sr(N__47320));
    defparam \phase_controller_inst1.state_2_LC_14_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_14_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_14_12_3 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_inst1.state_2_LC_14_12_3  (
            .in0(N__37520),
            .in1(N__34510),
            .in2(N__37565),
            .in3(N__36190),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47813),
            .ce(),
            .sr(N__47320));
    defparam \phase_controller_inst1.state_1_LC_14_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_14_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_14_12_4 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \phase_controller_inst1.state_1_LC_14_12_4  (
            .in0(N__34511),
            .in1(N__36191),
            .in2(N__38427),
            .in3(N__38395),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47813),
            .ce(),
            .sr(N__47320));
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_14_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_14_12_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_RNO_0_LC_14_12_5  (
            .in0(_gnd_net_),
            .in1(N__38417),
            .in2(_gnd_net_),
            .in3(N__38394),
            .lcout(),
            .ltout(\phase_controller_inst1.start_timer_tr_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_tr_LC_14_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_14_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_14_12_6 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_14_12_6  (
            .in0(N__38353),
            .in1(N__43020),
            .in2(N__34832),
            .in3(N__34829),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47813),
            .ce(),
            .sr(N__47320));
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_14_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_14_12_7 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_14_12_7  (
            .in0(N__42958),
            .in1(N__42907),
            .in2(_gnd_net_),
            .in3(N__43016),
            .lcout(\phase_controller_inst1.stoper_tr.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_14_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_14_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_14_13_1 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_LC_14_13_1  (
            .in0(N__34682),
            .in1(N__34761),
            .in2(N__34778),
            .in3(N__34717),
            .lcout(\phase_controller_inst2.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47807),
            .ce(),
            .sr(N__47325));
    defparam \phase_controller_inst2.stoper_tr.running_LC_14_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_LC_14_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.running_LC_14_13_3 .LUT_INIT=16'b1010001010101110;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_LC_14_13_3  (
            .in0(N__34736),
            .in1(N__34585),
            .in2(N__34745),
            .in3(N__34718),
            .lcout(\phase_controller_inst2.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47807),
            .ce(),
            .sr(N__47325));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNIP8O21_LC_14_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNIP8O21_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNIP8O21_LC_14_13_6 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNIP8O21_LC_14_13_6  (
            .in0(N__34716),
            .in1(N__34681),
            .in2(_gnd_net_),
            .in3(N__35539),
            .lcout(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_14_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_14_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_14_13_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_14_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34601),
            .in3(N__34584),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__34963),
            .in2(N__38324),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(N__43797),
            .in2(N__43835),
            .in3(N__38577),
            .lcout(\current_shift_inst.un38_control_input_5_1 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_14_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_14_2  (
            .in0(N__38578),
            .in1(N__44848),
            .in2(N__40679),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un38_control_input_5_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_14_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_14_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(N__34859),
            .in2(N__45041),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_14_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_14_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(N__44852),
            .in2(N__38309),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_14_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_14_14_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(N__38297),
            .in2(N__45042),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_14_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_14_14_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(N__44856),
            .in2(N__38477),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_14_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_14_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_LC_14_14_7  (
            .in0(_gnd_net_),
            .in1(N__38486),
            .in2(N__45043),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_14_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_14_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__38447),
            .in2(N__45044),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_14_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_14_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(N__44863),
            .in2(N__34850),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_14_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_14_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(N__43895),
            .in2(N__45045),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_14_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_14_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_LC_14_15_3  (
            .in0(_gnd_net_),
            .in1(N__44867),
            .in2(N__34841),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_14_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_14_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_LC_14_15_4  (
            .in0(_gnd_net_),
            .in1(N__34877),
            .in2(N__45046),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_14_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_14_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_LC_14_15_5  (
            .in0(_gnd_net_),
            .in1(N__44871),
            .in2(N__45401),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_14_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_14_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_LC_14_15_6  (
            .in0(_gnd_net_),
            .in1(N__34871),
            .in2(N__45047),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_14_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_14_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_LC_14_15_7  (
            .in0(_gnd_net_),
            .in1(N__44875),
            .in2(N__43475),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_14_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_14_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_LC_14_16_0  (
            .in0(_gnd_net_),
            .in1(N__44964),
            .in2(N__43199),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_14_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_14_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(N__43625),
            .in2(N__45132),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_14_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_14_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_LC_14_16_2  (
            .in0(_gnd_net_),
            .in1(N__44968),
            .in2(N__41129),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_14_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_14_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_LC_14_16_3  (
            .in0(_gnd_net_),
            .in1(N__34865),
            .in2(N__45133),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(N__44972),
            .in2(N__36650),
            .in3(N__34940),
            .lcout(\current_shift_inst.un38_control_input_0_s0_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(N__34937),
            .in2(N__45134),
            .in3(N__34928),
            .lcout(\current_shift_inst.un38_control_input_0_s0_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_16_6  (
            .in0(_gnd_net_),
            .in1(N__44976),
            .in2(N__36623),
            .in3(N__34925),
            .lcout(\current_shift_inst.un38_control_input_0_s0_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_16_7  (
            .in0(_gnd_net_),
            .in1(N__36614),
            .in2(N__45135),
            .in3(N__34922),
            .lcout(\current_shift_inst.un38_control_input_0_s0_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_17_0  (
            .in0(_gnd_net_),
            .in1(N__45010),
            .in2(N__45347),
            .in3(N__34919),
            .lcout(\current_shift_inst.un38_control_input_0_s0_24 ),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(N__34916),
            .in2(N__45143),
            .in3(N__34910),
            .lcout(\current_shift_inst.un38_control_input_0_s0_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(N__45014),
            .in2(N__44177),
            .in3(N__34907),
            .lcout(\current_shift_inst.un38_control_input_0_s0_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_17_3  (
            .in0(_gnd_net_),
            .in1(N__34904),
            .in2(N__45144),
            .in3(N__34895),
            .lcout(\current_shift_inst.un38_control_input_0_s0_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_17_4  (
            .in0(_gnd_net_),
            .in1(N__45018),
            .in2(N__34892),
            .in3(N__34880),
            .lcout(\current_shift_inst.un38_control_input_0_s0_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_17_5  (
            .in0(_gnd_net_),
            .in1(N__44129),
            .in2(N__45145),
            .in3(N__34982),
            .lcout(\current_shift_inst.un38_control_input_0_s0_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_14_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_14_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_14_17_6  (
            .in0(_gnd_net_),
            .in1(N__45022),
            .in2(N__44243),
            .in3(N__34979),
            .lcout(\current_shift_inst.un38_control_input_0_s0_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_RNO_0_11_LC_14_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_RNO_0_11_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_RNO_0_11_LC_14_17_7 .LUT_INIT=16'b1100010100110101;
    LogicCell40 \current_shift_inst.control_input_RNO_0_11_LC_14_17_7  (
            .in0(N__35027),
            .in1(N__34976),
            .in2(N__38747),
            .in3(N__34967),
            .lcout(\current_shift_inst.control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_14_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_14_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(N__34964),
            .in2(N__40636),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_14_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_14_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(N__43801),
            .in2(N__43778),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_14_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_14_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_LC_14_18_2  (
            .in0(_gnd_net_),
            .in1(N__44936),
            .in2(N__40664),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_14_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_14_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(N__34946),
            .in2(N__45125),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_14_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_14_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(N__44940),
            .in2(N__43232),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_14_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_14_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(N__38498),
            .in2(N__45126),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_14_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_14_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_LC_14_18_6  (
            .in0(_gnd_net_),
            .in1(N__44944),
            .in2(N__38465),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_14_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_14_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_LC_14_18_7  (
            .in0(_gnd_net_),
            .in1(N__38270),
            .in2(N__45127),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_14_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_14_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_LC_14_19_0  (
            .in0(_gnd_net_),
            .in1(N__44948),
            .in2(N__38288),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_19_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_14_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_14_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_LC_14_19_1  (
            .in0(_gnd_net_),
            .in1(N__41225),
            .in2(N__45128),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_14_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_14_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_LC_14_19_2  (
            .in0(_gnd_net_),
            .in1(N__44952),
            .in2(N__44114),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_14_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_14_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_LC_14_19_3  (
            .in0(_gnd_net_),
            .in1(N__37277),
            .in2(N__45129),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_14_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_14_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_LC_14_19_4  (
            .in0(_gnd_net_),
            .in1(N__44956),
            .in2(N__43586),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_14_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_14_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(N__41297),
            .in2(N__45130),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_14_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_14_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_LC_14_19_6  (
            .in0(_gnd_net_),
            .in1(N__44960),
            .in2(N__43526),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_14_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_14_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_LC_14_19_7  (
            .in0(_gnd_net_),
            .in1(N__37262),
            .in2(N__45131),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_14_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_14_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_LC_14_20_0  (
            .in0(_gnd_net_),
            .in1(N__37283),
            .in2(N__45136),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_20_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_14_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_14_20_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(N__44983),
            .in2(N__37271),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_14_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_14_20_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_LC_14_20_2  (
            .in0(_gnd_net_),
            .in1(N__41039),
            .in2(N__45137),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_14_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_14_20_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_LC_14_20_3  (
            .in0(_gnd_net_),
            .in1(N__44987),
            .in2(N__35018),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_14_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_14_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_14_20_4  (
            .in0(_gnd_net_),
            .in1(N__36767),
            .in2(N__45138),
            .in3(N__35003),
            .lcout(\current_shift_inst.un38_control_input_0_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_14_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_14_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_14_20_5  (
            .in0(_gnd_net_),
            .in1(N__44991),
            .in2(N__35000),
            .in3(N__34991),
            .lcout(\current_shift_inst.un38_control_input_0_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_14_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_14_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_14_20_6  (
            .in0(_gnd_net_),
            .in1(N__39098),
            .in2(N__45139),
            .in3(N__34988),
            .lcout(\current_shift_inst.un38_control_input_0_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_14_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_14_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_14_20_7  (
            .in0(_gnd_net_),
            .in1(N__44995),
            .in2(N__37637),
            .in3(N__34985),
            .lcout(\current_shift_inst.un38_control_input_0_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_14_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_14_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_14_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_14_21_0  (
            .in0(_gnd_net_),
            .in1(N__44996),
            .in2(N__45446),
            .in3(N__35069),
            .lcout(\current_shift_inst.un38_control_input_0_s1_24 ),
            .ltout(),
            .carryin(bfn_14_21_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_14_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_14_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_14_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_14_21_1  (
            .in0(_gnd_net_),
            .in1(N__44306),
            .in2(N__45140),
            .in3(N__35066),
            .lcout(\current_shift_inst.un38_control_input_0_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_14_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_14_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_14_21_2  (
            .in0(_gnd_net_),
            .in1(N__45000),
            .in2(N__35063),
            .in3(N__35054),
            .lcout(\current_shift_inst.un38_control_input_0_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_14_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_14_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_14_21_3  (
            .in0(_gnd_net_),
            .in1(N__40409),
            .in2(N__45141),
            .in3(N__35051),
            .lcout(\current_shift_inst.un38_control_input_0_s1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_14_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_14_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_14_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_14_21_4  (
            .in0(_gnd_net_),
            .in1(N__45004),
            .in2(N__35048),
            .in3(N__35039),
            .lcout(\current_shift_inst.un38_control_input_0_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_14_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_14_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_14_21_5  (
            .in0(_gnd_net_),
            .in1(N__39110),
            .in2(N__45142),
            .in3(N__35036),
            .lcout(\current_shift_inst.un38_control_input_0_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_14_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_14_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_14_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_14_21_6  (
            .in0(_gnd_net_),
            .in1(N__45008),
            .in2(N__44242),
            .in3(N__35033),
            .lcout(\current_shift_inst.un38_control_input_0_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_RNO_2_11_LC_14_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_RNO_2_11_LC_14_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_RNO_2_11_LC_14_21_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \current_shift_inst.control_input_RNO_2_11_LC_14_21_7  (
            .in0(N__45009),
            .in1(N__44646),
            .in2(_gnd_net_),
            .in3(N__35030),
            .lcout(\current_shift_inst.un38_control_input_0_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.S1_LC_14_22_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_14_22_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_14_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S1_LC_14_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37551),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47765),
            .ce(),
            .sr(N__47384));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_15_4_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_15_4_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_15_4_1 .LUT_INIT=16'b1111111011001110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_15_4_1  (
            .in0(N__42695),
            .in1(N__41582),
            .in2(N__41821),
            .in3(N__35207),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_15_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_15_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_15_7_0 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_15_7_0  (
            .in0(N__35174),
            .in1(N__37996),
            .in2(N__41825),
            .in3(N__40076),
            .lcout(elapsed_time_ns_1_RNIRBJF91_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2_1_LC_15_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2_1_LC_15_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2_1_LC_15_7_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2_1_LC_15_7_1  (
            .in0(_gnd_net_),
            .in1(N__42154),
            .in2(_gnd_net_),
            .in3(N__39564),
            .lcout(\phase_controller_inst1.stoper_tr.N_219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAKOL_31_LC_15_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAKOL_31_LC_15_7_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAKOL_31_LC_15_7_3 .LUT_INIT=16'b1111111110101000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAKOL_31_LC_15_7_3  (
            .in0(N__47469),
            .in1(N__35146),
            .in2(N__38174),
            .in3(N__35135),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFG4DM1_16_LC_15_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFG4DM1_16_LC_15_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFG4DM1_16_LC_15_7_4 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFG4DM1_16_LC_15_7_4  (
            .in0(N__41516),
            .in1(_gnd_net_),
            .in2(N__35129),
            .in3(_gnd_net_),
            .lcout(elapsed_time_ns_1_RNIFG4DM1_0_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_15_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_15_7_5 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_15_7_5  (
            .in0(N__40077),
            .in1(N__42366),
            .in2(N__41796),
            .in3(N__35126),
            .lcout(elapsed_time_ns_1_RNIDH2591_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIJ4DM1_19_LC_15_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIJ4DM1_19_LC_15_7_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIJ4DM1_19_LC_15_7_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIJ4DM1_19_LC_15_7_6  (
            .in0(_gnd_net_),
            .in1(N__35075),
            .in2(_gnd_net_),
            .in3(N__41496),
            .lcout(elapsed_time_ns_1_RNIIJ4DM1_0_19),
            .ltout(elapsed_time_ns_1_RNIIJ4DM1_0_19_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_15_7_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_15_7_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_15_7_7 .LUT_INIT=16'b1111111111011000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_15_7_7  (
            .in0(N__41743),
            .in1(N__35108),
            .in2(N__35078),
            .in3(N__41561),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_15_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_15_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_15_8_0 .LUT_INIT=16'b0011001100110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_14_LC_15_8_0  (
            .in0(N__38093),
            .in1(N__42527),
            .in2(N__39896),
            .in3(N__39735),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47845),
            .ce(N__43373),
            .sr(N__47294));
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_15_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_15_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_15_8_1 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_10_LC_15_8_1  (
            .in0(N__42523),
            .in1(N__37769),
            .in2(N__39764),
            .in3(N__38094),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47845),
            .ce(N__43373),
            .sr(N__47294));
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_15_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_15_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_15_8_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_11_LC_15_8_2  (
            .in0(N__38091),
            .in1(N__42525),
            .in2(N__37799),
            .in3(N__39742),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47845),
            .ce(N__43373),
            .sr(N__47294));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_15_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_15_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_15_8_3 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_15_8_3  (
            .in0(N__35285),
            .in1(N__37816),
            .in2(N__41768),
            .in3(N__40045),
            .lcout(elapsed_time_ns_1_RNISAHF91_0_13),
            .ltout(elapsed_time_ns_1_RNISAHF91_0_13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_15_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_15_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_15_8_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_13_LC_15_8_4  (
            .in0(N__38092),
            .in1(N__42526),
            .in2(N__35267),
            .in3(N__39734),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47845),
            .ce(N__43373),
            .sr(N__47294));
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_15_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_15_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_15_8_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_12_LC_15_8_5  (
            .in0(N__42524),
            .in1(N__37743),
            .in2(N__39765),
            .in3(N__38095),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47845),
            .ce(N__43373),
            .sr(N__47294));
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_15_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_15_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_15_8_6 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_19_LC_15_8_6  (
            .in0(N__39732),
            .in1(N__42528),
            .in2(_gnd_net_),
            .in3(N__39271),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47845),
            .ce(N__43373),
            .sr(N__47294));
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_15_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_15_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_15_8_7 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_18_LC_15_8_7  (
            .in0(N__42529),
            .in1(N__38246),
            .in2(_gnd_net_),
            .in3(N__39733),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47845),
            .ce(N__43373),
            .sr(N__47294));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_15_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_15_9_0 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_15_9_0  (
            .in0(N__40035),
            .in1(N__35264),
            .in2(N__41770),
            .in3(N__37982),
            .lcout(elapsed_time_ns_1_RNI3JIF91_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_15_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_15_9_1 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_15_9_1  (
            .in0(N__35246),
            .in1(N__35228),
            .in2(N__41750),
            .in3(N__40030),
            .lcout(elapsed_time_ns_1_RNIVEIF91_0_25),
            .ltout(elapsed_time_ns_1_RNIVEIF91_0_25_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6_15_LC_15_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6_15_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6_15_LC_15_9_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6_15_LC_15_9_2  (
            .in0(N__35413),
            .in1(N__35221),
            .in2(N__35210),
            .in3(N__35446),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_15_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_15_9_3 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_15_9_3  (
            .in0(N__41685),
            .in1(N__35414),
            .in2(N__35435),
            .in3(N__40032),
            .lcout(elapsed_time_ns_1_RNI2IIF91_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_15_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_15_9_4 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_15_9_4  (
            .in0(N__40031),
            .in1(N__41689),
            .in2(N__35405),
            .in3(N__37771),
            .lcout(elapsed_time_ns_1_RNIP7HF91_0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_15_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_15_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_15_9_5 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_15_9_5  (
            .in0(N__39513),
            .in1(N__35387),
            .in2(N__41752),
            .in3(N__40036),
            .lcout(elapsed_time_ns_1_RNIGK2591_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_15_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_15_9_6 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_15_9_6  (
            .in0(N__40033),
            .in1(N__41690),
            .in2(N__35363),
            .in3(N__37745),
            .lcout(elapsed_time_ns_1_RNIR9HF91_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_15_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_15_9_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_15_9_7 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_15_9_7  (
            .in0(N__37798),
            .in1(N__35339),
            .in2(N__41751),
            .in3(N__40034),
            .lcout(elapsed_time_ns_1_RNIQ8HF91_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_1_c_inv_LC_15_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_1_c_inv_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_1_c_inv_LC_15_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_1_c_inv_LC_15_10_0  (
            .in0(_gnd_net_),
            .in1(N__39629),
            .in2(N__35318),
            .in3(N__35755),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_15_10_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_2_c_inv_LC_15_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_2_c_inv_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_2_c_inv_LC_15_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_2_c_inv_LC_15_10_1  (
            .in0(_gnd_net_),
            .in1(N__39599),
            .in2(N__35309),
            .in3(N__35717),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_3_c_inv_LC_15_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_3_c_inv_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_3_c_inv_LC_15_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_3_c_inv_LC_15_10_2  (
            .in0(_gnd_net_),
            .in1(N__42128),
            .in2(N__35297),
            .in3(N__35687),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_4_c_inv_LC_15_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_4_c_inv_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_4_c_inv_LC_15_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_4_c_inv_LC_15_10_3  (
            .in0(_gnd_net_),
            .in1(N__35528),
            .in2(N__42551),
            .in3(N__35669),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_5_c_inv_LC_15_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_5_c_inv_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_5_c_inv_LC_15_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_5_c_inv_LC_15_10_4  (
            .in0(_gnd_net_),
            .in1(N__42344),
            .in2(N__35522),
            .in3(N__35651),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_6_c_inv_LC_15_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_6_c_inv_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_6_c_inv_LC_15_10_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_6_c_inv_LC_15_10_5  (
            .in0(N__35633),
            .in1(N__39455),
            .in2(N__35510),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_7_c_inv_LC_15_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_7_c_inv_LC_15_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_7_c_inv_LC_15_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_7_c_inv_LC_15_10_6  (
            .in0(_gnd_net_),
            .in1(N__39209),
            .in2(N__35498),
            .in3(N__36110),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_8_c_inv_LC_15_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_8_c_inv_LC_15_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_8_c_inv_LC_15_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_8_c_inv_LC_15_10_7  (
            .in0(_gnd_net_),
            .in1(N__39611),
            .in2(N__35489),
            .in3(N__36092),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_9_c_inv_LC_15_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_9_c_inv_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_9_c_inv_LC_15_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_9_c_inv_LC_15_11_0  (
            .in0(_gnd_net_),
            .in1(N__38048),
            .in2(N__35477),
            .in3(N__36074),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_15_11_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_10_c_inv_LC_15_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_10_c_inv_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_10_c_inv_LC_15_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_10_c_inv_LC_15_11_1  (
            .in0(_gnd_net_),
            .in1(N__37862),
            .in2(N__35468),
            .in3(N__36056),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_11_c_inv_LC_15_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_11_c_inv_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_11_c_inv_LC_15_11_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_11_c_inv_LC_15_11_2  (
            .in0(N__36038),
            .in1(N__35459),
            .in2(N__37850),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_12_c_inv_LC_15_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_12_c_inv_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_12_c_inv_LC_15_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_12_c_inv_LC_15_11_3  (
            .in0(_gnd_net_),
            .in1(N__35453),
            .in2(N__37838),
            .in3(N__36020),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_13_c_inv_LC_15_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_13_c_inv_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_13_c_inv_LC_15_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_13_c_inv_LC_15_11_4  (
            .in0(_gnd_net_),
            .in1(N__37826),
            .in2(N__35615),
            .in3(N__36002),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_14_c_inv_LC_15_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_14_c_inv_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_14_c_inv_LC_15_11_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_14_c_inv_LC_15_11_5  (
            .in0(N__35981),
            .in1(N__37916),
            .in2(N__35606),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_15_c_inv_LC_15_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_15_c_inv_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_15_c_inv_LC_15_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_15_c_inv_LC_15_11_6  (
            .in0(_gnd_net_),
            .in1(N__39221),
            .in2(N__35594),
            .in3(N__35963),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_16_c_inv_LC_15_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_16_c_inv_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_16_c_inv_LC_15_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_16_c_inv_LC_15_11_7  (
            .in0(_gnd_net_),
            .in1(N__39236),
            .in2(N__35585),
            .in3(N__36392),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_17_c_inv_LC_15_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_17_c_inv_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_17_c_inv_LC_15_12_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_17_c_inv_LC_15_12_0  (
            .in0(N__36374),
            .in1(N__38180),
            .in2(N__35576),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_15_12_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_18_c_inv_LC_15_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_18_c_inv_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_18_c_inv_LC_15_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_18_c_inv_LC_15_12_1  (
            .in0(_gnd_net_),
            .in1(N__38210),
            .in2(N__35567),
            .in3(N__36356),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_inv_LC_15_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_inv_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_inv_LC_15_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_inv_LC_15_12_2  (
            .in0(_gnd_net_),
            .in1(N__39251),
            .in2(N__35558),
            .in3(N__36335),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_LUT4_0_LC_15_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_LUT4_0_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_LUT4_0_LC_15_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_LUT4_0_LC_15_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35549),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_15_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_15_12_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_15_12_4  (
            .in0(N__36137),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5LMJQ_9_LC_15_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5LMJQ_9_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5LMJQ_9_LC_15_12_5 .LUT_INIT=16'b1111101111101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5LMJQ_9_LC_15_12_5  (
            .in0(N__35929),
            .in1(N__36944),
            .in2(N__35855),
            .in3(N__35822),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_15_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_15_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_15_13_0  (
            .in0(_gnd_net_),
            .in1(N__35765),
            .in2(N__35759),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_13_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_15_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_15_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_15_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_15_13_1  (
            .in0(N__42069),
            .in1(N__35716),
            .in2(_gnd_net_),
            .in3(N__35702),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__47814),
            .ce(),
            .sr(N__47321));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_15_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_15_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_15_13_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_15_13_2  (
            .in0(N__42081),
            .in1(N__35686),
            .in2(N__35699),
            .in3(N__35672),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__47814),
            .ce(),
            .sr(N__47321));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_15_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_15_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_15_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_15_13_3  (
            .in0(N__42070),
            .in1(N__35668),
            .in2(_gnd_net_),
            .in3(N__35654),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__47814),
            .ce(),
            .sr(N__47321));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_15_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_15_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_15_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_15_13_4  (
            .in0(N__42082),
            .in1(N__35650),
            .in2(_gnd_net_),
            .in3(N__35636),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__47814),
            .ce(),
            .sr(N__47321));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_15_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_15_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_15_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_15_13_5  (
            .in0(N__42071),
            .in1(N__35632),
            .in2(_gnd_net_),
            .in3(N__35618),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__47814),
            .ce(),
            .sr(N__47321));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_15_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_15_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_15_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_15_13_6  (
            .in0(N__42083),
            .in1(N__36109),
            .in2(_gnd_net_),
            .in3(N__36095),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__47814),
            .ce(),
            .sr(N__47321));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_15_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_15_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_15_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_15_13_7  (
            .in0(N__42072),
            .in1(N__36091),
            .in2(_gnd_net_),
            .in3(N__36077),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__47814),
            .ce(),
            .sr(N__47321));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_15_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_15_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_15_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_15_14_0  (
            .in0(N__42097),
            .in1(N__36073),
            .in2(_gnd_net_),
            .in3(N__36059),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_15_14_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__47808),
            .ce(),
            .sr(N__47326));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_15_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_15_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_15_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_15_14_1  (
            .in0(N__42089),
            .in1(N__36055),
            .in2(_gnd_net_),
            .in3(N__36041),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__47808),
            .ce(),
            .sr(N__47326));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_15_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_15_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_15_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_15_14_2  (
            .in0(N__42094),
            .in1(N__36037),
            .in2(_gnd_net_),
            .in3(N__36023),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__47808),
            .ce(),
            .sr(N__47326));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_15_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_15_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_15_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_15_14_3  (
            .in0(N__42090),
            .in1(N__36019),
            .in2(_gnd_net_),
            .in3(N__36005),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__47808),
            .ce(),
            .sr(N__47326));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_15_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_15_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_15_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_15_14_4  (
            .in0(N__42095),
            .in1(N__35998),
            .in2(_gnd_net_),
            .in3(N__35984),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__47808),
            .ce(),
            .sr(N__47326));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_15_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_15_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_15_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_15_14_5  (
            .in0(N__42091),
            .in1(N__35980),
            .in2(_gnd_net_),
            .in3(N__35966),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__47808),
            .ce(),
            .sr(N__47326));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_15_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_15_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_15_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_15_14_6  (
            .in0(N__42096),
            .in1(N__35959),
            .in2(_gnd_net_),
            .in3(N__35945),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__47808),
            .ce(),
            .sr(N__47326));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_15_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_15_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_15_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_15_14_7  (
            .in0(N__42092),
            .in1(N__36391),
            .in2(_gnd_net_),
            .in3(N__36377),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__47808),
            .ce(),
            .sr(N__47326));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_15_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_15_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_15_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_15_15_0  (
            .in0(N__42087),
            .in1(N__36373),
            .in2(_gnd_net_),
            .in3(N__36359),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_15_15_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__47802),
            .ce(),
            .sr(N__47329));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_15_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_15_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_15_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_15_15_1  (
            .in0(N__42093),
            .in1(N__36355),
            .in2(_gnd_net_),
            .in3(N__36341),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__47802),
            .ce(),
            .sr(N__47329));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_15_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_15_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_15_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_15_15_2  (
            .in0(N__42088),
            .in1(N__36334),
            .in2(_gnd_net_),
            .in3(N__36338),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47802),
            .ce(),
            .sr(N__47329));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_15_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_15_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_15_15_6 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_15_15_6  (
            .in0(N__36320),
            .in1(N__36308),
            .in2(N__36251),
            .in3(N__36180),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47802),
            .ce(),
            .sr(N__47329));
    defparam \current_shift_inst.control_input_0_LC_15_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_0_LC_15_16_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_0_LC_15_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_0_LC_15_16_0  (
            .in0(_gnd_net_),
            .in1(N__36779),
            .in2(N__36638),
            .in3(N__36637),
            .lcout(\current_shift_inst.control_inputZ0Z_0 ),
            .ltout(),
            .carryin(bfn_15_16_0_),
            .carryout(\current_shift_inst.control_input_1_cry_0 ),
            .clk(N__47796),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_1_LC_15_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_1_LC_15_16_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_1_LC_15_16_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.control_input_1_LC_15_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36746),
            .in3(N__36128),
            .lcout(\current_shift_inst.control_inputZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_0 ),
            .carryout(\current_shift_inst.control_input_1_cry_1 ),
            .clk(N__47796),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_2_LC_15_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_2_LC_15_16_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_2_LC_15_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_2_LC_15_16_2  (
            .in0(_gnd_net_),
            .in1(N__36719),
            .in2(_gnd_net_),
            .in3(N__36113),
            .lcout(\current_shift_inst.control_inputZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_1 ),
            .carryout(\current_shift_inst.control_input_1_cry_2 ),
            .clk(N__47796),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_3_LC_15_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_3_LC_15_16_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_3_LC_15_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_3_LC_15_16_3  (
            .in0(_gnd_net_),
            .in1(N__36692),
            .in2(_gnd_net_),
            .in3(N__36500),
            .lcout(\current_shift_inst.control_inputZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_2 ),
            .carryout(\current_shift_inst.control_input_1_cry_3 ),
            .clk(N__47796),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_4_LC_15_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_4_LC_15_16_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_4_LC_15_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_4_LC_15_16_4  (
            .in0(_gnd_net_),
            .in1(N__37349),
            .in2(_gnd_net_),
            .in3(N__36485),
            .lcout(\current_shift_inst.control_inputZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_3 ),
            .carryout(\current_shift_inst.control_input_1_cry_4 ),
            .clk(N__47796),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_5_LC_15_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_5_LC_15_16_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_5_LC_15_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_5_LC_15_16_5  (
            .in0(_gnd_net_),
            .in1(N__37322),
            .in2(_gnd_net_),
            .in3(N__36470),
            .lcout(\current_shift_inst.control_inputZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_4 ),
            .carryout(\current_shift_inst.control_input_1_cry_5 ),
            .clk(N__47796),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_6_LC_15_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_6_LC_15_16_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_6_LC_15_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_6_LC_15_16_6  (
            .in0(_gnd_net_),
            .in1(N__37292),
            .in2(_gnd_net_),
            .in3(N__36455),
            .lcout(\current_shift_inst.control_inputZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_5 ),
            .carryout(\current_shift_inst.control_input_1_cry_6 ),
            .clk(N__47796),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_7_LC_15_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_7_LC_15_16_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_7_LC_15_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_7_LC_15_16_7  (
            .in0(_gnd_net_),
            .in1(N__36593),
            .in2(_gnd_net_),
            .in3(N__36440),
            .lcout(\current_shift_inst.control_inputZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_6 ),
            .carryout(\current_shift_inst.control_input_1_cry_7 ),
            .clk(N__47796),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_8_LC_15_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_8_LC_15_17_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_8_LC_15_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_8_LC_15_17_0  (
            .in0(_gnd_net_),
            .in1(N__36566),
            .in2(_gnd_net_),
            .in3(N__36425),
            .lcout(\current_shift_inst.control_inputZ0Z_8 ),
            .ltout(),
            .carryin(bfn_15_17_0_),
            .carryout(\current_shift_inst.control_input_1_cry_8 ),
            .clk(N__47791),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_9_LC_15_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_9_LC_15_17_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_9_LC_15_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_9_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(N__36542),
            .in2(_gnd_net_),
            .in3(N__36410),
            .lcout(\current_shift_inst.control_inputZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_8 ),
            .carryout(\current_shift_inst.control_input_1_cry_9 ),
            .clk(N__47791),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_10_LC_15_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_10_LC_15_17_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_10_LC_15_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_10_LC_15_17_2  (
            .in0(_gnd_net_),
            .in1(N__36518),
            .in2(_gnd_net_),
            .in3(N__36395),
            .lcout(\current_shift_inst.control_inputZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_9 ),
            .carryout(\current_shift_inst.control_input_1_cry_10 ),
            .clk(N__47791),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_11_LC_15_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_11_LC_15_17_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_11_LC_15_17_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.control_input_11_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(N__36683),
            .in2(_gnd_net_),
            .in3(N__36674),
            .lcout(\current_shift_inst.control_inputZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47791),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_17_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_17_4  (
            .in0(N__44618),
            .in1(N__46817),
            .in2(N__45202),
            .in3(N__41071),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_15_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_15_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38740),
            .lcout(\current_shift_inst.N_1609_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_15_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_15_17_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_15_17_6  (
            .in0(N__44619),
            .in1(N__46692),
            .in2(N__45201),
            .in3(N__40942),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_15_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_15_17_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_15_17_7  (
            .in0(N__45098),
            .in1(N__44620),
            .in2(N__46628),
            .in3(N__40911),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_15_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_15_18_0 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_15_18_0  (
            .in0(N__36608),
            .in1(N__36602),
            .in2(_gnd_net_),
            .in3(N__38733),
            .lcout(\current_shift_inst.control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_15_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_15_18_1 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_15_18_1  (
            .in0(N__38734),
            .in1(N__36584),
            .in2(_gnd_net_),
            .in3(N__36572),
            .lcout(\current_shift_inst.control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_15_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_15_18_2 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_15_18_2  (
            .in0(N__36560),
            .in1(N__36554),
            .in2(_gnd_net_),
            .in3(N__38735),
            .lcout(\current_shift_inst.control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_15_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_15_18_3 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_15_18_3  (
            .in0(N__38736),
            .in1(N__36536),
            .in2(_gnd_net_),
            .in3(N__36524),
            .lcout(\current_shift_inst.control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI81DJ11_2_LC_15_18_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI81DJ11_2_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI81DJ11_2_LC_15_18_4 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI81DJ11_2_LC_15_18_4  (
            .in0(N__37157),
            .in1(N__36998),
            .in2(N__37200),
            .in3(N__37243),
            .lcout(elapsed_time_ns_1_RNI81DJ11_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_18_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_18_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_18_5  (
            .in0(N__37229),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47786),
            .ce(N__37178),
            .sr(N__47339));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO1ND11_20_LC_15_18_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO1ND11_20_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO1ND11_20_LC_15_18_6 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO1ND11_20_LC_15_18_6  (
            .in0(N__37156),
            .in1(N__36808),
            .in2(N__37025),
            .in3(N__36997),
            .lcout(elapsed_time_ns_1_RNIO1ND11_0_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_15_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_15_19_0 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_15_19_0  (
            .in0(N__36794),
            .in1(N__36785),
            .in2(_gnd_net_),
            .in3(N__38723),
            .lcout(\current_shift_inst.control_input_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_15_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_15_19_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_15_19_1  (
            .in0(N__46813),
            .in1(N__44653),
            .in2(N__45263),
            .in3(N__41075),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_15_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_15_19_2 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_15_19_2  (
            .in0(N__36761),
            .in1(N__38724),
            .in2(_gnd_net_),
            .in3(N__36752),
            .lcout(\current_shift_inst.control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_15_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_15_19_3 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_15_19_3  (
            .in0(N__38725),
            .in1(N__36734),
            .in2(_gnd_net_),
            .in3(N__36725),
            .lcout(\current_shift_inst.control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_15_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_15_19_4 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_15_19_4  (
            .in0(N__36707),
            .in1(N__36701),
            .in2(_gnd_net_),
            .in3(N__38726),
            .lcout(\current_shift_inst.control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_15_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_15_19_5 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_15_19_5  (
            .in0(N__38728),
            .in1(N__37367),
            .in2(_gnd_net_),
            .in3(N__37358),
            .lcout(\current_shift_inst.control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_15_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_15_19_6 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_15_19_6  (
            .in0(N__37340),
            .in1(N__37331),
            .in2(_gnd_net_),
            .in3(N__38727),
            .lcout(\current_shift_inst.control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_15_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_15_19_7 .LUT_INIT=16'b0000101001011111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_15_19_7  (
            .in0(N__38729),
            .in1(_gnd_net_),
            .in2(N__37313),
            .in3(N__37301),
            .lcout(\current_shift_inst.control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_15_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_15_20_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_15_20_0  (
            .in0(N__44649),
            .in1(N__45209),
            .in2(N__46112),
            .in3(N__43709),
            .lcout(\current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_15_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_15_20_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_15_20_2  (
            .in0(N__44065),
            .in1(N__46693),
            .in2(_gnd_net_),
            .in3(N__40943),
            .lcout(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_15_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_15_20_3 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_15_20_3  (
            .in0(N__45207),
            .in1(N__44647),
            .in2(N__41215),
            .in3(N__46423),
            .lcout(\current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_15_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_15_20_4 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_15_20_4  (
            .in0(N__44650),
            .in1(N__46054),
            .in2(N__43667),
            .in3(N__45210),
            .lcout(\current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_15_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_15_20_5 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_15_20_5  (
            .in0(N__46620),
            .in1(N__40912),
            .in2(_gnd_net_),
            .in3(N__44066),
            .lcout(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_15_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_15_20_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_15_20_6  (
            .in0(N__44648),
            .in1(N__45208),
            .in2(N__46169),
            .in3(N__43504),
            .lcout(\current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_15_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_15_20_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_15_20_7  (
            .in0(N__45206),
            .in1(N__44651),
            .in2(N__46627),
            .in3(N__40913),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.stop_timer_s1_LC_15_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_LC_15_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.stop_timer_s1_LC_15_21_0 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \current_shift_inst.stop_timer_s1_LC_15_21_0  (
            .in0(N__37543),
            .in1(N__37423),
            .in2(N__37459),
            .in3(N__37600),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47774),
            .ce(),
            .sr(N__47369));
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_15_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_15_21_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNII51H_LC_15_21_1  (
            .in0(_gnd_net_),
            .in1(N__39142),
            .in2(_gnd_net_),
            .in3(N__37418),
            .lcout(\current_shift_inst.timer_s1.N_166_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.start_timer_s1_LC_15_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_15_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.start_timer_s1_LC_15_21_3 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_15_21_3  (
            .in0(N__37599),
            .in1(N__37452),
            .in2(_gnd_net_),
            .in3(N__37547),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47774),
            .ce(),
            .sr(N__47369));
    defparam \phase_controller_inst1.state_3_LC_15_21_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_15_21_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_15_21_6 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \phase_controller_inst1.state_3_LC_15_21_6  (
            .in0(N__38357),
            .in1(N__37519),
            .in2(N__37552),
            .in3(N__37586),
            .lcout(state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47774),
            .ce(),
            .sr(N__47369));
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_15_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_15_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_15_21_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_1_LC_15_21_7  (
            .in0(_gnd_net_),
            .in1(N__37542),
            .in2(_gnd_net_),
            .in3(N__37518),
            .lcout(\phase_controller_inst1.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_15_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_15_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_15_22_5 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIEOIK_LC_15_22_5  (
            .in0(N__39143),
            .in1(N__37419),
            .in2(_gnd_net_),
            .in3(N__37451),
            .lcout(\current_shift_inst.timer_s1.N_167_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_LC_16_6_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_16_6_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_16_6_0 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_16_6_0  (
            .in0(N__37469),
            .in1(N__39126),
            .in2(_gnd_net_),
            .in3(N__37433),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47866),
            .ce(),
            .sr(N__47281));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKL65B1_3_LC_16_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKL65B1_3_LC_16_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKL65B1_3_LC_16_7_0 .LUT_INIT=16'b1111111011110010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKL65B1_3_LC_16_7_0  (
            .in0(N__42164),
            .in1(N__41803),
            .in2(N__41497),
            .in3(N__37397),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRHL2M1_3_LC_16_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRHL2M1_3_LC_16_7_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRHL2M1_3_LC_16_7_1 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRHL2M1_3_LC_16_7_1  (
            .in0(N__41584),
            .in1(_gnd_net_),
            .in2(N__37697),
            .in3(_gnd_net_),
            .lcout(elapsed_time_ns_1_RNIRHL2M1_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_16_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_16_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_16_7_2 .LUT_INIT=16'b1111110011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_16_7_2  (
            .in0(N__38195),
            .in1(N__41583),
            .in2(N__37694),
            .in3(N__41804),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGH4DM1_17_LC_16_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGH4DM1_17_LC_16_7_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGH4DM1_17_LC_16_7_3 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGH4DM1_17_LC_16_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37670),
            .in3(N__41480),
            .lcout(elapsed_time_ns_1_RNIGH4DM1_0_17),
            .ltout(elapsed_time_ns_1_RNIGH4DM1_0_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_9_LC_16_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_9_LC_16_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_9_LC_16_7_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_9_LC_16_7_4  (
            .in0(N__38238),
            .in1(N__41845),
            .in2(N__37667),
            .in3(N__39269),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_16_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_16_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_16_7_5 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_16_7_5  (
            .in0(N__42567),
            .in1(N__37664),
            .in2(N__41822),
            .in3(N__40075),
            .lcout(elapsed_time_ns_1_RNICG2591_0_4),
            .ltout(elapsed_time_ns_1_RNICG2591_0_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3_2_LC_16_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3_2_LC_16_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3_2_LC_16_7_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3_2_LC_16_7_6  (
            .in0(N__38196),
            .in1(N__41846),
            .in2(N__37646),
            .in3(N__42360),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_2_LC_16_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_2_LC_16_7_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_2_LC_16_7_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_2_LC_16_7_7  (
            .in0(N__39270),
            .in1(N__38237),
            .in2(N__37643),
            .in3(N__39946),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDE4DM1_14_LC_16_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDE4DM1_14_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDE4DM1_14_LC_16_8_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDE4DM1_14_LC_16_8_0  (
            .in0(_gnd_net_),
            .in1(N__37868),
            .in2(_gnd_net_),
            .in3(N__41479),
            .lcout(elapsed_time_ns_1_RNIDE4DM1_0_14),
            .ltout(elapsed_time_ns_1_RNIDE4DM1_0_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_10_LC_16_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_10_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_10_LC_16_8_1 .LUT_INIT=16'b0011001100110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_a2_10_LC_16_8_1  (
            .in0(_gnd_net_),
            .in1(N__39839),
            .in2(N__37640),
            .in3(N__39806),
            .lcout(\phase_controller_inst1.stoper_tr.N_241 ),
            .ltout(\phase_controller_inst1.stoper_tr.N_241_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_16_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_16_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_16_8_2 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_14_LC_16_8_2  (
            .in0(N__42520),
            .in1(N__39892),
            .in2(N__37919),
            .in3(N__39754),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47857),
            .ce(N__42116),
            .sr(N__47287));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_16_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_16_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_16_8_3 .LUT_INIT=16'b1111101011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_16_8_3  (
            .in0(N__41586),
            .in1(N__39891),
            .in2(N__37907),
            .in3(N__41809),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_16_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_16_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_16_8_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_10_LC_16_8_4  (
            .in0(N__42518),
            .in1(N__37770),
            .in2(N__38108),
            .in3(N__39752),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47857),
            .ce(N__42116),
            .sr(N__47287));
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_16_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_16_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_16_8_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_11_LC_16_8_5  (
            .in0(N__38089),
            .in1(N__42521),
            .in2(N__39766),
            .in3(N__37797),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47857),
            .ce(N__42116),
            .sr(N__47287));
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_16_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_16_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_16_8_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_12_LC_16_8_6  (
            .in0(N__42519),
            .in1(N__37744),
            .in2(N__38109),
            .in3(N__39753),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47857),
            .ce(N__42116),
            .sr(N__47287));
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_16_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_16_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_16_8_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_13_LC_16_8_7  (
            .in0(N__38090),
            .in1(N__42522),
            .in2(N__39767),
            .in3(N__37817),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47857),
            .ce(N__42116),
            .sr(N__47287));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_3_LC_16_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_3_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_3_LC_16_9_1 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_3_LC_16_9_1  (
            .in0(N__39477),
            .in1(N__42452),
            .in2(N__39756),
            .in3(N__39551),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_2_LC_16_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_2_LC_16_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_2_LC_16_9_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_2_LC_16_9_2  (
            .in0(N__37815),
            .in1(N__37793),
            .in2(N__37772),
            .in3(N__37742),
            .lcout(\phase_controller_inst1.stoper_tr.N_244 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_16_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_16_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_16_9_3 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_16_9_3  (
            .in0(N__37721),
            .in1(N__42621),
            .in2(N__41816),
            .in3(N__40059),
            .lcout(elapsed_time_ns_1_RNIFJ2591_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_16_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_16_9_4 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_16_9_4  (
            .in0(N__40058),
            .in1(N__37949),
            .in2(N__38042),
            .in3(N__41786),
            .lcout(elapsed_time_ns_1_RNISBIF91_0_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_16_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_16_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_16_9_5 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_16_9_5  (
            .in0(N__38021),
            .in1(N__38003),
            .in2(N__41815),
            .in3(N__40057),
            .lcout(elapsed_time_ns_1_RNIRAIF91_0_21),
            .ltout(elapsed_time_ns_1_RNIRAIF91_0_21_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7_15_LC_16_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7_15_LC_16_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7_15_LC_16_9_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7_15_LC_16_9_6  (
            .in0(N__37997),
            .in1(N__37981),
            .in2(N__37970),
            .in3(N__37967),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_15_LC_16_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_15_LC_16_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_15_LC_16_9_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_o5_15_LC_16_9_7  (
            .in0(N__37948),
            .in1(N__37940),
            .in2(N__37934),
            .in3(N__37931),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_16_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_16_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_16_10_0 .LUT_INIT=16'b0011001100110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_9_LC_16_10_0  (
            .in0(N__39755),
            .in1(N__38117),
            .in2(N__39925),
            .in3(N__38111),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47837),
            .ce(N__43367),
            .sr(N__47302));
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_16_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_16_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_16_10_1 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_17_LC_16_10_1  (
            .in0(N__39743),
            .in1(N__42510),
            .in2(_gnd_net_),
            .in3(N__38204),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47837),
            .ce(N__43367),
            .sr(N__47302));
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_16_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_16_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_16_10_2 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_16_LC_16_10_2  (
            .in0(N__41860),
            .in1(N__42450),
            .in2(_gnd_net_),
            .in3(N__39745),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47837),
            .ce(N__43367),
            .sr(N__47302));
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_16_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_16_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_16_10_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_15_LC_16_10_3  (
            .in0(N__39744),
            .in1(N__39845),
            .in2(N__39811),
            .in3(N__42511),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47837),
            .ce(N__43367),
            .sr(N__47302));
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_16_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_16_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_16_10_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_8_LC_16_10_4  (
            .in0(N__42289),
            .in1(N__42451),
            .in2(_gnd_net_),
            .in3(N__39509),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47837),
            .ce(N__43367),
            .sr(N__47302));
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_16_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_16_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_16_10_5 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_3_LC_16_10_5  (
            .in0(N__42231),
            .in1(N__42290),
            .in2(N__42332),
            .in3(N__42169),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47837),
            .ce(N__43367),
            .sr(N__47302));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0_9_LC_16_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0_9_LC_16_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0_9_LC_16_10_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0_9_LC_16_10_6  (
            .in0(N__39918),
            .in1(N__39802),
            .in2(_gnd_net_),
            .in3(N__39863),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHI4DM1_18_LC_16_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHI4DM1_18_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHI4DM1_18_LC_16_11_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHI4DM1_18_LC_16_11_2  (
            .in0(_gnd_net_),
            .in1(N__38258),
            .in2(_gnd_net_),
            .in3(N__41504),
            .lcout(elapsed_time_ns_1_RNIHI4DM1_0_18),
            .ltout(elapsed_time_ns_1_RNIHI4DM1_0_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_16_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_16_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_16_11_3 .LUT_INIT=16'b0000000011111010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_18_LC_16_11_3  (
            .in0(N__39758),
            .in1(_gnd_net_),
            .in2(N__38213),
            .in3(N__42433),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47829),
            .ce(N__42119),
            .sr(N__47306));
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_16_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_16_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_16_11_4 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_17_LC_16_11_4  (
            .in0(N__42432),
            .in1(N__38203),
            .in2(_gnd_net_),
            .in3(N__39760),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47829),
            .ce(N__42119),
            .sr(N__47306));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_16_11_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_16_11_5 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_16_11_5  (
            .in0(N__38169),
            .in1(N__42431),
            .in2(N__41823),
            .in3(N__40078),
            .lcout(elapsed_time_ns_1_RNISCJF91_0_31),
            .ltout(elapsed_time_ns_1_RNISCJF91_0_31_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1_9_LC_16_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1_9_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1_9_LC_16_11_6 .LUT_INIT=16'b1111000011111110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1_9_LC_16_11_6  (
            .in0(N__38126),
            .in1(N__39950),
            .in2(N__38120),
            .in3(N__39757),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_16_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_16_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_16_11_7 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_9_LC_16_11_7  (
            .in0(N__39759),
            .in1(N__38110),
            .in2(N__38051),
            .in3(N__39926),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47829),
            .ce(N__42119),
            .sr(N__47306));
    defparam \phase_controller_inst1.state_0_LC_16_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_16_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_16_12_0 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \phase_controller_inst1.state_0_LC_16_12_0  (
            .in0(N__38335),
            .in1(N__38428),
            .in2(N__38369),
            .in3(N__38399),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47824),
            .ce(),
            .sr(N__47312));
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_16_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_16_12_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNI7NN7_0_LC_16_12_1  (
            .in0(_gnd_net_),
            .in1(N__38334),
            .in2(_gnd_net_),
            .in3(N__38365),
            .lcout(\phase_controller_inst1.N_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_16_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_16_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_16_12_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_16_12_2  (
            .in0(N__38336),
            .in1(N__43024),
            .in2(N__42975),
            .in3(N__42878),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47824),
            .ce(),
            .sr(N__47312));
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_16_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_16_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_16_12_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_LC_16_12_3  (
            .in0(_gnd_net_),
            .in1(N__43023),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47824),
            .ce(),
            .sr(N__47312));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_16_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_16_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_16_12_5 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_16_12_5  (
            .in0(N__42840),
            .in1(N__42865),
            .in2(N__42795),
            .in3(N__43351),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47824),
            .ce(),
            .sr(N__47312));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_16_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_16_13_0 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_16_13_0  (
            .in0(N__44417),
            .in1(N__40646),
            .in2(_gnd_net_),
            .in3(N__40480),
            .lcout(\current_shift_inst.un38_control_input_cry_0_s0_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_16_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_16_14_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_16_14_0  (
            .in0(N__44426),
            .in1(N__45842),
            .in2(N__45176),
            .in3(N__43249),
            .lcout(\current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_16_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_16_14_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_16_14_1  (
            .in0(N__44422),
            .in1(N__45051),
            .in2(N__45767),
            .in3(N__40732),
            .lcout(\current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_16_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_16_14_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_16_14_2  (
            .in0(N__45061),
            .in1(N__44424),
            .in2(N__45548),
            .in3(N__40879),
            .lcout(\current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_16_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_16_14_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_16_14_3  (
            .in0(N__44421),
            .in1(N__45060),
            .in2(N__45622),
            .in3(N__40697),
            .lcout(\current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_16_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_16_14_4 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_16_14_4  (
            .in0(N__40733),
            .in1(N__45763),
            .in2(N__45177),
            .in3(N__44420),
            .lcout(\current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_16_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_16_14_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_16_14_5  (
            .in0(N__44423),
            .in1(N__45059),
            .in2(N__45623),
            .in3(N__40696),
            .lcout(\current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_16_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_16_14_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_16_14_6  (
            .in0(N__44427),
            .in1(N__45691),
            .in2(N__45178),
            .in3(N__40714),
            .lcout(\current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_16_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_16_14_7 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_16_14_7  (
            .in0(N__40715),
            .in1(N__45058),
            .in2(N__45692),
            .in3(N__44425),
            .lcout(\current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_15_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_15_0  (
            .in0(N__44081),
            .in1(N__45838),
            .in2(_gnd_net_),
            .in3(N__43248),
            .lcout(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_15_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_15_1  (
            .in0(N__45916),
            .in1(N__44080),
            .in2(_gnd_net_),
            .in3(N__40762),
            .lcout(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_16_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_16_15_2 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_16_15_2  (
            .in0(N__44534),
            .in1(N__45181),
            .in2(N__40880),
            .in3(N__45544),
            .lcout(\current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_15_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_15_3  (
            .in0(N__45984),
            .in1(N__44079),
            .in2(_gnd_net_),
            .in3(N__40792),
            .lcout(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_16_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_16_15_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_16_15_4  (
            .in0(N__44083),
            .in1(N__45682),
            .in2(_gnd_net_),
            .in3(N__40713),
            .lcout(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_15_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_15_5  (
            .in0(N__45610),
            .in1(N__44084),
            .in2(_gnd_net_),
            .in3(N__40695),
            .lcout(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_15_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_15_6  (
            .in0(N__44082),
            .in1(N__45757),
            .in2(_gnd_net_),
            .in3(N__40731),
            .lcout(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_15_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_15_7  (
            .in0(N__45543),
            .in1(N__44085),
            .in2(_gnd_net_),
            .in3(N__40875),
            .lcout(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_16_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_16_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_LC_16_16_0  (
            .in0(_gnd_net_),
            .in1(N__38582),
            .in2(N__38558),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_16_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_16_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_16_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_LC_16_16_1  (
            .in0(_gnd_net_),
            .in1(N__39035),
            .in2(N__43733),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_0 ),
            .carryout(\current_shift_inst.un10_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_16_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_16_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_LC_16_16_2  (
            .in0(_gnd_net_),
            .in1(N__38531),
            .in2(N__39064),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_1 ),
            .carryout(\current_shift_inst.un10_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_16_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_16_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_LC_16_16_3  (
            .in0(_gnd_net_),
            .in1(N__39039),
            .in2(N__38525),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_2 ),
            .carryout(\current_shift_inst.un10_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_16_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_16_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_LC_16_16_4  (
            .in0(_gnd_net_),
            .in1(N__38513),
            .in2(N__39065),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_3 ),
            .carryout(\current_shift_inst.un10_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_16_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_16_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_LC_16_16_5  (
            .in0(_gnd_net_),
            .in1(N__39043),
            .in2(N__38507),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_4 ),
            .carryout(\current_shift_inst.un10_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_16_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_16_16_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_LC_16_16_6  (
            .in0(_gnd_net_),
            .in1(N__38624),
            .in2(N__39066),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_5 ),
            .carryout(\current_shift_inst.un10_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_16_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_16_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_16_16_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_LC_16_16_7  (
            .in0(_gnd_net_),
            .in1(N__39047),
            .in2(N__38618),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_6 ),
            .carryout(\current_shift_inst.un10_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_16_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_16_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_LC_16_17_0  (
            .in0(_gnd_net_),
            .in1(N__39030),
            .in2(N__38609),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_17_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_16_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_16_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_LC_16_17_1  (
            .in0(_gnd_net_),
            .in1(N__39034),
            .in2(N__43856),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_8 ),
            .carryout(\current_shift_inst.un10_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_16_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_16_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_LC_16_17_2  (
            .in0(_gnd_net_),
            .in1(N__39027),
            .in2(N__43907),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_9 ),
            .carryout(\current_shift_inst.un10_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_16_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_16_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_LC_16_17_3  (
            .in0(_gnd_net_),
            .in1(N__39031),
            .in2(N__41177),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_10 ),
            .carryout(\current_shift_inst.un10_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_16_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_16_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_LC_16_17_4  (
            .in0(_gnd_net_),
            .in1(N__39028),
            .in2(N__41246),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_11 ),
            .carryout(\current_shift_inst.un10_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_16_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_16_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_LC_16_17_5  (
            .in0(_gnd_net_),
            .in1(N__39032),
            .in2(N__43568),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_12 ),
            .carryout(\current_shift_inst.un10_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_16_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_16_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_LC_16_17_6  (
            .in0(_gnd_net_),
            .in1(N__39029),
            .in2(N__38597),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_13 ),
            .carryout(\current_shift_inst.un10_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_16_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_16_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_LC_16_17_7  (
            .in0(_gnd_net_),
            .in1(N__39033),
            .in2(N__43214),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_14 ),
            .carryout(\current_shift_inst.un10_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_16_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_16_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_LC_16_18_0  (
            .in0(_gnd_net_),
            .in1(N__39011),
            .in2(N__43682),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_18_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_16_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_16_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_LC_16_18_1  (
            .in0(_gnd_net_),
            .in1(N__41027),
            .in2(N__39060),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_16 ),
            .carryout(\current_shift_inst.un10_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_16_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_16_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_LC_16_18_2  (
            .in0(_gnd_net_),
            .in1(N__39015),
            .in2(N__38684),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_17 ),
            .carryout(\current_shift_inst.un10_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_16_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_16_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_LC_16_18_3  (
            .in0(_gnd_net_),
            .in1(N__38672),
            .in2(N__39061),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_18 ),
            .carryout(\current_shift_inst.un10_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_16_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_16_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_LC_16_18_4  (
            .in0(_gnd_net_),
            .in1(N__39019),
            .in2(N__41048),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_19 ),
            .carryout(\current_shift_inst.un10_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_16_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_16_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_LC_16_18_5  (
            .in0(_gnd_net_),
            .in1(N__38657),
            .in2(N__39062),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_20 ),
            .carryout(\current_shift_inst.un10_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_16_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_16_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_LC_16_18_6  (
            .in0(_gnd_net_),
            .in1(N__39023),
            .in2(N__38645),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_21 ),
            .carryout(\current_shift_inst.un10_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_16_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_16_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_LC_16_18_7  (
            .in0(_gnd_net_),
            .in1(N__38633),
            .in2(N__39063),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_22 ),
            .carryout(\current_shift_inst.un10_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_16_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_16_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_LC_16_19_0  (
            .in0(_gnd_net_),
            .in1(N__38850),
            .in2(N__41234),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_19_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_16_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_16_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_LC_16_19_1  (
            .in0(_gnd_net_),
            .in1(N__44213),
            .in2(N__38922),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_24 ),
            .carryout(\current_shift_inst.un10_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_16_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_16_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_LC_16_19_2  (
            .in0(_gnd_net_),
            .in1(N__38854),
            .in2(N__41021),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_25 ),
            .carryout(\current_shift_inst.un10_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_16_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_16_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_LC_16_19_3  (
            .in0(_gnd_net_),
            .in1(N__40397),
            .in2(N__38923),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_26 ),
            .carryout(\current_shift_inst.un10_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_16_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_16_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_LC_16_19_4  (
            .in0(_gnd_net_),
            .in1(N__38858),
            .in2(N__41261),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_27 ),
            .carryout(\current_shift_inst.un10_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_16_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_16_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_LC_16_19_5  (
            .in0(_gnd_net_),
            .in1(N__41252),
            .in2(N__38924),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_28 ),
            .carryout(\current_shift_inst.un10_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_16_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_16_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_LC_16_19_6  (
            .in0(_gnd_net_),
            .in1(N__38862),
            .in2(N__44270),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_29 ),
            .carryout(\current_shift_inst.un10_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_16_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_16_19_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_16_19_7  (
            .in0(_gnd_net_),
            .in1(N__44611),
            .in2(_gnd_net_),
            .in3(N__38750),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_16_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_16_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_16_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39141),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_16_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_16_20_2 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_16_20_2  (
            .in0(N__44654),
            .in1(N__47915),
            .in2(N__44159),
            .in3(N__45257),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_20_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_20_5  (
            .in0(N__44652),
            .in1(N__46694),
            .in2(N__45287),
            .in3(N__40941),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.counter_0_LC_16_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_16_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_16_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_16_21_0  (
            .in0(N__39402),
            .in1(N__46008),
            .in2(_gnd_net_),
            .in3(N__39089),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_16_21_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__47778),
            .ce(N__39310),
            .sr(N__47361));
    defparam \current_shift_inst.timer_s1.counter_1_LC_16_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_16_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_16_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_16_21_1  (
            .in0(N__39406),
            .in1(N__45936),
            .in2(_gnd_net_),
            .in3(N__39086),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__47778),
            .ce(N__39310),
            .sr(N__47361));
    defparam \current_shift_inst.timer_s1.counter_2_LC_16_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_16_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_16_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_16_21_2  (
            .in0(N__39403),
            .in1(N__45861),
            .in2(_gnd_net_),
            .in3(N__39083),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__47778),
            .ce(N__39310),
            .sr(N__47361));
    defparam \current_shift_inst.timer_s1.counter_3_LC_16_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_16_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_16_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_16_21_3  (
            .in0(N__39407),
            .in1(N__45781),
            .in2(_gnd_net_),
            .in3(N__39080),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__47778),
            .ce(N__39310),
            .sr(N__47361));
    defparam \current_shift_inst.timer_s1.counter_4_LC_16_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_16_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_16_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_16_21_4  (
            .in0(N__39404),
            .in1(N__45708),
            .in2(_gnd_net_),
            .in3(N__39077),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__47778),
            .ce(N__39310),
            .sr(N__47361));
    defparam \current_shift_inst.timer_s1.counter_5_LC_16_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_16_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_16_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_16_21_5  (
            .in0(N__39408),
            .in1(N__45639),
            .in2(_gnd_net_),
            .in3(N__39074),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__47778),
            .ce(N__39310),
            .sr(N__47361));
    defparam \current_shift_inst.timer_s1.counter_6_LC_16_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_16_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_16_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_16_21_6  (
            .in0(N__39405),
            .in1(N__45564),
            .in2(_gnd_net_),
            .in3(N__39071),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__47778),
            .ce(N__39310),
            .sr(N__47361));
    defparam \current_shift_inst.timer_s1.counter_7_LC_16_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_16_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_16_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_16_21_7  (
            .in0(N__39409),
            .in1(N__45504),
            .in2(_gnd_net_),
            .in3(N__39170),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__47778),
            .ce(N__39310),
            .sr(N__47361));
    defparam \current_shift_inst.timer_s1.counter_8_LC_16_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_16_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_16_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_16_22_0  (
            .in0(N__39421),
            .in1(N__46512),
            .in2(_gnd_net_),
            .in3(N__39167),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_16_22_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__47775),
            .ce(N__39302),
            .sr(N__47370));
    defparam \current_shift_inst.timer_s1.counter_9_LC_16_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_16_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_16_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_16_22_1  (
            .in0(N__39431),
            .in1(N__46446),
            .in2(_gnd_net_),
            .in3(N__39164),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__47775),
            .ce(N__39302),
            .sr(N__47370));
    defparam \current_shift_inst.timer_s1.counter_10_LC_16_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_16_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_16_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_16_22_2  (
            .in0(N__39418),
            .in1(N__46383),
            .in2(_gnd_net_),
            .in3(N__39161),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__47775),
            .ce(N__39302),
            .sr(N__47370));
    defparam \current_shift_inst.timer_s1.counter_11_LC_16_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_16_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_16_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_16_22_3  (
            .in0(N__39428),
            .in1(N__46312),
            .in2(_gnd_net_),
            .in3(N__39158),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__47775),
            .ce(N__39302),
            .sr(N__47370));
    defparam \current_shift_inst.timer_s1.counter_12_LC_16_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_16_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_16_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_16_22_4  (
            .in0(N__39419),
            .in1(N__46257),
            .in2(_gnd_net_),
            .in3(N__39155),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__47775),
            .ce(N__39302),
            .sr(N__47370));
    defparam \current_shift_inst.timer_s1.counter_13_LC_16_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_16_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_16_22_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_16_22_5  (
            .in0(N__39429),
            .in1(N__46183),
            .in2(_gnd_net_),
            .in3(N__39152),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__47775),
            .ce(N__39302),
            .sr(N__47370));
    defparam \current_shift_inst.timer_s1.counter_14_LC_16_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_16_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_16_22_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_16_22_6  (
            .in0(N__39420),
            .in1(N__46126),
            .in2(_gnd_net_),
            .in3(N__39149),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__47775),
            .ce(N__39302),
            .sr(N__47370));
    defparam \current_shift_inst.timer_s1.counter_15_LC_16_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_16_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_16_22_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_16_22_7  (
            .in0(N__39430),
            .in1(N__46069),
            .in2(_gnd_net_),
            .in3(N__39146),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__47775),
            .ce(N__39302),
            .sr(N__47370));
    defparam \current_shift_inst.timer_s1.counter_16_LC_16_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_16_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_16_23_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_16_23_0  (
            .in0(N__39410),
            .in1(N__46968),
            .in2(_gnd_net_),
            .in3(N__39197),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_16_23_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__47770),
            .ce(N__39311),
            .sr(N__47377));
    defparam \current_shift_inst.timer_s1.counter_17_LC_16_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_16_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_16_23_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_16_23_1  (
            .in0(N__39422),
            .in1(N__46896),
            .in2(_gnd_net_),
            .in3(N__39194),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__47770),
            .ce(N__39311),
            .sr(N__47377));
    defparam \current_shift_inst.timer_s1.counter_18_LC_16_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_16_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_16_23_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_16_23_2  (
            .in0(N__39411),
            .in1(N__46839),
            .in2(_gnd_net_),
            .in3(N__39191),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__47770),
            .ce(N__39311),
            .sr(N__47377));
    defparam \current_shift_inst.timer_s1.counter_19_LC_16_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_16_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_16_23_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_16_23_3  (
            .in0(N__39423),
            .in1(N__46765),
            .in2(_gnd_net_),
            .in3(N__39188),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__47770),
            .ce(N__39311),
            .sr(N__47377));
    defparam \current_shift_inst.timer_s1.counter_20_LC_16_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_16_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_16_23_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_16_23_4  (
            .in0(N__39412),
            .in1(N__46710),
            .in2(_gnd_net_),
            .in3(N__39185),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__47770),
            .ce(N__39311),
            .sr(N__47377));
    defparam \current_shift_inst.timer_s1.counter_21_LC_16_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_16_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_16_23_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_16_23_5  (
            .in0(N__39424),
            .in1(N__46642),
            .in2(_gnd_net_),
            .in3(N__39182),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__47770),
            .ce(N__39311),
            .sr(N__47377));
    defparam \current_shift_inst.timer_s1.counter_22_LC_16_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_16_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_16_23_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_16_23_6  (
            .in0(N__39413),
            .in1(N__46579),
            .in2(_gnd_net_),
            .in3(N__39179),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__47770),
            .ce(N__39311),
            .sr(N__47377));
    defparam \current_shift_inst.timer_s1.counter_23_LC_16_23_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_16_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_16_23_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_16_23_7  (
            .in0(N__39425),
            .in1(N__48256),
            .in2(_gnd_net_),
            .in3(N__39176),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__47770),
            .ce(N__39311),
            .sr(N__47377));
    defparam \current_shift_inst.timer_s1.counter_24_LC_16_24_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_16_24_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_16_24_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_16_24_0  (
            .in0(N__39414),
            .in1(N__48189),
            .in2(_gnd_net_),
            .in3(N__39173),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_16_24_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__47766),
            .ce(N__39303),
            .sr(N__47385));
    defparam \current_shift_inst.timer_s1.counter_25_LC_16_24_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_16_24_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_16_24_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_16_24_1  (
            .in0(N__39426),
            .in1(N__48108),
            .in2(_gnd_net_),
            .in3(N__39443),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__47766),
            .ce(N__39303),
            .sr(N__47385));
    defparam \current_shift_inst.timer_s1.counter_26_LC_16_24_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_16_24_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_16_24_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_16_24_2  (
            .in0(N__39415),
            .in1(N__48024),
            .in2(_gnd_net_),
            .in3(N__39440),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__47766),
            .ce(N__39303),
            .sr(N__47385));
    defparam \current_shift_inst.timer_s1.counter_27_LC_16_24_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_16_24_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_16_24_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_16_24_3  (
            .in0(N__39427),
            .in1(N__47931),
            .in2(_gnd_net_),
            .in3(N__39437),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__47766),
            .ce(N__39303),
            .sr(N__47385));
    defparam \current_shift_inst.timer_s1.counter_28_LC_16_24_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_16_24_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_16_24_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_16_24_4  (
            .in0(N__39416),
            .in1(N__48043),
            .in2(_gnd_net_),
            .in3(N__39434),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__47766),
            .ce(N__39303),
            .sr(N__47385));
    defparam \current_shift_inst.timer_s1.counter_29_LC_16_24_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_16_24_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_16_24_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_16_24_5  (
            .in0(N__47956),
            .in1(N__39417),
            .in2(_gnd_net_),
            .in3(N__39314),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47766),
            .ce(N__39303),
            .sr(N__47385));
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_17_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_17_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_17_7_2 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_19_LC_17_7_2  (
            .in0(N__39761),
            .in1(N__42512),
            .in2(_gnd_net_),
            .in3(N__39275),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47867),
            .ce(N__42117),
            .sr(N__47282));
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_17_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_17_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_17_7_3 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_16_LC_17_7_3  (
            .in0(N__42515),
            .in1(N__41856),
            .in2(_gnd_net_),
            .in3(N__39763),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47867),
            .ce(N__42117),
            .sr(N__47282));
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_17_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_17_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_17_7_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_15_LC_17_7_4  (
            .in0(N__39762),
            .in1(N__39840),
            .in2(N__39815),
            .in3(N__42514),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47867),
            .ce(N__42117),
            .sr(N__47282));
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_17_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_17_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_17_7_5 .LUT_INIT=16'b0100000001000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_7_LC_17_7_5  (
            .in0(N__42516),
            .in1(N__42306),
            .in2(N__42626),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47867),
            .ce(N__42117),
            .sr(N__47282));
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_17_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_17_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_17_7_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_8_LC_17_7_6  (
            .in0(N__42304),
            .in1(N__42513),
            .in2(_gnd_net_),
            .in3(N__39521),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47867),
            .ce(N__42117),
            .sr(N__47282));
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_17_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_17_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_17_7_7 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_2_LC_17_7_7  (
            .in0(N__42517),
            .in1(N__42305),
            .in2(N__42239),
            .in3(N__42662),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47867),
            .ce(N__42117),
            .sr(N__47282));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5_1_LC_17_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5_1_LC_17_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5_1_LC_17_8_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5_1_LC_17_8_1  (
            .in0(N__39714),
            .in1(N__39587),
            .in2(N__39482),
            .in3(N__39550),
            .lcout(\phase_controller_inst1.stoper_tr.N_235 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_0_2_LC_17_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_0_2_LC_17_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_0_2_LC_17_8_3 .LUT_INIT=16'b0101110101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_0_2_LC_17_8_3  (
            .in0(N__39575),
            .in1(N__39478),
            .in2(N__42165),
            .in3(N__39549),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUKL2M1_6_LC_17_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUKL2M1_6_LC_17_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUKL2M1_6_LC_17_8_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUKL2M1_6_LC_17_8_4  (
            .in0(_gnd_net_),
            .in1(N__41498),
            .in2(_gnd_net_),
            .in3(N__39533),
            .lcout(elapsed_time_ns_1_RNIUKL2M1_0_6),
            .ltout(elapsed_time_ns_1_RNIUKL2M1_0_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_2_LC_17_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_2_LC_17_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_2_LC_17_8_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_2_LC_17_8_5  (
            .in0(N__39520),
            .in1(N__42614),
            .in2(N__39485),
            .in3(N__39862),
            .lcout(\phase_controller_inst1.stoper_tr.N_247 ),
            .ltout(\phase_controller_inst1.stoper_tr.N_247_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_6_LC_17_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_6_LC_17_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_6_LC_17_8_6 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_6_LC_17_8_6  (
            .in0(_gnd_net_),
            .in1(N__39807),
            .in2(N__39461),
            .in3(N__39713),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_17_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_17_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_17_8_7 .LUT_INIT=16'b0000001000000011;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_6_LC_17_8_7  (
            .in0(N__42690),
            .in1(N__42467),
            .in2(N__39458),
            .in3(N__42303),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47863),
            .ce(N__42098),
            .sr(N__47283));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_17_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_17_9_0 .LUT_INIT=16'b1110111111101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_17_9_0  (
            .in0(N__41585),
            .in1(N__40133),
            .in2(N__41811),
            .in3(N__39917),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_17_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_17_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_17_9_1 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_17_9_1  (
            .in0(N__40103),
            .in1(N__39800),
            .in2(N__41810),
            .in3(N__40056),
            .lcout(elapsed_time_ns_1_RNIUCHF91_0_15),
            .ltout(elapsed_time_ns_1_RNIUCHF91_0_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_9_LC_17_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_9_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_9_LC_17_9_2 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_9_LC_17_9_2  (
            .in0(_gnd_net_),
            .in1(N__39889),
            .in2(N__39953),
            .in3(N__39916),
            .lcout(\phase_controller_inst1.stoper_tr.N_251 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1OL2M1_9_LC_17_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1OL2M1_9_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1OL2M1_9_LC_17_9_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1OL2M1_9_LC_17_9_3  (
            .in0(_gnd_net_),
            .in1(N__39932),
            .in2(_gnd_net_),
            .in3(N__41499),
            .lcout(elapsed_time_ns_1_RNI1OL2M1_0_9),
            .ltout(elapsed_time_ns_1_RNI1OL2M1_0_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_6_LC_17_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_6_LC_17_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_6_LC_17_9_4 .LUT_INIT=16'b0011111100110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_6_LC_17_9_4  (
            .in0(_gnd_net_),
            .in1(N__39890),
            .in2(N__39866),
            .in3(N__39861),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.N_211_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_6_LC_17_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_6_LC_17_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_6_LC_17_9_5 .LUT_INIT=16'b0000000010111010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_6_LC_17_9_5  (
            .in0(N__39844),
            .in1(N__39801),
            .in2(N__39770),
            .in3(N__39715),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_0_6 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_1_LC_17_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_1_LC_17_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_1_LC_17_9_6 .LUT_INIT=16'b1111111100110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_1_LC_17_9_6  (
            .in0(_gnd_net_),
            .in1(N__41430),
            .in2(N__39635),
            .in3(N__42453),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_17_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_17_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_17_9_7 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_1_LC_17_9_7  (
            .in0(N__41431),
            .in1(N__42224),
            .in2(N__39632),
            .in3(N__41413),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47858),
            .ce(N__42118),
            .sr(N__47288));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_1_c_inv_LC_17_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_1_c_inv_LC_17_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_1_c_inv_LC_17_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_1_c_inv_LC_17_10_0  (
            .in0(_gnd_net_),
            .in1(N__39617),
            .in2(N__41393),
            .in3(N__42796),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_2_c_inv_LC_17_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_2_c_inv_LC_17_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_2_c_inv_LC_17_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_2_c_inv_LC_17_10_1  (
            .in0(_gnd_net_),
            .in1(N__42647),
            .in2(N__40229),
            .in3(N__42763),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_3_c_inv_LC_17_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_3_c_inv_LC_17_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_3_c_inv_LC_17_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_3_c_inv_LC_17_10_2  (
            .in0(_gnd_net_),
            .in1(N__40220),
            .in2(N__40214),
            .in3(N__42739),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_4_c_inv_LC_17_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_4_c_inv_LC_17_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_4_c_inv_LC_17_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_4_c_inv_LC_17_10_3  (
            .in0(_gnd_net_),
            .in1(N__42641),
            .in2(N__40205),
            .in3(N__42724),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_5_c_inv_LC_17_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_5_c_inv_LC_17_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_5_c_inv_LC_17_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_5_c_inv_LC_17_10_4  (
            .in0(_gnd_net_),
            .in1(N__40196),
            .in2(N__42635),
            .in3(N__42709),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_6_c_inv_LC_17_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_6_c_inv_LC_17_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_6_c_inv_LC_17_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_6_c_inv_LC_17_10_5  (
            .in0(_gnd_net_),
            .in1(N__40190),
            .in2(N__42671),
            .in3(N__43180),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_7_c_inv_LC_17_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_7_c_inv_LC_17_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_7_c_inv_LC_17_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_7_c_inv_LC_17_10_6  (
            .in0(_gnd_net_),
            .in1(N__42593),
            .in2(N__40181),
            .in3(N__43165),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_8_c_inv_LC_17_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_8_c_inv_LC_17_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_8_c_inv_LC_17_10_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_8_c_inv_LC_17_10_7  (
            .in0(N__43150),
            .in1(N__40172),
            .in2(N__40160),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_9_c_inv_LC_17_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_9_c_inv_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_9_c_inv_LC_17_11_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_9_c_inv_LC_17_11_0  (
            .in0(N__43135),
            .in1(N__40148),
            .in2(N__40142),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_10_c_inv_LC_17_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_10_c_inv_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_10_c_inv_LC_17_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_10_c_inv_LC_17_11_1  (
            .in0(_gnd_net_),
            .in1(N__40370),
            .in2(N__40385),
            .in3(N__43120),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_11_c_inv_LC_17_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_11_c_inv_LC_17_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_11_c_inv_LC_17_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_11_c_inv_LC_17_11_2  (
            .in0(_gnd_net_),
            .in1(N__40364),
            .in2(N__40352),
            .in3(N__43105),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_12_c_inv_LC_17_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_12_c_inv_LC_17_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_12_c_inv_LC_17_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_12_c_inv_LC_17_11_3  (
            .in0(_gnd_net_),
            .in1(N__40343),
            .in2(N__40331),
            .in3(N__43090),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_13_c_inv_LC_17_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_13_c_inv_LC_17_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_13_c_inv_LC_17_11_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_13_c_inv_LC_17_11_4  (
            .in0(N__43075),
            .in1(N__40322),
            .in2(N__40310),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_14_c_inv_LC_17_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_14_c_inv_LC_17_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_14_c_inv_LC_17_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_14_c_inv_LC_17_11_5  (
            .in0(_gnd_net_),
            .in1(N__40286),
            .in2(N__40301),
            .in3(N__43447),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_15_c_inv_LC_17_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_15_c_inv_LC_17_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_15_c_inv_LC_17_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_15_c_inv_LC_17_11_6  (
            .in0(_gnd_net_),
            .in1(N__40280),
            .in2(N__40274),
            .in3(N__43432),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_16_c_inv_LC_17_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_16_c_inv_LC_17_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_16_c_inv_LC_17_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_16_c_inv_LC_17_11_7  (
            .in0(_gnd_net_),
            .in1(N__40265),
            .in2(N__40259),
            .in3(N__43417),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_17_c_inv_LC_17_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_17_c_inv_LC_17_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_17_c_inv_LC_17_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_17_c_inv_LC_17_12_0  (
            .in0(_gnd_net_),
            .in1(N__40250),
            .in2(N__40238),
            .in3(N__43402),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_17_12_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_18_c_inv_LC_17_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_18_c_inv_LC_17_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_18_c_inv_LC_17_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_18_c_inv_LC_17_12_1  (
            .in0(_gnd_net_),
            .in1(N__40454),
            .in2(N__40442),
            .in3(N__43387),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_inv_LC_17_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_inv_LC_17_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_inv_LC_17_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_inv_LC_17_12_2  (
            .in0(_gnd_net_),
            .in1(N__40433),
            .in2(N__40421),
            .in3(N__43261),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_LUT4_0_LC_17_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_LUT4_0_LC_17_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_LUT4_0_LC_17_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_LUT4_0_LC_17_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40412),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNISF8I2_LC_17_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNISF8I2_LC_17_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNISF8I2_LC_17_12_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNISF8I2_LC_17_12_4  (
            .in0(_gnd_net_),
            .in1(N__42839),
            .in2(_gnd_net_),
            .in3(N__42864),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNISF8IZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_17_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_17_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_17_12_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_17_12_5  (
            .in0(N__43022),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42945),
            .lcout(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIM28A1_LC_17_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIM28A1_LC_17_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIM28A1_LC_17_12_7 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIM28A1_LC_17_12_7  (
            .in0(N__43021),
            .in1(N__42944),
            .in2(_gnd_net_),
            .in3(N__43054),
            .lcout(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_17_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_17_13_0 .LUT_INIT=16'b1100010111000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_17_13_0  (
            .in0(N__48086),
            .in1(N__41107),
            .in2(N__44480),
            .in3(N__45198),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_17_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_17_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_17_13_1 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_17_13_1  (
            .in0(N__41106),
            .in1(N__48085),
            .in2(_gnd_net_),
            .in3(N__44413),
            .lcout(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_17_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_17_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_17_13_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_17_13_2  (
            .in0(N__47019),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47825),
            .ce(N__47516),
            .sr(N__47313));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_17_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_17_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_17_13_3 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_17_13_3  (
            .in0(N__45199),
            .in1(N__44412),
            .in2(N__45989),
            .in3(N__40798),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_17_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_17_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_17_13_4 .LUT_INIT=16'b1010001110100011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_17_13_4  (
            .in0(N__40799),
            .in1(N__45985),
            .in2(N__44479),
            .in3(N__45200),
            .lcout(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_17_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_17_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_17_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_17_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40827),
            .lcout(\current_shift_inst.un4_control_input1_1 ),
            .ltout(\current_shift_inst.un4_control_input1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_17_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_17_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_17_13_7 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_17_13_7  (
            .in0(_gnd_net_),
            .in1(N__44408),
            .in2(N__40640),
            .in3(N__40479),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_17_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_17_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_17_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40612),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_17_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_17_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_17_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40547),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_17_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_17_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_17_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40475),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_17_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_17_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_17_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_17_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46019),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47819),
            .ce(N__47515),
            .sr(N__47316));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_17_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_17_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_17_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_17_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45836),
            .lcout(\current_shift_inst.un4_control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_17_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_17_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_17_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_17_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45756),
            .lcout(\current_shift_inst.un4_control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_15_0  (
            .in0(_gnd_net_),
            .in1(N__43817),
            .in2(N__40828),
            .in3(N__40826),
            .lcout(\current_shift_inst.un4_control_input1_2 ),
            .ltout(),
            .carryin(bfn_17_15_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_15_1  (
            .in0(_gnd_net_),
            .in1(N__43841),
            .in2(_gnd_net_),
            .in3(N__40781),
            .lcout(\current_shift_inst.un4_control_input1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_15_2  (
            .in0(_gnd_net_),
            .in1(N__43460),
            .in2(_gnd_net_),
            .in3(N__40751),
            .lcout(\current_shift_inst.un4_control_input1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_15_3  (
            .in0(_gnd_net_),
            .in1(N__40748),
            .in2(_gnd_net_),
            .in3(N__40742),
            .lcout(\current_shift_inst.un4_control_input1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_15_4  (
            .in0(_gnd_net_),
            .in1(N__40739),
            .in2(_gnd_net_),
            .in3(N__40718),
            .lcout(\current_shift_inst.un4_control_input1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_15_5  (
            .in0(_gnd_net_),
            .in1(N__44294),
            .in2(_gnd_net_),
            .in3(N__40700),
            .lcout(\current_shift_inst.un4_control_input1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_15_6  (
            .in0(_gnd_net_),
            .in1(N__43454),
            .in2(_gnd_net_),
            .in3(N__40682),
            .lcout(\current_shift_inst.un4_control_input1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_15_7  (
            .in0(_gnd_net_),
            .in1(N__44282),
            .in2(_gnd_net_),
            .in3(N__40862),
            .lcout(\current_shift_inst.un4_control_input1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_16_0  (
            .in0(_gnd_net_),
            .in1(N__45383),
            .in2(_gnd_net_),
            .in3(N__40859),
            .lcout(\current_shift_inst.un4_control_input1_10 ),
            .ltout(),
            .carryin(bfn_17_16_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_16_1  (
            .in0(_gnd_net_),
            .in1(N__41366),
            .in2(_gnd_net_),
            .in3(N__40856),
            .lcout(\current_shift_inst.un4_control_input1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_16_2  (
            .in0(_gnd_net_),
            .in1(N__44165),
            .in2(_gnd_net_),
            .in3(N__40853),
            .lcout(\current_shift_inst.un4_control_input1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_16_3  (
            .in0(_gnd_net_),
            .in1(N__41165),
            .in2(_gnd_net_),
            .in3(N__40850),
            .lcout(\current_shift_inst.un4_control_input1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_16_4  (
            .in0(_gnd_net_),
            .in1(N__44120),
            .in2(_gnd_net_),
            .in3(N__40847),
            .lcout(\current_shift_inst.un4_control_input1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_16_5  (
            .in0(_gnd_net_),
            .in1(N__41357),
            .in2(_gnd_net_),
            .in3(N__40844),
            .lcout(\current_shift_inst.un4_control_input1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_16_6  (
            .in0(_gnd_net_),
            .in1(N__41324),
            .in2(_gnd_net_),
            .in3(N__40841),
            .lcout(\current_shift_inst.un4_control_input1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_16_7  (
            .in0(_gnd_net_),
            .in1(N__41306),
            .in2(_gnd_net_),
            .in3(N__40838),
            .lcout(\current_shift_inst.un4_control_input1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_17_0  (
            .in0(_gnd_net_),
            .in1(N__45374),
            .in2(_gnd_net_),
            .in3(N__41009),
            .lcout(\current_shift_inst.un4_control_input1_18 ),
            .ltout(),
            .carryin(bfn_17_17_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_17_1  (
            .in0(_gnd_net_),
            .in1(N__41345),
            .in2(_gnd_net_),
            .in3(N__41006),
            .lcout(\current_shift_inst.un4_control_input1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_17_2  (
            .in0(_gnd_net_),
            .in1(N__41384),
            .in2(_gnd_net_),
            .in3(N__40976),
            .lcout(\current_shift_inst.un4_control_input1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_17_3  (
            .in0(_gnd_net_),
            .in1(N__43718),
            .in2(_gnd_net_),
            .in3(N__40973),
            .lcout(\current_shift_inst.un4_control_input1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_17_4  (
            .in0(_gnd_net_),
            .in1(N__41375),
            .in2(_gnd_net_),
            .in3(N__40946),
            .lcout(\current_shift_inst.un4_control_input1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_17_5  (
            .in0(_gnd_net_),
            .in1(N__45329),
            .in2(_gnd_net_),
            .in3(N__40916),
            .lcout(\current_shift_inst.un4_control_input1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_17_6  (
            .in0(_gnd_net_),
            .in1(N__41942),
            .in2(_gnd_net_),
            .in3(N__40889),
            .lcout(\current_shift_inst.un4_control_input1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_17_7  (
            .in0(_gnd_net_),
            .in1(N__41315),
            .in2(_gnd_net_),
            .in3(N__40886),
            .lcout(\current_shift_inst.un4_control_input1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_18_0  (
            .in0(_gnd_net_),
            .in1(N__41951),
            .in2(_gnd_net_),
            .in3(N__40883),
            .lcout(\current_shift_inst.un4_control_input1_26 ),
            .ltout(),
            .carryin(bfn_17_18_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_18_1  (
            .in0(_gnd_net_),
            .in1(N__41333),
            .in2(_gnd_net_),
            .in3(N__41114),
            .lcout(\current_shift_inst.un4_control_input1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_18_2  (
            .in0(_gnd_net_),
            .in1(N__41915),
            .in2(_gnd_net_),
            .in3(N__41087),
            .lcout(\current_shift_inst.un4_control_input1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_18_3  (
            .in0(_gnd_net_),
            .in1(N__41933),
            .in2(_gnd_net_),
            .in3(N__41084),
            .lcout(\current_shift_inst.un4_control_input1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_18_4  (
            .in0(_gnd_net_),
            .in1(N__41924),
            .in2(_gnd_net_),
            .in3(N__41081),
            .lcout(\current_shift_inst.un4_control_input1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41078),
            .lcout(\current_shift_inst.un4_control_input1_31_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_17_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_17_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_17_18_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_17_18_6  (
            .in0(N__46805),
            .in1(N__44092),
            .in2(_gnd_net_),
            .in3(N__41064),
            .lcout(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_17_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_17_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_17_18_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_17_18_7  (
            .in0(N__44609),
            .in1(N__46945),
            .in2(N__45253),
            .in3(N__41148),
            .lcout(\current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_19_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_19_0  (
            .in0(N__44088),
            .in1(N__46046),
            .in2(_gnd_net_),
            .in3(N__43650),
            .lcout(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_17_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_17_19_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_17_19_1  (
            .in0(N__44592),
            .in1(_gnd_net_),
            .in2(N__48159),
            .in3(N__44193),
            .lcout(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_17_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_17_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_17_19_2 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_17_19_2  (
            .in0(N__45258),
            .in1(N__44591),
            .in2(N__45428),
            .in3(N__46292),
            .lcout(\current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_19_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_19_3  (
            .in0(N__44593),
            .in1(N__47991),
            .in2(_gnd_net_),
            .in3(N__41272),
            .lcout(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_17_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_17_19_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_17_19_4  (
            .in0(N__47907),
            .in1(N__44594),
            .in2(_gnd_net_),
            .in3(N__44145),
            .lcout(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_19_5 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_19_5  (
            .in0(N__43611),
            .in1(N__44087),
            .in2(_gnd_net_),
            .in3(N__46344),
            .lcout(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_17_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_17_19_6 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_17_19_6  (
            .in0(_gnd_net_),
            .in1(N__46558),
            .in2(N__44098),
            .in3(N__45368),
            .lcout(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_17_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_17_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_17_19_7 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_17_19_7  (
            .in0(N__44590),
            .in1(N__45259),
            .in2(N__43886),
            .in3(N__45477),
            .lcout(\current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_17_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_17_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_17_20_0 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_17_20_0  (
            .in0(N__41208),
            .in1(N__44086),
            .in2(_gnd_net_),
            .in3(N__46412),
            .lcout(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46343),
            .lcout(\current_shift_inst.un4_control_input_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_17_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_17_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_17_20_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_17_20_3  (
            .in0(N__44610),
            .in1(N__46935),
            .in2(N__45288),
            .in3(N__41155),
            .lcout(\current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_20_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_20_4  (
            .in0(N__46858),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_17_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_17_20_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_17_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46735),
            .lcout(\current_shift_inst.un4_control_input_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_17_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_17_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_17_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46473),
            .lcout(\current_shift_inst.un4_control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_17_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_17_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_17_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46215),
            .lcout(\current_shift_inst.un4_control_input_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_21_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46929),
            .lcout(\current_shift_inst.un4_control_input_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48140),
            .lcout(\current_shift_inst.un4_control_input_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_17_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_17_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_17_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46154),
            .lcout(\current_shift_inst.un4_control_input_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_21_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46542),
            .lcout(\current_shift_inst.un4_control_input_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_17_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_17_21_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_17_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46095),
            .lcout(\current_shift_inst.un4_control_input_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_21_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48219),
            .lcout(\current_shift_inst.un4_control_input_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_21_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46605),
            .lcout(\current_shift_inst.un4_control_input_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_21_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47981),
            .lcout(\current_shift_inst.un4_control_input_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_22_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47897),
            .lcout(\current_shift_inst.un4_control_input_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_17_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_17_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_17_22_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_17_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48066),
            .lcout(\current_shift_inst.un4_control_input_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_18_7_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_18_7_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_18_7_7 .LUT_INIT=16'b1101111111001110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_18_7_7  (
            .in0(N__41805),
            .in1(N__41587),
            .in2(N__41906),
            .in3(N__41432),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_18_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_18_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_18_8_1 .LUT_INIT=16'b1111111110101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_18_8_1  (
            .in0(N__41885),
            .in1(N__41861),
            .in2(N__41824),
            .in3(N__41588),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPFL2M1_1_LC_18_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPFL2M1_1_LC_18_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPFL2M1_1_LC_18_9_1 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPFL2M1_1_LC_18_9_1  (
            .in0(N__41503),
            .in1(N__41441),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(elapsed_time_ns_1_RNIPFL2M1_0_1),
            .ltout(elapsed_time_ns_1_RNIPFL2M1_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_18_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_18_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_18_9_2 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_1_LC_18_9_2  (
            .in0(N__42220),
            .in1(N__41414),
            .in2(N__41402),
            .in3(N__41399),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47864),
            .ce(N__43368),
            .sr(N__47284));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_18_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_18_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_18_9_3 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_LC_18_9_3  (
            .in0(N__42534),
            .in1(N__42296),
            .in2(N__42240),
            .in3(N__42691),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47864),
            .ce(N__43368),
            .sr(N__47284));
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_18_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_18_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_18_9_4 .LUT_INIT=16'b0000000000110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_2_LC_18_9_4  (
            .in0(N__42221),
            .in1(N__42661),
            .in2(N__42307),
            .in3(N__42536),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47864),
            .ce(N__43368),
            .sr(N__47284));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_18_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_18_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_18_9_5 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_LC_18_9_5  (
            .in0(N__42533),
            .in1(N__42295),
            .in2(N__42586),
            .in3(N__42223),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47864),
            .ce(N__43368),
            .sr(N__47284));
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_18_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_18_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_18_9_6 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_5_LC_18_9_6  (
            .in0(N__42222),
            .in1(N__42535),
            .in2(N__42308),
            .in3(N__42377),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47864),
            .ce(N__43368),
            .sr(N__47284));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_18_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_18_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_18_9_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_LC_18_9_7  (
            .in0(N__42532),
            .in1(N__42294),
            .in2(_gnd_net_),
            .in3(N__42625),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47864),
            .ce(N__43368),
            .sr(N__47284));
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_18_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_18_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_18_10_0 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_4_LC_18_10_0  (
            .in0(N__42530),
            .in1(N__42232),
            .in2(N__42587),
            .in3(N__42293),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47859),
            .ce(N__42115),
            .sr(N__47289));
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_18_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_18_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_18_10_1 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_5_LC_18_10_1  (
            .in0(N__42291),
            .in1(N__42531),
            .in2(N__42241),
            .in3(N__42373),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47859),
            .ce(N__42115),
            .sr(N__47289));
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_18_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_18_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_18_10_2 .LUT_INIT=16'b1111111010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_3_LC_18_10_2  (
            .in0(N__42331),
            .in1(N__42292),
            .in2(N__42242),
            .in3(N__42170),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47859),
            .ce(N__42115),
            .sr(N__47289));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIM28A1_0_LC_18_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIM28A1_0_LC_18_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIM28A1_0_LC_18_10_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIM28A1_0_LC_18_10_3  (
            .in0(N__43061),
            .in1(N__42971),
            .in2(_gnd_net_),
            .in3(N__43030),
            .lcout(\phase_controller_inst1.stoper_tr.running_1_sqmuxa ),
            .ltout(\phase_controller_inst1.stoper_tr.running_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_18_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_18_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_18_10_4 .LUT_INIT=16'b0000111100000111;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_18_10_4  (
            .in0(N__43031),
            .in1(N__42979),
            .in2(N__42914),
            .in3(N__42911),
            .lcout(\phase_controller_inst1.stoper_tr.un1_start_latched2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_18_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_18_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_18_10_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_18_10_7  (
            .in0(N__42866),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42844),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_18_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_18_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_18_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_18_11_0  (
            .in0(_gnd_net_),
            .in1(N__42806),
            .in2(N__42800),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_11_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_18_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_18_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_18_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_18_11_1  (
            .in0(N__43333),
            .in1(N__42764),
            .in2(_gnd_net_),
            .in3(N__42752),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__47846),
            .ce(),
            .sr(N__47295));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_18_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_18_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_18_11_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_18_11_2  (
            .in0(N__43337),
            .in1(N__42749),
            .in2(N__42743),
            .in3(N__42728),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__47846),
            .ce(),
            .sr(N__47295));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_18_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_18_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_18_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_18_11_3  (
            .in0(N__43334),
            .in1(N__42725),
            .in2(_gnd_net_),
            .in3(N__42713),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__47846),
            .ce(),
            .sr(N__47295));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_18_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_18_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_18_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_18_11_4  (
            .in0(N__43338),
            .in1(N__42710),
            .in2(_gnd_net_),
            .in3(N__42698),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__47846),
            .ce(),
            .sr(N__47295));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_18_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_18_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_18_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_18_11_5  (
            .in0(N__43335),
            .in1(N__43181),
            .in2(_gnd_net_),
            .in3(N__43169),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__47846),
            .ce(),
            .sr(N__47295));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_18_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_18_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_18_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_18_11_6  (
            .in0(N__43339),
            .in1(N__43166),
            .in2(_gnd_net_),
            .in3(N__43154),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__47846),
            .ce(),
            .sr(N__47295));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_18_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_18_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_18_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_18_11_7  (
            .in0(N__43336),
            .in1(N__43151),
            .in2(_gnd_net_),
            .in3(N__43139),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__47846),
            .ce(),
            .sr(N__47295));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_18_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_18_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_18_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_18_12_0  (
            .in0(N__43372),
            .in1(N__43136),
            .in2(_gnd_net_),
            .in3(N__43124),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_18_12_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__47838),
            .ce(),
            .sr(N__47303));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_18_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_18_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_18_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_18_12_1  (
            .in0(N__43326),
            .in1(N__43121),
            .in2(_gnd_net_),
            .in3(N__43109),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__47838),
            .ce(),
            .sr(N__47303));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_18_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_18_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_18_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_18_12_2  (
            .in0(N__43369),
            .in1(N__43106),
            .in2(_gnd_net_),
            .in3(N__43094),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__47838),
            .ce(),
            .sr(N__47303));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_18_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_18_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_18_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_18_12_3  (
            .in0(N__43327),
            .in1(N__43091),
            .in2(_gnd_net_),
            .in3(N__43079),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__47838),
            .ce(),
            .sr(N__47303));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_18_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_18_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_18_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_18_12_4  (
            .in0(N__43370),
            .in1(N__43076),
            .in2(_gnd_net_),
            .in3(N__43064),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__47838),
            .ce(),
            .sr(N__47303));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_18_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_18_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_18_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_18_12_5  (
            .in0(N__43328),
            .in1(N__43448),
            .in2(_gnd_net_),
            .in3(N__43436),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__47838),
            .ce(),
            .sr(N__47303));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_18_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_18_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_18_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_18_12_6  (
            .in0(N__43371),
            .in1(N__43433),
            .in2(_gnd_net_),
            .in3(N__43421),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__47838),
            .ce(),
            .sr(N__47303));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_18_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_18_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_18_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_18_12_7  (
            .in0(N__43329),
            .in1(N__43418),
            .in2(_gnd_net_),
            .in3(N__43406),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__47838),
            .ce(),
            .sr(N__47303));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_18_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_18_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_18_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_18_13_0  (
            .in0(N__43330),
            .in1(N__43403),
            .in2(_gnd_net_),
            .in3(N__43391),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_18_13_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__47830),
            .ce(),
            .sr(N__47307));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_18_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_18_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_18_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_18_13_1  (
            .in0(N__43332),
            .in1(N__43388),
            .in2(_gnd_net_),
            .in3(N__43376),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__47830),
            .ce(),
            .sr(N__47307));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_18_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_18_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_18_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_18_13_2  (
            .in0(N__43331),
            .in1(N__43262),
            .in2(_gnd_net_),
            .in3(N__43265),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47830),
            .ce(),
            .sr(N__47307));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_18_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_18_14_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_18_14_1  (
            .in0(N__44418),
            .in1(N__45837),
            .in2(N__45180),
            .in3(N__43250),
            .lcout(\current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_18_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_18_14_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_18_14_2  (
            .in0(N__44075),
            .in1(N__46164),
            .in2(_gnd_net_),
            .in3(N__43497),
            .lcout(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_18_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_18_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_18_14_3 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_18_14_3  (
            .in0(N__45065),
            .in1(N__44456),
            .in2(N__43708),
            .in3(N__46111),
            .lcout(\current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_18_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_18_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_18_14_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_18_14_4  (
            .in0(N__46812),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_18_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_18_14_5 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_18_14_5  (
            .in0(N__43701),
            .in1(N__44076),
            .in2(_gnd_net_),
            .in3(N__46110),
            .lcout(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_18_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_18_14_6 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_18_14_6  (
            .in0(N__44457),
            .in1(N__46055),
            .in2(N__43663),
            .in3(N__45066),
            .lcout(\current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_18_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_18_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_18_14_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_18_14_7  (
            .in0(N__44419),
            .in1(N__46351),
            .in2(N__45179),
            .in3(N__43612),
            .lcout(\current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_18_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_18_15_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_18_15_0  (
            .in0(N__46298),
            .in1(N__44094),
            .in2(_gnd_net_),
            .in3(N__45417),
            .lcout(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_18_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_18_15_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_18_15_1  (
            .in0(N__46227),
            .in1(N__44477),
            .in2(N__45264),
            .in3(N__43545),
            .lcout(\current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_18_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_18_15_2 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_18_15_2  (
            .in0(N__44478),
            .in1(N__45215),
            .in2(N__43508),
            .in3(N__46165),
            .lcout(\current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_18_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_18_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_18_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_18_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45899),
            .lcout(\current_shift_inst.un4_control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_18_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_18_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_18_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_18_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45603),
            .lcout(\current_shift_inst.un4_control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_18_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_18_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_18_15_5 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_18_15_5  (
            .in0(N__45211),
            .in1(N__44476),
            .in2(N__46490),
            .in3(N__43927),
            .lcout(\current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_18_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_18_15_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_18_15_6  (
            .in0(N__45478),
            .in1(N__44093),
            .in2(_gnd_net_),
            .in3(N__43872),
            .lcout(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_18_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_18_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_18_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_18_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45975),
            .lcout(\current_shift_inst.un4_control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_18_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_18_16_0 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_18_16_0  (
            .in0(N__44463),
            .in1(N__43759),
            .in2(N__43811),
            .in3(N__43747),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45950),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47815),
            .ce(N__47514),
            .sr(N__47322));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43745),
            .lcout(\current_shift_inst.un4_control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_16_3 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_16_3  (
            .in0(N__43748),
            .in1(N__44464),
            .in2(N__43763),
            .in3(N__43810),
            .lcout(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_18_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_18_16_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_18_16_4  (
            .in0(N__44078),
            .in1(N__43758),
            .in2(_gnd_net_),
            .in3(N__43746),
            .lcout(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_18_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_18_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_18_16_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_18_16_5  (
            .in0(_gnd_net_),
            .in1(N__44465),
            .in2(_gnd_net_),
            .in3(N__44254),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_18_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_18_16_6 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_18_16_6  (
            .in0(N__44255),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44579),
            .lcout(\current_shift_inst.un4_control_input_0_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_18_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_18_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_18_16_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_18_16_7  (
            .in0(N__44578),
            .in1(N__48237),
            .in2(_gnd_net_),
            .in3(N__45316),
            .lcout(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_18_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_18_17_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_18_17_0  (
            .in0(N__45267),
            .in1(N__44576),
            .in2(N__48166),
            .in3(N__44197),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46419),
            .lcout(\current_shift_inst.un4_control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_18_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_18_17_2 .LUT_INIT=16'b1111000000110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_18_17_2  (
            .in0(N__45265),
            .in1(N__47914),
            .in2(N__44155),
            .in3(N__44577),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_18_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_18_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_18_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46293),
            .lcout(\current_shift_inst.un4_control_input_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_18_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_18_17_4 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_18_17_4  (
            .in0(N__46483),
            .in1(N__43931),
            .in2(N__45289),
            .in3(N__44573),
            .lcout(\current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_18_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_18_17_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_18_17_5  (
            .in0(N__44099),
            .in1(N__46482),
            .in2(_gnd_net_),
            .in3(N__43923),
            .lcout(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_18_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_18_17_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_18_17_6  (
            .in0(N__45266),
            .in1(N__44575),
            .in2(N__46565),
            .in3(N__45366),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_18_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_18_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_18_17_7 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_18_17_7  (
            .in0(N__44574),
            .in1(N__45271),
            .in2(N__45424),
            .in3(N__46294),
            .lcout(\current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_18_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_18_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_18_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45470),
            .lcout(\current_shift_inst.un4_control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_18_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_18_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_18_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46050),
            .lcout(\current_shift_inst.un4_control_input_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_18_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_18_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_18_18_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_18_18_3  (
            .in0(N__44644),
            .in1(N__46557),
            .in2(N__45290),
            .in3(N__45367),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_18_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_18_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_18_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46682),
            .lcout(\current_shift_inst.un4_control_input_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_18_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_18_18_5 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_18_18_5  (
            .in0(N__48238),
            .in1(N__45315),
            .in2(N__45291),
            .in3(N__44645),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_18_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_18_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_18_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_18_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45669),
            .lcout(\current_shift_inst.un4_control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_18_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_18_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_18_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_18_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45529),
            .lcout(\current_shift_inst.un4_control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_18_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_18_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_18_19_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_18_19_0  (
            .in0(_gnd_net_),
            .in1(N__46018),
            .in2(N__45868),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_18_19_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__47797),
            .ce(N__47513),
            .sr(N__47332));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_18_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_18_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_18_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_18_19_1  (
            .in0(_gnd_net_),
            .in1(N__45946),
            .in2(N__45793),
            .in3(N__45872),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__47797),
            .ce(N__47513),
            .sr(N__47332));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_18_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_18_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_18_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_18_19_2  (
            .in0(_gnd_net_),
            .in1(N__45715),
            .in2(N__45869),
            .in3(N__45797),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__47797),
            .ce(N__47513),
            .sr(N__47332));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_18_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_18_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_18_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_18_19_3  (
            .in0(_gnd_net_),
            .in1(N__45646),
            .in2(N__45794),
            .in3(N__45722),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__47797),
            .ce(N__47513),
            .sr(N__47332));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_18_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_18_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_18_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_18_19_4  (
            .in0(_gnd_net_),
            .in1(N__45571),
            .in2(N__45719),
            .in3(N__45653),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__47797),
            .ce(N__47513),
            .sr(N__47332));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_18_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_18_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_18_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_18_19_5  (
            .in0(_gnd_net_),
            .in1(N__45511),
            .in2(N__45650),
            .in3(N__45578),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__47797),
            .ce(N__47513),
            .sr(N__47332));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_18_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_18_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_18_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_18_19_6  (
            .in0(_gnd_net_),
            .in1(N__46519),
            .in2(N__45575),
            .in3(N__45518),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__47797),
            .ce(N__47513),
            .sr(N__47332));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_18_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_18_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_18_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_18_19_7  (
            .in0(_gnd_net_),
            .in1(N__46453),
            .in2(N__45515),
            .in3(N__45449),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__47797),
            .ce(N__47513),
            .sr(N__47332));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_18_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_18_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_18_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_18_20_0  (
            .in0(_gnd_net_),
            .in1(N__46384),
            .in2(N__46523),
            .in3(N__46460),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_18_20_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__47792),
            .ce(N__47512),
            .sr(N__47334));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_18_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_18_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_18_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_18_20_1  (
            .in0(_gnd_net_),
            .in1(N__46318),
            .in2(N__46457),
            .in3(N__46391),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__47792),
            .ce(N__47512),
            .sr(N__47334));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_18_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_18_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_18_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_18_20_2  (
            .in0(_gnd_net_),
            .in1(N__46264),
            .in2(N__46388),
            .in3(N__46322),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__47792),
            .ce(N__47512),
            .sr(N__47334));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_18_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_18_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_18_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_18_20_3  (
            .in0(_gnd_net_),
            .in1(N__46319),
            .in2(N__46195),
            .in3(N__46271),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__47792),
            .ce(N__47512),
            .sr(N__47334));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_18_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_18_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_18_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_18_20_4  (
            .in0(_gnd_net_),
            .in1(N__46132),
            .in2(N__46268),
            .in3(N__46199),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__47792),
            .ce(N__47512),
            .sr(N__47334));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_18_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_18_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_18_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_18_20_5  (
            .in0(_gnd_net_),
            .in1(N__46075),
            .in2(N__46196),
            .in3(N__46136),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__47792),
            .ce(N__47512),
            .sr(N__47334));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_18_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_18_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_18_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_18_20_6  (
            .in0(_gnd_net_),
            .in1(N__46133),
            .in2(N__46981),
            .in3(N__46079),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__47792),
            .ce(N__47512),
            .sr(N__47334));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_18_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_18_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_18_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_18_20_7  (
            .in0(_gnd_net_),
            .in1(N__46076),
            .in2(N__46909),
            .in3(N__46022),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__47792),
            .ce(N__47512),
            .sr(N__47334));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_18_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_18_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_18_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_18_21_0  (
            .in0(_gnd_net_),
            .in1(N__46840),
            .in2(N__46982),
            .in3(N__46913),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_18_21_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__47787),
            .ce(N__47511),
            .sr(N__47340));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_18_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_18_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_18_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_18_21_1  (
            .in0(_gnd_net_),
            .in1(N__46771),
            .in2(N__46910),
            .in3(N__46847),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__47787),
            .ce(N__47511),
            .sr(N__47340));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_18_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_18_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_18_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_18_21_2  (
            .in0(_gnd_net_),
            .in1(N__46717),
            .in2(N__46844),
            .in3(N__46775),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__47787),
            .ce(N__47511),
            .sr(N__47340));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_18_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_18_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_18_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_18_21_3  (
            .in0(_gnd_net_),
            .in1(N__46772),
            .in2(N__46654),
            .in3(N__46724),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__47787),
            .ce(N__47511),
            .sr(N__47340));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_18_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_18_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_18_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_18_21_4  (
            .in0(_gnd_net_),
            .in1(N__46585),
            .in2(N__46721),
            .in3(N__46658),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__47787),
            .ce(N__47511),
            .sr(N__47340));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_18_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_18_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_18_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_18_21_5  (
            .in0(_gnd_net_),
            .in1(N__48262),
            .in2(N__46655),
            .in3(N__46589),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__47787),
            .ce(N__47511),
            .sr(N__47340));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_18_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_18_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_18_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_18_21_6  (
            .in0(_gnd_net_),
            .in1(N__46586),
            .in2(N__48202),
            .in3(N__46526),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__47787),
            .ce(N__47511),
            .sr(N__47340));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_18_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_18_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_18_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_18_21_7  (
            .in0(_gnd_net_),
            .in1(N__48263),
            .in2(N__48121),
            .in3(N__48206),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__47787),
            .ce(N__47511),
            .sr(N__47340));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_18_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_18_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_18_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_18_22_0  (
            .in0(_gnd_net_),
            .in1(N__48025),
            .in2(N__48203),
            .in3(N__48125),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_18_22_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__47783),
            .ce(N__47510),
            .sr(N__47351));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_18_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_18_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_18_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_18_22_1  (
            .in0(_gnd_net_),
            .in1(N__47938),
            .in2(N__48122),
            .in3(N__48050),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__47783),
            .ce(N__47510),
            .sr(N__47351));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_18_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_18_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_18_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_18_22_2  (
            .in0(_gnd_net_),
            .in1(N__48047),
            .in2(N__48029),
            .in3(N__47963),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__47783),
            .ce(N__47510),
            .sr(N__47351));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_18_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_18_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_18_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_18_22_3  (
            .in0(_gnd_net_),
            .in1(N__47960),
            .in2(N__47942),
            .in3(N__47879),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__47783),
            .ce(N__47510),
            .sr(N__47351));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_18_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_18_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_18_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_18_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47024),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // MAIN
