// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Feb 27 2025 18:59:42

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    rgb_g,
    T01,
    start_stop,
    s2_phy,
    T23,
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    clock_output,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    T45,
    T12,
    s4_phy,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    output rgb_g;
    output T01;
    input start_stop;
    output s2_phy;
    output T23;
    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    output clock_output;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output T45;
    output T12;
    output s4_phy;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__49535;
    wire N__49534;
    wire N__49533;
    wire N__49524;
    wire N__49523;
    wire N__49522;
    wire N__49515;
    wire N__49514;
    wire N__49513;
    wire N__49506;
    wire N__49505;
    wire N__49504;
    wire N__49497;
    wire N__49496;
    wire N__49495;
    wire N__49488;
    wire N__49487;
    wire N__49486;
    wire N__49479;
    wire N__49478;
    wire N__49477;
    wire N__49470;
    wire N__49469;
    wire N__49468;
    wire N__49461;
    wire N__49460;
    wire N__49459;
    wire N__49452;
    wire N__49451;
    wire N__49450;
    wire N__49443;
    wire N__49442;
    wire N__49441;
    wire N__49434;
    wire N__49433;
    wire N__49432;
    wire N__49425;
    wire N__49424;
    wire N__49423;
    wire N__49416;
    wire N__49415;
    wire N__49414;
    wire N__49407;
    wire N__49406;
    wire N__49405;
    wire N__49398;
    wire N__49397;
    wire N__49396;
    wire N__49389;
    wire N__49388;
    wire N__49387;
    wire N__49380;
    wire N__49379;
    wire N__49378;
    wire N__49361;
    wire N__49358;
    wire N__49355;
    wire N__49352;
    wire N__49349;
    wire N__49346;
    wire N__49345;
    wire N__49342;
    wire N__49339;
    wire N__49336;
    wire N__49331;
    wire N__49330;
    wire N__49329;
    wire N__49322;
    wire N__49319;
    wire N__49318;
    wire N__49317;
    wire N__49316;
    wire N__49313;
    wire N__49304;
    wire N__49301;
    wire N__49300;
    wire N__49297;
    wire N__49294;
    wire N__49289;
    wire N__49288;
    wire N__49285;
    wire N__49282;
    wire N__49281;
    wire N__49276;
    wire N__49273;
    wire N__49268;
    wire N__49265;
    wire N__49262;
    wire N__49259;
    wire N__49256;
    wire N__49253;
    wire N__49252;
    wire N__49249;
    wire N__49246;
    wire N__49243;
    wire N__49238;
    wire N__49235;
    wire N__49234;
    wire N__49233;
    wire N__49230;
    wire N__49225;
    wire N__49222;
    wire N__49219;
    wire N__49214;
    wire N__49211;
    wire N__49208;
    wire N__49207;
    wire N__49204;
    wire N__49203;
    wire N__49200;
    wire N__49195;
    wire N__49192;
    wire N__49187;
    wire N__49184;
    wire N__49181;
    wire N__49178;
    wire N__49177;
    wire N__49176;
    wire N__49173;
    wire N__49168;
    wire N__49163;
    wire N__49160;
    wire N__49159;
    wire N__49158;
    wire N__49153;
    wire N__49150;
    wire N__49145;
    wire N__49142;
    wire N__49139;
    wire N__49136;
    wire N__49133;
    wire N__49130;
    wire N__49127;
    wire N__49126;
    wire N__49125;
    wire N__49122;
    wire N__49117;
    wire N__49116;
    wire N__49111;
    wire N__49108;
    wire N__49103;
    wire N__49100;
    wire N__49097;
    wire N__49094;
    wire N__49091;
    wire N__49088;
    wire N__49087;
    wire N__49084;
    wire N__49083;
    wire N__49080;
    wire N__49077;
    wire N__49074;
    wire N__49067;
    wire N__49066;
    wire N__49065;
    wire N__49064;
    wire N__49063;
    wire N__49062;
    wire N__49059;
    wire N__49056;
    wire N__49055;
    wire N__49054;
    wire N__49051;
    wire N__49050;
    wire N__49045;
    wire N__49042;
    wire N__49039;
    wire N__49036;
    wire N__49031;
    wire N__49026;
    wire N__49021;
    wire N__49018;
    wire N__49015;
    wire N__49010;
    wire N__49007;
    wire N__49004;
    wire N__49001;
    wire N__48998;
    wire N__48995;
    wire N__48990;
    wire N__48987;
    wire N__48980;
    wire N__48979;
    wire N__48978;
    wire N__48977;
    wire N__48976;
    wire N__48973;
    wire N__48968;
    wire N__48963;
    wire N__48962;
    wire N__48961;
    wire N__48960;
    wire N__48959;
    wire N__48958;
    wire N__48953;
    wire N__48950;
    wire N__48947;
    wire N__48940;
    wire N__48937;
    wire N__48930;
    wire N__48927;
    wire N__48924;
    wire N__48919;
    wire N__48916;
    wire N__48913;
    wire N__48908;
    wire N__48907;
    wire N__48904;
    wire N__48901;
    wire N__48900;
    wire N__48897;
    wire N__48894;
    wire N__48891;
    wire N__48888;
    wire N__48883;
    wire N__48878;
    wire N__48875;
    wire N__48872;
    wire N__48871;
    wire N__48870;
    wire N__48869;
    wire N__48868;
    wire N__48867;
    wire N__48864;
    wire N__48859;
    wire N__48852;
    wire N__48851;
    wire N__48846;
    wire N__48843;
    wire N__48840;
    wire N__48833;
    wire N__48830;
    wire N__48827;
    wire N__48826;
    wire N__48825;
    wire N__48820;
    wire N__48817;
    wire N__48812;
    wire N__48809;
    wire N__48808;
    wire N__48807;
    wire N__48806;
    wire N__48805;
    wire N__48804;
    wire N__48803;
    wire N__48802;
    wire N__48801;
    wire N__48800;
    wire N__48799;
    wire N__48798;
    wire N__48797;
    wire N__48796;
    wire N__48795;
    wire N__48794;
    wire N__48793;
    wire N__48792;
    wire N__48791;
    wire N__48790;
    wire N__48789;
    wire N__48788;
    wire N__48787;
    wire N__48786;
    wire N__48785;
    wire N__48784;
    wire N__48783;
    wire N__48782;
    wire N__48781;
    wire N__48780;
    wire N__48779;
    wire N__48778;
    wire N__48777;
    wire N__48776;
    wire N__48775;
    wire N__48774;
    wire N__48773;
    wire N__48772;
    wire N__48771;
    wire N__48770;
    wire N__48769;
    wire N__48768;
    wire N__48767;
    wire N__48766;
    wire N__48765;
    wire N__48764;
    wire N__48763;
    wire N__48762;
    wire N__48761;
    wire N__48760;
    wire N__48759;
    wire N__48758;
    wire N__48757;
    wire N__48756;
    wire N__48755;
    wire N__48754;
    wire N__48753;
    wire N__48752;
    wire N__48751;
    wire N__48750;
    wire N__48749;
    wire N__48748;
    wire N__48747;
    wire N__48746;
    wire N__48745;
    wire N__48744;
    wire N__48743;
    wire N__48742;
    wire N__48741;
    wire N__48740;
    wire N__48739;
    wire N__48738;
    wire N__48737;
    wire N__48736;
    wire N__48735;
    wire N__48734;
    wire N__48733;
    wire N__48732;
    wire N__48731;
    wire N__48730;
    wire N__48729;
    wire N__48728;
    wire N__48727;
    wire N__48726;
    wire N__48725;
    wire N__48724;
    wire N__48723;
    wire N__48722;
    wire N__48721;
    wire N__48720;
    wire N__48719;
    wire N__48718;
    wire N__48717;
    wire N__48716;
    wire N__48715;
    wire N__48714;
    wire N__48713;
    wire N__48712;
    wire N__48711;
    wire N__48710;
    wire N__48709;
    wire N__48708;
    wire N__48707;
    wire N__48706;
    wire N__48705;
    wire N__48704;
    wire N__48703;
    wire N__48702;
    wire N__48701;
    wire N__48700;
    wire N__48699;
    wire N__48698;
    wire N__48697;
    wire N__48696;
    wire N__48695;
    wire N__48694;
    wire N__48693;
    wire N__48692;
    wire N__48691;
    wire N__48690;
    wire N__48689;
    wire N__48688;
    wire N__48687;
    wire N__48686;
    wire N__48685;
    wire N__48684;
    wire N__48683;
    wire N__48682;
    wire N__48681;
    wire N__48680;
    wire N__48679;
    wire N__48678;
    wire N__48677;
    wire N__48676;
    wire N__48675;
    wire N__48674;
    wire N__48673;
    wire N__48672;
    wire N__48671;
    wire N__48670;
    wire N__48669;
    wire N__48668;
    wire N__48667;
    wire N__48666;
    wire N__48665;
    wire N__48664;
    wire N__48663;
    wire N__48662;
    wire N__48661;
    wire N__48660;
    wire N__48659;
    wire N__48658;
    wire N__48657;
    wire N__48656;
    wire N__48655;
    wire N__48654;
    wire N__48653;
    wire N__48652;
    wire N__48651;
    wire N__48650;
    wire N__48649;
    wire N__48648;
    wire N__48647;
    wire N__48646;
    wire N__48643;
    wire N__48314;
    wire N__48311;
    wire N__48310;
    wire N__48309;
    wire N__48308;
    wire N__48305;
    wire N__48302;
    wire N__48299;
    wire N__48296;
    wire N__48293;
    wire N__48290;
    wire N__48287;
    wire N__48286;
    wire N__48283;
    wire N__48282;
    wire N__48281;
    wire N__48280;
    wire N__48279;
    wire N__48278;
    wire N__48277;
    wire N__48276;
    wire N__48275;
    wire N__48274;
    wire N__48273;
    wire N__48272;
    wire N__48271;
    wire N__48270;
    wire N__48269;
    wire N__48268;
    wire N__48267;
    wire N__48266;
    wire N__48265;
    wire N__48264;
    wire N__48263;
    wire N__48262;
    wire N__48261;
    wire N__48260;
    wire N__48259;
    wire N__48258;
    wire N__48257;
    wire N__48256;
    wire N__48255;
    wire N__48254;
    wire N__48253;
    wire N__48252;
    wire N__48251;
    wire N__48250;
    wire N__48249;
    wire N__48248;
    wire N__48247;
    wire N__48246;
    wire N__48245;
    wire N__48244;
    wire N__48243;
    wire N__48242;
    wire N__48241;
    wire N__48240;
    wire N__48239;
    wire N__48238;
    wire N__48237;
    wire N__48236;
    wire N__48235;
    wire N__48234;
    wire N__48233;
    wire N__48232;
    wire N__48231;
    wire N__48230;
    wire N__48229;
    wire N__48228;
    wire N__48227;
    wire N__48226;
    wire N__48225;
    wire N__48224;
    wire N__48223;
    wire N__48222;
    wire N__48221;
    wire N__48220;
    wire N__48219;
    wire N__48218;
    wire N__48217;
    wire N__48216;
    wire N__48215;
    wire N__48214;
    wire N__48213;
    wire N__48212;
    wire N__48211;
    wire N__48210;
    wire N__48209;
    wire N__48208;
    wire N__48207;
    wire N__48206;
    wire N__48205;
    wire N__48204;
    wire N__48203;
    wire N__48202;
    wire N__48201;
    wire N__48200;
    wire N__48199;
    wire N__48198;
    wire N__48197;
    wire N__48196;
    wire N__48195;
    wire N__48194;
    wire N__48193;
    wire N__48192;
    wire N__48191;
    wire N__48190;
    wire N__48189;
    wire N__48188;
    wire N__48187;
    wire N__48186;
    wire N__48185;
    wire N__48184;
    wire N__48183;
    wire N__48182;
    wire N__48181;
    wire N__48180;
    wire N__48179;
    wire N__48178;
    wire N__48177;
    wire N__48176;
    wire N__48175;
    wire N__48174;
    wire N__48173;
    wire N__48172;
    wire N__48171;
    wire N__48170;
    wire N__48169;
    wire N__48168;
    wire N__48167;
    wire N__48166;
    wire N__48165;
    wire N__48164;
    wire N__48163;
    wire N__48162;
    wire N__48161;
    wire N__48160;
    wire N__48159;
    wire N__48158;
    wire N__48157;
    wire N__48156;
    wire N__48155;
    wire N__48154;
    wire N__48153;
    wire N__48152;
    wire N__48151;
    wire N__48150;
    wire N__48149;
    wire N__48148;
    wire N__48147;
    wire N__48146;
    wire N__48145;
    wire N__48144;
    wire N__48143;
    wire N__48142;
    wire N__48141;
    wire N__48140;
    wire N__48139;
    wire N__48138;
    wire N__48137;
    wire N__48136;
    wire N__48135;
    wire N__48134;
    wire N__48133;
    wire N__48132;
    wire N__48131;
    wire N__48130;
    wire N__48129;
    wire N__48128;
    wire N__48127;
    wire N__48126;
    wire N__48125;
    wire N__48124;
    wire N__48123;
    wire N__48122;
    wire N__48121;
    wire N__47786;
    wire N__47783;
    wire N__47780;
    wire N__47777;
    wire N__47774;
    wire N__47773;
    wire N__47772;
    wire N__47765;
    wire N__47762;
    wire N__47759;
    wire N__47758;
    wire N__47757;
    wire N__47754;
    wire N__47749;
    wire N__47746;
    wire N__47743;
    wire N__47740;
    wire N__47737;
    wire N__47734;
    wire N__47731;
    wire N__47726;
    wire N__47723;
    wire N__47722;
    wire N__47721;
    wire N__47718;
    wire N__47713;
    wire N__47710;
    wire N__47705;
    wire N__47704;
    wire N__47701;
    wire N__47698;
    wire N__47695;
    wire N__47692;
    wire N__47691;
    wire N__47688;
    wire N__47685;
    wire N__47682;
    wire N__47679;
    wire N__47674;
    wire N__47671;
    wire N__47666;
    wire N__47665;
    wire N__47664;
    wire N__47661;
    wire N__47656;
    wire N__47653;
    wire N__47648;
    wire N__47645;
    wire N__47642;
    wire N__47639;
    wire N__47636;
    wire N__47635;
    wire N__47632;
    wire N__47629;
    wire N__47626;
    wire N__47621;
    wire N__47620;
    wire N__47617;
    wire N__47614;
    wire N__47609;
    wire N__47606;
    wire N__47605;
    wire N__47604;
    wire N__47601;
    wire N__47598;
    wire N__47595;
    wire N__47590;
    wire N__47587;
    wire N__47584;
    wire N__47581;
    wire N__47578;
    wire N__47573;
    wire N__47572;
    wire N__47571;
    wire N__47568;
    wire N__47565;
    wire N__47562;
    wire N__47559;
    wire N__47556;
    wire N__47553;
    wire N__47546;
    wire N__47545;
    wire N__47544;
    wire N__47543;
    wire N__47542;
    wire N__47541;
    wire N__47540;
    wire N__47539;
    wire N__47538;
    wire N__47537;
    wire N__47532;
    wire N__47517;
    wire N__47514;
    wire N__47509;
    wire N__47504;
    wire N__47501;
    wire N__47498;
    wire N__47495;
    wire N__47492;
    wire N__47489;
    wire N__47486;
    wire N__47483;
    wire N__47480;
    wire N__47477;
    wire N__47476;
    wire N__47475;
    wire N__47474;
    wire N__47473;
    wire N__47472;
    wire N__47471;
    wire N__47470;
    wire N__47469;
    wire N__47464;
    wire N__47463;
    wire N__47448;
    wire N__47445;
    wire N__47442;
    wire N__47439;
    wire N__47434;
    wire N__47431;
    wire N__47428;
    wire N__47425;
    wire N__47422;
    wire N__47419;
    wire N__47414;
    wire N__47411;
    wire N__47408;
    wire N__47405;
    wire N__47404;
    wire N__47401;
    wire N__47396;
    wire N__47395;
    wire N__47392;
    wire N__47389;
    wire N__47386;
    wire N__47381;
    wire N__47380;
    wire N__47377;
    wire N__47372;
    wire N__47371;
    wire N__47368;
    wire N__47365;
    wire N__47362;
    wire N__47357;
    wire N__47354;
    wire N__47351;
    wire N__47348;
    wire N__47347;
    wire N__47346;
    wire N__47343;
    wire N__47340;
    wire N__47337;
    wire N__47334;
    wire N__47331;
    wire N__47324;
    wire N__47323;
    wire N__47320;
    wire N__47319;
    wire N__47316;
    wire N__47313;
    wire N__47310;
    wire N__47307;
    wire N__47304;
    wire N__47299;
    wire N__47298;
    wire N__47295;
    wire N__47292;
    wire N__47289;
    wire N__47282;
    wire N__47281;
    wire N__47276;
    wire N__47273;
    wire N__47270;
    wire N__47269;
    wire N__47266;
    wire N__47263;
    wire N__47260;
    wire N__47257;
    wire N__47254;
    wire N__47251;
    wire N__47248;
    wire N__47245;
    wire N__47240;
    wire N__47237;
    wire N__47234;
    wire N__47231;
    wire N__47230;
    wire N__47227;
    wire N__47226;
    wire N__47223;
    wire N__47220;
    wire N__47217;
    wire N__47210;
    wire N__47209;
    wire N__47206;
    wire N__47205;
    wire N__47202;
    wire N__47199;
    wire N__47196;
    wire N__47195;
    wire N__47192;
    wire N__47189;
    wire N__47186;
    wire N__47183;
    wire N__47178;
    wire N__47175;
    wire N__47172;
    wire N__47165;
    wire N__47164;
    wire N__47163;
    wire N__47162;
    wire N__47161;
    wire N__47160;
    wire N__47157;
    wire N__47154;
    wire N__47151;
    wire N__47148;
    wire N__47147;
    wire N__47146;
    wire N__47145;
    wire N__47144;
    wire N__47143;
    wire N__47142;
    wire N__47141;
    wire N__47140;
    wire N__47139;
    wire N__47138;
    wire N__47137;
    wire N__47136;
    wire N__47135;
    wire N__47134;
    wire N__47133;
    wire N__47132;
    wire N__47131;
    wire N__47130;
    wire N__47125;
    wire N__47124;
    wire N__47123;
    wire N__47122;
    wire N__47121;
    wire N__47120;
    wire N__47119;
    wire N__47118;
    wire N__47117;
    wire N__47116;
    wire N__47115;
    wire N__47114;
    wire N__47113;
    wire N__47112;
    wire N__47111;
    wire N__47110;
    wire N__47109;
    wire N__47108;
    wire N__47107;
    wire N__47106;
    wire N__47103;
    wire N__47096;
    wire N__47091;
    wire N__47090;
    wire N__47089;
    wire N__47088;
    wire N__47085;
    wire N__47084;
    wire N__47083;
    wire N__47082;
    wire N__47081;
    wire N__47072;
    wire N__47067;
    wire N__47066;
    wire N__47065;
    wire N__47064;
    wire N__47063;
    wire N__47062;
    wire N__47061;
    wire N__47060;
    wire N__47059;
    wire N__47058;
    wire N__47057;
    wire N__47056;
    wire N__47055;
    wire N__47054;
    wire N__47053;
    wire N__47052;
    wire N__47051;
    wire N__47048;
    wire N__47045;
    wire N__47034;
    wire N__47029;
    wire N__47026;
    wire N__47021;
    wire N__47018;
    wire N__47013;
    wire N__47004;
    wire N__46995;
    wire N__46994;
    wire N__46993;
    wire N__46992;
    wire N__46991;
    wire N__46990;
    wire N__46985;
    wire N__46978;
    wire N__46977;
    wire N__46976;
    wire N__46975;
    wire N__46974;
    wire N__46971;
    wire N__46964;
    wire N__46957;
    wire N__46954;
    wire N__46949;
    wire N__46946;
    wire N__46943;
    wire N__46940;
    wire N__46937;
    wire N__46936;
    wire N__46935;
    wire N__46934;
    wire N__46933;
    wire N__46932;
    wire N__46931;
    wire N__46930;
    wire N__46929;
    wire N__46928;
    wire N__46927;
    wire N__46926;
    wire N__46925;
    wire N__46924;
    wire N__46923;
    wire N__46922;
    wire N__46921;
    wire N__46916;
    wire N__46907;
    wire N__46900;
    wire N__46893;
    wire N__46884;
    wire N__46877;
    wire N__46870;
    wire N__46861;
    wire N__46850;
    wire N__46845;
    wire N__46842;
    wire N__46841;
    wire N__46834;
    wire N__46823;
    wire N__46814;
    wire N__46811;
    wire N__46808;
    wire N__46801;
    wire N__46796;
    wire N__46785;
    wire N__46776;
    wire N__46773;
    wire N__46764;
    wire N__46757;
    wire N__46750;
    wire N__46747;
    wire N__46740;
    wire N__46715;
    wire N__46714;
    wire N__46709;
    wire N__46706;
    wire N__46703;
    wire N__46702;
    wire N__46701;
    wire N__46700;
    wire N__46699;
    wire N__46698;
    wire N__46697;
    wire N__46696;
    wire N__46695;
    wire N__46694;
    wire N__46691;
    wire N__46688;
    wire N__46687;
    wire N__46686;
    wire N__46685;
    wire N__46684;
    wire N__46683;
    wire N__46682;
    wire N__46681;
    wire N__46680;
    wire N__46679;
    wire N__46678;
    wire N__46677;
    wire N__46676;
    wire N__46675;
    wire N__46672;
    wire N__46669;
    wire N__46666;
    wire N__46665;
    wire N__46664;
    wire N__46663;
    wire N__46662;
    wire N__46661;
    wire N__46658;
    wire N__46657;
    wire N__46648;
    wire N__46643;
    wire N__46640;
    wire N__46637;
    wire N__46628;
    wire N__46619;
    wire N__46616;
    wire N__46615;
    wire N__46614;
    wire N__46611;
    wire N__46610;
    wire N__46609;
    wire N__46608;
    wire N__46607;
    wire N__46606;
    wire N__46605;
    wire N__46604;
    wire N__46603;
    wire N__46602;
    wire N__46601;
    wire N__46598;
    wire N__46595;
    wire N__46594;
    wire N__46593;
    wire N__46592;
    wire N__46591;
    wire N__46590;
    wire N__46589;
    wire N__46586;
    wire N__46583;
    wire N__46580;
    wire N__46571;
    wire N__46568;
    wire N__46565;
    wire N__46562;
    wire N__46557;
    wire N__46554;
    wire N__46547;
    wire N__46544;
    wire N__46541;
    wire N__46538;
    wire N__46531;
    wire N__46522;
    wire N__46515;
    wire N__46512;
    wire N__46509;
    wire N__46500;
    wire N__46497;
    wire N__46494;
    wire N__46477;
    wire N__46474;
    wire N__46471;
    wire N__46468;
    wire N__46465;
    wire N__46454;
    wire N__46451;
    wire N__46448;
    wire N__46439;
    wire N__46436;
    wire N__46427;
    wire N__46422;
    wire N__46415;
    wire N__46414;
    wire N__46413;
    wire N__46410;
    wire N__46407;
    wire N__46400;
    wire N__46397;
    wire N__46396;
    wire N__46395;
    wire N__46394;
    wire N__46391;
    wire N__46388;
    wire N__46385;
    wire N__46382;
    wire N__46379;
    wire N__46374;
    wire N__46371;
    wire N__46368;
    wire N__46365;
    wire N__46362;
    wire N__46355;
    wire N__46354;
    wire N__46353;
    wire N__46350;
    wire N__46347;
    wire N__46344;
    wire N__46337;
    wire N__46336;
    wire N__46335;
    wire N__46332;
    wire N__46329;
    wire N__46326;
    wire N__46323;
    wire N__46320;
    wire N__46319;
    wire N__46316;
    wire N__46313;
    wire N__46310;
    wire N__46307;
    wire N__46298;
    wire N__46295;
    wire N__46292;
    wire N__46291;
    wire N__46288;
    wire N__46287;
    wire N__46284;
    wire N__46281;
    wire N__46278;
    wire N__46271;
    wire N__46268;
    wire N__46267;
    wire N__46264;
    wire N__46261;
    wire N__46256;
    wire N__46253;
    wire N__46250;
    wire N__46247;
    wire N__46246;
    wire N__46243;
    wire N__46242;
    wire N__46239;
    wire N__46238;
    wire N__46235;
    wire N__46232;
    wire N__46229;
    wire N__46228;
    wire N__46225;
    wire N__46222;
    wire N__46219;
    wire N__46216;
    wire N__46213;
    wire N__46202;
    wire N__46201;
    wire N__46198;
    wire N__46195;
    wire N__46192;
    wire N__46191;
    wire N__46190;
    wire N__46189;
    wire N__46186;
    wire N__46183;
    wire N__46178;
    wire N__46175;
    wire N__46168;
    wire N__46163;
    wire N__46160;
    wire N__46159;
    wire N__46156;
    wire N__46153;
    wire N__46150;
    wire N__46149;
    wire N__46146;
    wire N__46143;
    wire N__46140;
    wire N__46137;
    wire N__46130;
    wire N__46129;
    wire N__46124;
    wire N__46121;
    wire N__46118;
    wire N__46117;
    wire N__46116;
    wire N__46115;
    wire N__46114;
    wire N__46113;
    wire N__46112;
    wire N__46111;
    wire N__46110;
    wire N__46109;
    wire N__46108;
    wire N__46107;
    wire N__46082;
    wire N__46079;
    wire N__46076;
    wire N__46075;
    wire N__46072;
    wire N__46069;
    wire N__46068;
    wire N__46065;
    wire N__46062;
    wire N__46059;
    wire N__46056;
    wire N__46053;
    wire N__46048;
    wire N__46045;
    wire N__46044;
    wire N__46041;
    wire N__46038;
    wire N__46035;
    wire N__46028;
    wire N__46025;
    wire N__46024;
    wire N__46021;
    wire N__46020;
    wire N__46017;
    wire N__46014;
    wire N__46011;
    wire N__46004;
    wire N__46001;
    wire N__46000;
    wire N__45997;
    wire N__45996;
    wire N__45993;
    wire N__45990;
    wire N__45987;
    wire N__45980;
    wire N__45977;
    wire N__45976;
    wire N__45975;
    wire N__45974;
    wire N__45971;
    wire N__45968;
    wire N__45965;
    wire N__45962;
    wire N__45957;
    wire N__45954;
    wire N__45949;
    wire N__45944;
    wire N__45941;
    wire N__45938;
    wire N__45935;
    wire N__45932;
    wire N__45929;
    wire N__45926;
    wire N__45923;
    wire N__45920;
    wire N__45919;
    wire N__45914;
    wire N__45911;
    wire N__45908;
    wire N__45907;
    wire N__45904;
    wire N__45901;
    wire N__45896;
    wire N__45895;
    wire N__45892;
    wire N__45891;
    wire N__45888;
    wire N__45885;
    wire N__45882;
    wire N__45875;
    wire N__45874;
    wire N__45873;
    wire N__45870;
    wire N__45867;
    wire N__45864;
    wire N__45861;
    wire N__45858;
    wire N__45851;
    wire N__45850;
    wire N__45847;
    wire N__45844;
    wire N__45841;
    wire N__45836;
    wire N__45833;
    wire N__45830;
    wire N__45829;
    wire N__45826;
    wire N__45823;
    wire N__45820;
    wire N__45817;
    wire N__45814;
    wire N__45811;
    wire N__45806;
    wire N__45803;
    wire N__45802;
    wire N__45799;
    wire N__45796;
    wire N__45791;
    wire N__45788;
    wire N__45787;
    wire N__45786;
    wire N__45785;
    wire N__45782;
    wire N__45777;
    wire N__45774;
    wire N__45771;
    wire N__45768;
    wire N__45765;
    wire N__45758;
    wire N__45755;
    wire N__45752;
    wire N__45749;
    wire N__45746;
    wire N__45745;
    wire N__45744;
    wire N__45737;
    wire N__45734;
    wire N__45733;
    wire N__45730;
    wire N__45729;
    wire N__45728;
    wire N__45725;
    wire N__45718;
    wire N__45713;
    wire N__45712;
    wire N__45711;
    wire N__45710;
    wire N__45707;
    wire N__45700;
    wire N__45695;
    wire N__45692;
    wire N__45689;
    wire N__45686;
    wire N__45683;
    wire N__45680;
    wire N__45677;
    wire N__45674;
    wire N__45671;
    wire N__45668;
    wire N__45665;
    wire N__45662;
    wire N__45659;
    wire N__45656;
    wire N__45653;
    wire N__45650;
    wire N__45647;
    wire N__45644;
    wire N__45641;
    wire N__45638;
    wire N__45635;
    wire N__45632;
    wire N__45629;
    wire N__45626;
    wire N__45623;
    wire N__45620;
    wire N__45617;
    wire N__45614;
    wire N__45611;
    wire N__45610;
    wire N__45607;
    wire N__45606;
    wire N__45603;
    wire N__45598;
    wire N__45593;
    wire N__45592;
    wire N__45589;
    wire N__45584;
    wire N__45581;
    wire N__45578;
    wire N__45577;
    wire N__45576;
    wire N__45573;
    wire N__45568;
    wire N__45563;
    wire N__45560;
    wire N__45557;
    wire N__45554;
    wire N__45551;
    wire N__45550;
    wire N__45547;
    wire N__45544;
    wire N__45541;
    wire N__45540;
    wire N__45535;
    wire N__45532;
    wire N__45527;
    wire N__45524;
    wire N__45523;
    wire N__45522;
    wire N__45519;
    wire N__45516;
    wire N__45513;
    wire N__45508;
    wire N__45507;
    wire N__45504;
    wire N__45501;
    wire N__45498;
    wire N__45491;
    wire N__45488;
    wire N__45485;
    wire N__45482;
    wire N__45479;
    wire N__45476;
    wire N__45475;
    wire N__45472;
    wire N__45469;
    wire N__45464;
    wire N__45461;
    wire N__45458;
    wire N__45455;
    wire N__45454;
    wire N__45451;
    wire N__45448;
    wire N__45443;
    wire N__45440;
    wire N__45437;
    wire N__45434;
    wire N__45431;
    wire N__45428;
    wire N__45425;
    wire N__45422;
    wire N__45421;
    wire N__45418;
    wire N__45415;
    wire N__45410;
    wire N__45407;
    wire N__45404;
    wire N__45401;
    wire N__45398;
    wire N__45395;
    wire N__45392;
    wire N__45391;
    wire N__45388;
    wire N__45385;
    wire N__45380;
    wire N__45377;
    wire N__45374;
    wire N__45371;
    wire N__45368;
    wire N__45365;
    wire N__45362;
    wire N__45359;
    wire N__45356;
    wire N__45353;
    wire N__45350;
    wire N__45347;
    wire N__45344;
    wire N__45341;
    wire N__45338;
    wire N__45335;
    wire N__45332;
    wire N__45329;
    wire N__45326;
    wire N__45323;
    wire N__45320;
    wire N__45317;
    wire N__45314;
    wire N__45311;
    wire N__45308;
    wire N__45305;
    wire N__45302;
    wire N__45299;
    wire N__45296;
    wire N__45293;
    wire N__45290;
    wire N__45287;
    wire N__45284;
    wire N__45283;
    wire N__45280;
    wire N__45277;
    wire N__45272;
    wire N__45269;
    wire N__45266;
    wire N__45265;
    wire N__45262;
    wire N__45259;
    wire N__45254;
    wire N__45251;
    wire N__45248;
    wire N__45245;
    wire N__45242;
    wire N__45239;
    wire N__45236;
    wire N__45233;
    wire N__45230;
    wire N__45229;
    wire N__45226;
    wire N__45223;
    wire N__45218;
    wire N__45215;
    wire N__45212;
    wire N__45209;
    wire N__45206;
    wire N__45203;
    wire N__45202;
    wire N__45199;
    wire N__45196;
    wire N__45191;
    wire N__45188;
    wire N__45185;
    wire N__45182;
    wire N__45179;
    wire N__45176;
    wire N__45175;
    wire N__45172;
    wire N__45169;
    wire N__45164;
    wire N__45161;
    wire N__45158;
    wire N__45155;
    wire N__45152;
    wire N__45149;
    wire N__45146;
    wire N__45145;
    wire N__45142;
    wire N__45139;
    wire N__45136;
    wire N__45131;
    wire N__45128;
    wire N__45125;
    wire N__45122;
    wire N__45121;
    wire N__45118;
    wire N__45115;
    wire N__45110;
    wire N__45107;
    wire N__45104;
    wire N__45101;
    wire N__45098;
    wire N__45095;
    wire N__45092;
    wire N__45089;
    wire N__45088;
    wire N__45085;
    wire N__45082;
    wire N__45077;
    wire N__45076;
    wire N__45073;
    wire N__45072;
    wire N__45069;
    wire N__45066;
    wire N__45063;
    wire N__45056;
    wire N__45055;
    wire N__45052;
    wire N__45049;
    wire N__45048;
    wire N__45045;
    wire N__45042;
    wire N__45039;
    wire N__45036;
    wire N__45033;
    wire N__45030;
    wire N__45029;
    wire N__45026;
    wire N__45023;
    wire N__45020;
    wire N__45017;
    wire N__45008;
    wire N__45005;
    wire N__45004;
    wire N__45003;
    wire N__45002;
    wire N__44999;
    wire N__44996;
    wire N__44993;
    wire N__44990;
    wire N__44987;
    wire N__44982;
    wire N__44979;
    wire N__44976;
    wire N__44971;
    wire N__44966;
    wire N__44965;
    wire N__44964;
    wire N__44961;
    wire N__44958;
    wire N__44955;
    wire N__44952;
    wire N__44945;
    wire N__44942;
    wire N__44941;
    wire N__44938;
    wire N__44937;
    wire N__44934;
    wire N__44931;
    wire N__44928;
    wire N__44921;
    wire N__44920;
    wire N__44919;
    wire N__44916;
    wire N__44915;
    wire N__44912;
    wire N__44909;
    wire N__44906;
    wire N__44903;
    wire N__44898;
    wire N__44893;
    wire N__44890;
    wire N__44887;
    wire N__44882;
    wire N__44879;
    wire N__44878;
    wire N__44877;
    wire N__44874;
    wire N__44871;
    wire N__44868;
    wire N__44865;
    wire N__44862;
    wire N__44855;
    wire N__44854;
    wire N__44853;
    wire N__44850;
    wire N__44849;
    wire N__44846;
    wire N__44843;
    wire N__44840;
    wire N__44837;
    wire N__44834;
    wire N__44831;
    wire N__44826;
    wire N__44823;
    wire N__44818;
    wire N__44813;
    wire N__44810;
    wire N__44809;
    wire N__44806;
    wire N__44805;
    wire N__44802;
    wire N__44799;
    wire N__44796;
    wire N__44789;
    wire N__44788;
    wire N__44787;
    wire N__44784;
    wire N__44781;
    wire N__44778;
    wire N__44773;
    wire N__44770;
    wire N__44767;
    wire N__44766;
    wire N__44763;
    wire N__44760;
    wire N__44757;
    wire N__44750;
    wire N__44747;
    wire N__44746;
    wire N__44741;
    wire N__44738;
    wire N__44735;
    wire N__44734;
    wire N__44733;
    wire N__44730;
    wire N__44727;
    wire N__44724;
    wire N__44721;
    wire N__44718;
    wire N__44715;
    wire N__44712;
    wire N__44709;
    wire N__44702;
    wire N__44699;
    wire N__44696;
    wire N__44693;
    wire N__44690;
    wire N__44687;
    wire N__44686;
    wire N__44683;
    wire N__44680;
    wire N__44675;
    wire N__44672;
    wire N__44669;
    wire N__44666;
    wire N__44663;
    wire N__44660;
    wire N__44657;
    wire N__44654;
    wire N__44651;
    wire N__44650;
    wire N__44647;
    wire N__44644;
    wire N__44639;
    wire N__44636;
    wire N__44633;
    wire N__44632;
    wire N__44631;
    wire N__44628;
    wire N__44627;
    wire N__44624;
    wire N__44621;
    wire N__44618;
    wire N__44613;
    wire N__44606;
    wire N__44603;
    wire N__44600;
    wire N__44597;
    wire N__44594;
    wire N__44591;
    wire N__44590;
    wire N__44587;
    wire N__44584;
    wire N__44579;
    wire N__44578;
    wire N__44577;
    wire N__44572;
    wire N__44569;
    wire N__44564;
    wire N__44563;
    wire N__44560;
    wire N__44557;
    wire N__44554;
    wire N__44551;
    wire N__44546;
    wire N__44543;
    wire N__44540;
    wire N__44537;
    wire N__44534;
    wire N__44531;
    wire N__44528;
    wire N__44525;
    wire N__44522;
    wire N__44519;
    wire N__44516;
    wire N__44513;
    wire N__44510;
    wire N__44509;
    wire N__44506;
    wire N__44503;
    wire N__44498;
    wire N__44495;
    wire N__44492;
    wire N__44491;
    wire N__44488;
    wire N__44485;
    wire N__44480;
    wire N__44477;
    wire N__44476;
    wire N__44473;
    wire N__44470;
    wire N__44467;
    wire N__44464;
    wire N__44459;
    wire N__44456;
    wire N__44455;
    wire N__44452;
    wire N__44449;
    wire N__44444;
    wire N__44441;
    wire N__44438;
    wire N__44435;
    wire N__44432;
    wire N__44429;
    wire N__44426;
    wire N__44423;
    wire N__44420;
    wire N__44419;
    wire N__44416;
    wire N__44413;
    wire N__44408;
    wire N__44405;
    wire N__44402;
    wire N__44399;
    wire N__44396;
    wire N__44395;
    wire N__44394;
    wire N__44391;
    wire N__44388;
    wire N__44385;
    wire N__44382;
    wire N__44379;
    wire N__44372;
    wire N__44371;
    wire N__44368;
    wire N__44367;
    wire N__44364;
    wire N__44361;
    wire N__44358;
    wire N__44351;
    wire N__44350;
    wire N__44349;
    wire N__44346;
    wire N__44345;
    wire N__44342;
    wire N__44339;
    wire N__44336;
    wire N__44333;
    wire N__44330;
    wire N__44327;
    wire N__44324;
    wire N__44321;
    wire N__44318;
    wire N__44315;
    wire N__44310;
    wire N__44303;
    wire N__44302;
    wire N__44299;
    wire N__44298;
    wire N__44297;
    wire N__44294;
    wire N__44291;
    wire N__44288;
    wire N__44285;
    wire N__44282;
    wire N__44279;
    wire N__44276;
    wire N__44273;
    wire N__44268;
    wire N__44263;
    wire N__44258;
    wire N__44257;
    wire N__44254;
    wire N__44253;
    wire N__44250;
    wire N__44247;
    wire N__44244;
    wire N__44237;
    wire N__44234;
    wire N__44233;
    wire N__44232;
    wire N__44231;
    wire N__44226;
    wire N__44223;
    wire N__44220;
    wire N__44217;
    wire N__44214;
    wire N__44211;
    wire N__44208;
    wire N__44203;
    wire N__44198;
    wire N__44197;
    wire N__44196;
    wire N__44193;
    wire N__44188;
    wire N__44183;
    wire N__44180;
    wire N__44179;
    wire N__44174;
    wire N__44171;
    wire N__44168;
    wire N__44165;
    wire N__44164;
    wire N__44163;
    wire N__44160;
    wire N__44157;
    wire N__44152;
    wire N__44147;
    wire N__44146;
    wire N__44141;
    wire N__44138;
    wire N__44137;
    wire N__44136;
    wire N__44133;
    wire N__44126;
    wire N__44123;
    wire N__44120;
    wire N__44117;
    wire N__44116;
    wire N__44113;
    wire N__44112;
    wire N__44109;
    wire N__44108;
    wire N__44105;
    wire N__44102;
    wire N__44099;
    wire N__44096;
    wire N__44095;
    wire N__44092;
    wire N__44089;
    wire N__44086;
    wire N__44083;
    wire N__44080;
    wire N__44075;
    wire N__44072;
    wire N__44069;
    wire N__44066;
    wire N__44057;
    wire N__44056;
    wire N__44055;
    wire N__44052;
    wire N__44049;
    wire N__44046;
    wire N__44043;
    wire N__44042;
    wire N__44039;
    wire N__44036;
    wire N__44033;
    wire N__44030;
    wire N__44027;
    wire N__44018;
    wire N__44017;
    wire N__44016;
    wire N__44013;
    wire N__44010;
    wire N__44007;
    wire N__44000;
    wire N__43999;
    wire N__43996;
    wire N__43995;
    wire N__43992;
    wire N__43989;
    wire N__43986;
    wire N__43985;
    wire N__43978;
    wire N__43975;
    wire N__43970;
    wire N__43967;
    wire N__43966;
    wire N__43965;
    wire N__43964;
    wire N__43961;
    wire N__43958;
    wire N__43955;
    wire N__43952;
    wire N__43949;
    wire N__43940;
    wire N__43939;
    wire N__43938;
    wire N__43935;
    wire N__43934;
    wire N__43931;
    wire N__43928;
    wire N__43925;
    wire N__43922;
    wire N__43919;
    wire N__43916;
    wire N__43911;
    wire N__43908;
    wire N__43905;
    wire N__43902;
    wire N__43895;
    wire N__43892;
    wire N__43889;
    wire N__43886;
    wire N__43883;
    wire N__43880;
    wire N__43877;
    wire N__43874;
    wire N__43873;
    wire N__43870;
    wire N__43869;
    wire N__43868;
    wire N__43865;
    wire N__43862;
    wire N__43859;
    wire N__43856;
    wire N__43853;
    wire N__43848;
    wire N__43845;
    wire N__43842;
    wire N__43839;
    wire N__43832;
    wire N__43829;
    wire N__43828;
    wire N__43825;
    wire N__43824;
    wire N__43821;
    wire N__43818;
    wire N__43815;
    wire N__43808;
    wire N__43805;
    wire N__43802;
    wire N__43801;
    wire N__43798;
    wire N__43795;
    wire N__43790;
    wire N__43789;
    wire N__43788;
    wire N__43785;
    wire N__43780;
    wire N__43775;
    wire N__43772;
    wire N__43771;
    wire N__43770;
    wire N__43767;
    wire N__43764;
    wire N__43761;
    wire N__43756;
    wire N__43751;
    wire N__43748;
    wire N__43747;
    wire N__43746;
    wire N__43741;
    wire N__43738;
    wire N__43735;
    wire N__43730;
    wire N__43727;
    wire N__43724;
    wire N__43723;
    wire N__43722;
    wire N__43717;
    wire N__43714;
    wire N__43711;
    wire N__43706;
    wire N__43703;
    wire N__43702;
    wire N__43701;
    wire N__43696;
    wire N__43693;
    wire N__43690;
    wire N__43685;
    wire N__43682;
    wire N__43681;
    wire N__43678;
    wire N__43677;
    wire N__43672;
    wire N__43669;
    wire N__43666;
    wire N__43661;
    wire N__43658;
    wire N__43655;
    wire N__43652;
    wire N__43649;
    wire N__43646;
    wire N__43643;
    wire N__43640;
    wire N__43637;
    wire N__43634;
    wire N__43631;
    wire N__43628;
    wire N__43625;
    wire N__43622;
    wire N__43619;
    wire N__43618;
    wire N__43617;
    wire N__43614;
    wire N__43611;
    wire N__43608;
    wire N__43605;
    wire N__43600;
    wire N__43597;
    wire N__43592;
    wire N__43589;
    wire N__43588;
    wire N__43585;
    wire N__43582;
    wire N__43581;
    wire N__43580;
    wire N__43575;
    wire N__43570;
    wire N__43565;
    wire N__43564;
    wire N__43561;
    wire N__43560;
    wire N__43559;
    wire N__43556;
    wire N__43553;
    wire N__43550;
    wire N__43547;
    wire N__43544;
    wire N__43539;
    wire N__43536;
    wire N__43533;
    wire N__43530;
    wire N__43527;
    wire N__43520;
    wire N__43519;
    wire N__43518;
    wire N__43515;
    wire N__43512;
    wire N__43509;
    wire N__43506;
    wire N__43499;
    wire N__43498;
    wire N__43497;
    wire N__43494;
    wire N__43491;
    wire N__43488;
    wire N__43481;
    wire N__43480;
    wire N__43477;
    wire N__43474;
    wire N__43473;
    wire N__43472;
    wire N__43469;
    wire N__43466;
    wire N__43463;
    wire N__43460;
    wire N__43457;
    wire N__43454;
    wire N__43449;
    wire N__43442;
    wire N__43439;
    wire N__43436;
    wire N__43433;
    wire N__43430;
    wire N__43427;
    wire N__43424;
    wire N__43421;
    wire N__43418;
    wire N__43415;
    wire N__43412;
    wire N__43409;
    wire N__43406;
    wire N__43405;
    wire N__43402;
    wire N__43401;
    wire N__43398;
    wire N__43395;
    wire N__43392;
    wire N__43385;
    wire N__43384;
    wire N__43383;
    wire N__43380;
    wire N__43377;
    wire N__43374;
    wire N__43371;
    wire N__43368;
    wire N__43365;
    wire N__43362;
    wire N__43359;
    wire N__43358;
    wire N__43355;
    wire N__43352;
    wire N__43349;
    wire N__43346;
    wire N__43337;
    wire N__43334;
    wire N__43333;
    wire N__43330;
    wire N__43327;
    wire N__43322;
    wire N__43319;
    wire N__43318;
    wire N__43317;
    wire N__43312;
    wire N__43309;
    wire N__43306;
    wire N__43303;
    wire N__43300;
    wire N__43299;
    wire N__43296;
    wire N__43293;
    wire N__43290;
    wire N__43283;
    wire N__43282;
    wire N__43277;
    wire N__43274;
    wire N__43273;
    wire N__43272;
    wire N__43269;
    wire N__43266;
    wire N__43263;
    wire N__43260;
    wire N__43257;
    wire N__43250;
    wire N__43249;
    wire N__43246;
    wire N__43245;
    wire N__43242;
    wire N__43239;
    wire N__43236;
    wire N__43233;
    wire N__43232;
    wire N__43229;
    wire N__43224;
    wire N__43221;
    wire N__43218;
    wire N__43215;
    wire N__43212;
    wire N__43205;
    wire N__43204;
    wire N__43199;
    wire N__43196;
    wire N__43193;
    wire N__43192;
    wire N__43187;
    wire N__43184;
    wire N__43181;
    wire N__43178;
    wire N__43177;
    wire N__43174;
    wire N__43173;
    wire N__43170;
    wire N__43167;
    wire N__43164;
    wire N__43157;
    wire N__43156;
    wire N__43155;
    wire N__43152;
    wire N__43149;
    wire N__43146;
    wire N__43145;
    wire N__43142;
    wire N__43139;
    wire N__43136;
    wire N__43133;
    wire N__43124;
    wire N__43123;
    wire N__43118;
    wire N__43115;
    wire N__43112;
    wire N__43111;
    wire N__43106;
    wire N__43103;
    wire N__43100;
    wire N__43097;
    wire N__43094;
    wire N__43093;
    wire N__43090;
    wire N__43087;
    wire N__43084;
    wire N__43079;
    wire N__43076;
    wire N__43073;
    wire N__43070;
    wire N__43069;
    wire N__43068;
    wire N__43067;
    wire N__43064;
    wire N__43061;
    wire N__43058;
    wire N__43057;
    wire N__43054;
    wire N__43047;
    wire N__43044;
    wire N__43037;
    wire N__43034;
    wire N__43031;
    wire N__43028;
    wire N__43025;
    wire N__43024;
    wire N__43021;
    wire N__43018;
    wire N__43013;
    wire N__43010;
    wire N__43007;
    wire N__43006;
    wire N__43003;
    wire N__43000;
    wire N__42999;
    wire N__42996;
    wire N__42993;
    wire N__42990;
    wire N__42987;
    wire N__42984;
    wire N__42981;
    wire N__42978;
    wire N__42973;
    wire N__42968;
    wire N__42967;
    wire N__42966;
    wire N__42963;
    wire N__42962;
    wire N__42959;
    wire N__42956;
    wire N__42953;
    wire N__42950;
    wire N__42947;
    wire N__42942;
    wire N__42941;
    wire N__42936;
    wire N__42933;
    wire N__42930;
    wire N__42929;
    wire N__42926;
    wire N__42921;
    wire N__42918;
    wire N__42913;
    wire N__42908;
    wire N__42907;
    wire N__42904;
    wire N__42901;
    wire N__42898;
    wire N__42895;
    wire N__42890;
    wire N__42889;
    wire N__42884;
    wire N__42881;
    wire N__42880;
    wire N__42875;
    wire N__42872;
    wire N__42869;
    wire N__42868;
    wire N__42863;
    wire N__42860;
    wire N__42859;
    wire N__42854;
    wire N__42851;
    wire N__42850;
    wire N__42845;
    wire N__42842;
    wire N__42841;
    wire N__42836;
    wire N__42833;
    wire N__42832;
    wire N__42827;
    wire N__42824;
    wire N__42823;
    wire N__42820;
    wire N__42817;
    wire N__42812;
    wire N__42809;
    wire N__42808;
    wire N__42805;
    wire N__42802;
    wire N__42797;
    wire N__42794;
    wire N__42791;
    wire N__42790;
    wire N__42787;
    wire N__42784;
    wire N__42779;
    wire N__42776;
    wire N__42773;
    wire N__42772;
    wire N__42769;
    wire N__42766;
    wire N__42763;
    wire N__42758;
    wire N__42755;
    wire N__42754;
    wire N__42751;
    wire N__42748;
    wire N__42745;
    wire N__42740;
    wire N__42739;
    wire N__42734;
    wire N__42731;
    wire N__42730;
    wire N__42725;
    wire N__42722;
    wire N__42721;
    wire N__42716;
    wire N__42713;
    wire N__42710;
    wire N__42709;
    wire N__42708;
    wire N__42705;
    wire N__42700;
    wire N__42699;
    wire N__42696;
    wire N__42693;
    wire N__42690;
    wire N__42687;
    wire N__42684;
    wire N__42677;
    wire N__42674;
    wire N__42671;
    wire N__42668;
    wire N__42667;
    wire N__42664;
    wire N__42661;
    wire N__42656;
    wire N__42653;
    wire N__42652;
    wire N__42649;
    wire N__42646;
    wire N__42641;
    wire N__42638;
    wire N__42635;
    wire N__42634;
    wire N__42633;
    wire N__42630;
    wire N__42627;
    wire N__42624;
    wire N__42619;
    wire N__42616;
    wire N__42613;
    wire N__42610;
    wire N__42607;
    wire N__42604;
    wire N__42601;
    wire N__42598;
    wire N__42593;
    wire N__42590;
    wire N__42587;
    wire N__42586;
    wire N__42583;
    wire N__42580;
    wire N__42575;
    wire N__42572;
    wire N__42569;
    wire N__42566;
    wire N__42563;
    wire N__42560;
    wire N__42557;
    wire N__42554;
    wire N__42553;
    wire N__42552;
    wire N__42549;
    wire N__42546;
    wire N__42543;
    wire N__42540;
    wire N__42533;
    wire N__42530;
    wire N__42527;
    wire N__42524;
    wire N__42523;
    wire N__42522;
    wire N__42519;
    wire N__42516;
    wire N__42513;
    wire N__42512;
    wire N__42507;
    wire N__42504;
    wire N__42501;
    wire N__42494;
    wire N__42491;
    wire N__42488;
    wire N__42487;
    wire N__42486;
    wire N__42483;
    wire N__42480;
    wire N__42477;
    wire N__42474;
    wire N__42473;
    wire N__42470;
    wire N__42465;
    wire N__42462;
    wire N__42455;
    wire N__42452;
    wire N__42449;
    wire N__42446;
    wire N__42445;
    wire N__42442;
    wire N__42441;
    wire N__42438;
    wire N__42435;
    wire N__42432;
    wire N__42425;
    wire N__42422;
    wire N__42419;
    wire N__42418;
    wire N__42417;
    wire N__42414;
    wire N__42413;
    wire N__42408;
    wire N__42405;
    wire N__42402;
    wire N__42399;
    wire N__42392;
    wire N__42389;
    wire N__42388;
    wire N__42385;
    wire N__42384;
    wire N__42381;
    wire N__42380;
    wire N__42377;
    wire N__42374;
    wire N__42371;
    wire N__42368;
    wire N__42365;
    wire N__42356;
    wire N__42355;
    wire N__42352;
    wire N__42349;
    wire N__42348;
    wire N__42345;
    wire N__42344;
    wire N__42341;
    wire N__42340;
    wire N__42337;
    wire N__42334;
    wire N__42331;
    wire N__42328;
    wire N__42325;
    wire N__42322;
    wire N__42319;
    wire N__42316;
    wire N__42313;
    wire N__42310;
    wire N__42307;
    wire N__42302;
    wire N__42299;
    wire N__42294;
    wire N__42287;
    wire N__42284;
    wire N__42281;
    wire N__42278;
    wire N__42277;
    wire N__42274;
    wire N__42271;
    wire N__42266;
    wire N__42263;
    wire N__42262;
    wire N__42259;
    wire N__42258;
    wire N__42255;
    wire N__42252;
    wire N__42249;
    wire N__42242;
    wire N__42241;
    wire N__42236;
    wire N__42233;
    wire N__42232;
    wire N__42227;
    wire N__42224;
    wire N__42221;
    wire N__42220;
    wire N__42217;
    wire N__42216;
    wire N__42213;
    wire N__42210;
    wire N__42207;
    wire N__42200;
    wire N__42199;
    wire N__42194;
    wire N__42193;
    wire N__42192;
    wire N__42189;
    wire N__42186;
    wire N__42183;
    wire N__42180;
    wire N__42175;
    wire N__42170;
    wire N__42169;
    wire N__42166;
    wire N__42165;
    wire N__42164;
    wire N__42161;
    wire N__42158;
    wire N__42155;
    wire N__42152;
    wire N__42145;
    wire N__42142;
    wire N__42137;
    wire N__42134;
    wire N__42131;
    wire N__42128;
    wire N__42125;
    wire N__42122;
    wire N__42119;
    wire N__42116;
    wire N__42115;
    wire N__42112;
    wire N__42109;
    wire N__42104;
    wire N__42103;
    wire N__42102;
    wire N__42101;
    wire N__42098;
    wire N__42091;
    wire N__42086;
    wire N__42083;
    wire N__42080;
    wire N__42077;
    wire N__42076;
    wire N__42073;
    wire N__42072;
    wire N__42071;
    wire N__42066;
    wire N__42061;
    wire N__42058;
    wire N__42053;
    wire N__42050;
    wire N__42049;
    wire N__42046;
    wire N__42043;
    wire N__42038;
    wire N__42035;
    wire N__42032;
    wire N__42029;
    wire N__42026;
    wire N__42025;
    wire N__42020;
    wire N__42019;
    wire N__42016;
    wire N__42013;
    wire N__42010;
    wire N__42005;
    wire N__42004;
    wire N__42001;
    wire N__41998;
    wire N__41995;
    wire N__41992;
    wire N__41987;
    wire N__41986;
    wire N__41983;
    wire N__41980;
    wire N__41977;
    wire N__41972;
    wire N__41971;
    wire N__41968;
    wire N__41965;
    wire N__41960;
    wire N__41957;
    wire N__41954;
    wire N__41951;
    wire N__41948;
    wire N__41945;
    wire N__41944;
    wire N__41943;
    wire N__41942;
    wire N__41939;
    wire N__41936;
    wire N__41933;
    wire N__41930;
    wire N__41927;
    wire N__41924;
    wire N__41921;
    wire N__41914;
    wire N__41911;
    wire N__41906;
    wire N__41903;
    wire N__41902;
    wire N__41901;
    wire N__41900;
    wire N__41899;
    wire N__41898;
    wire N__41897;
    wire N__41896;
    wire N__41895;
    wire N__41894;
    wire N__41893;
    wire N__41892;
    wire N__41891;
    wire N__41890;
    wire N__41889;
    wire N__41888;
    wire N__41887;
    wire N__41886;
    wire N__41885;
    wire N__41884;
    wire N__41883;
    wire N__41882;
    wire N__41881;
    wire N__41880;
    wire N__41879;
    wire N__41878;
    wire N__41875;
    wire N__41868;
    wire N__41865;
    wire N__41862;
    wire N__41861;
    wire N__41860;
    wire N__41859;
    wire N__41858;
    wire N__41857;
    wire N__41856;
    wire N__41855;
    wire N__41854;
    wire N__41853;
    wire N__41852;
    wire N__41851;
    wire N__41850;
    wire N__41849;
    wire N__41844;
    wire N__41841;
    wire N__41834;
    wire N__41833;
    wire N__41832;
    wire N__41829;
    wire N__41826;
    wire N__41825;
    wire N__41822;
    wire N__41821;
    wire N__41820;
    wire N__41817;
    wire N__41816;
    wire N__41815;
    wire N__41814;
    wire N__41811;
    wire N__41806;
    wire N__41803;
    wire N__41796;
    wire N__41795;
    wire N__41794;
    wire N__41793;
    wire N__41792;
    wire N__41791;
    wire N__41790;
    wire N__41789;
    wire N__41788;
    wire N__41787;
    wire N__41786;
    wire N__41785;
    wire N__41784;
    wire N__41783;
    wire N__41782;
    wire N__41781;
    wire N__41780;
    wire N__41779;
    wire N__41776;
    wire N__41775;
    wire N__41774;
    wire N__41773;
    wire N__41772;
    wire N__41771;
    wire N__41770;
    wire N__41769;
    wire N__41768;
    wire N__41765;
    wire N__41762;
    wire N__41757;
    wire N__41752;
    wire N__41749;
    wire N__41744;
    wire N__41743;
    wire N__41742;
    wire N__41733;
    wire N__41728;
    wire N__41723;
    wire N__41718;
    wire N__41711;
    wire N__41706;
    wire N__41701;
    wire N__41698;
    wire N__41695;
    wire N__41690;
    wire N__41687;
    wire N__41684;
    wire N__41679;
    wire N__41676;
    wire N__41669;
    wire N__41668;
    wire N__41667;
    wire N__41666;
    wire N__41665;
    wire N__41664;
    wire N__41663;
    wire N__41662;
    wire N__41661;
    wire N__41660;
    wire N__41659;
    wire N__41658;
    wire N__41657;
    wire N__41656;
    wire N__41655;
    wire N__41654;
    wire N__41653;
    wire N__41652;
    wire N__41651;
    wire N__41648;
    wire N__41635;
    wire N__41628;
    wire N__41623;
    wire N__41620;
    wire N__41613;
    wire N__41610;
    wire N__41607;
    wire N__41596;
    wire N__41589;
    wire N__41584;
    wire N__41577;
    wire N__41574;
    wire N__41569;
    wire N__41562;
    wire N__41551;
    wire N__41548;
    wire N__41543;
    wire N__41534;
    wire N__41531;
    wire N__41524;
    wire N__41513;
    wire N__41500;
    wire N__41497;
    wire N__41492;
    wire N__41485;
    wire N__41482;
    wire N__41477;
    wire N__41474;
    wire N__41471;
    wire N__41462;
    wire N__41447;
    wire N__41420;
    wire N__41419;
    wire N__41416;
    wire N__41415;
    wire N__41412;
    wire N__41409;
    wire N__41406;
    wire N__41403;
    wire N__41400;
    wire N__41393;
    wire N__41390;
    wire N__41387;
    wire N__41386;
    wire N__41383;
    wire N__41380;
    wire N__41375;
    wire N__41372;
    wire N__41371;
    wire N__41368;
    wire N__41367;
    wire N__41364;
    wire N__41361;
    wire N__41358;
    wire N__41351;
    wire N__41350;
    wire N__41345;
    wire N__41342;
    wire N__41339;
    wire N__41338;
    wire N__41333;
    wire N__41330;
    wire N__41327;
    wire N__41324;
    wire N__41321;
    wire N__41318;
    wire N__41315;
    wire N__41314;
    wire N__41311;
    wire N__41308;
    wire N__41305;
    wire N__41304;
    wire N__41301;
    wire N__41298;
    wire N__41297;
    wire N__41294;
    wire N__41291;
    wire N__41288;
    wire N__41285;
    wire N__41280;
    wire N__41273;
    wire N__41270;
    wire N__41269;
    wire N__41266;
    wire N__41263;
    wire N__41260;
    wire N__41259;
    wire N__41258;
    wire N__41255;
    wire N__41252;
    wire N__41249;
    wire N__41246;
    wire N__41239;
    wire N__41234;
    wire N__41231;
    wire N__41228;
    wire N__41225;
    wire N__41224;
    wire N__41221;
    wire N__41218;
    wire N__41215;
    wire N__41212;
    wire N__41211;
    wire N__41208;
    wire N__41207;
    wire N__41204;
    wire N__41201;
    wire N__41198;
    wire N__41195;
    wire N__41192;
    wire N__41183;
    wire N__41180;
    wire N__41179;
    wire N__41176;
    wire N__41173;
    wire N__41170;
    wire N__41169;
    wire N__41168;
    wire N__41165;
    wire N__41162;
    wire N__41159;
    wire N__41156;
    wire N__41153;
    wire N__41144;
    wire N__41141;
    wire N__41140;
    wire N__41137;
    wire N__41136;
    wire N__41133;
    wire N__41130;
    wire N__41127;
    wire N__41124;
    wire N__41121;
    wire N__41120;
    wire N__41115;
    wire N__41112;
    wire N__41109;
    wire N__41106;
    wire N__41099;
    wire N__41096;
    wire N__41093;
    wire N__41092;
    wire N__41089;
    wire N__41088;
    wire N__41085;
    wire N__41082;
    wire N__41079;
    wire N__41078;
    wire N__41075;
    wire N__41072;
    wire N__41069;
    wire N__41066;
    wire N__41063;
    wire N__41054;
    wire N__41051;
    wire N__41050;
    wire N__41047;
    wire N__41046;
    wire N__41043;
    wire N__41042;
    wire N__41041;
    wire N__41040;
    wire N__41037;
    wire N__41036;
    wire N__41035;
    wire N__41034;
    wire N__41033;
    wire N__41032;
    wire N__41031;
    wire N__41028;
    wire N__41025;
    wire N__41022;
    wire N__41017;
    wire N__41014;
    wire N__41013;
    wire N__41012;
    wire N__41011;
    wire N__41010;
    wire N__41009;
    wire N__41008;
    wire N__41007;
    wire N__41006;
    wire N__41005;
    wire N__41004;
    wire N__41003;
    wire N__41002;
    wire N__41001;
    wire N__41000;
    wire N__40999;
    wire N__40998;
    wire N__40997;
    wire N__40996;
    wire N__40995;
    wire N__40992;
    wire N__40989;
    wire N__40980;
    wire N__40977;
    wire N__40972;
    wire N__40971;
    wire N__40968;
    wire N__40965;
    wire N__40962;
    wire N__40959;
    wire N__40956;
    wire N__40949;
    wire N__40946;
    wire N__40931;
    wire N__40920;
    wire N__40917;
    wire N__40908;
    wire N__40905;
    wire N__40898;
    wire N__40895;
    wire N__40874;
    wire N__40873;
    wire N__40872;
    wire N__40871;
    wire N__40870;
    wire N__40869;
    wire N__40868;
    wire N__40867;
    wire N__40866;
    wire N__40863;
    wire N__40862;
    wire N__40859;
    wire N__40858;
    wire N__40855;
    wire N__40854;
    wire N__40851;
    wire N__40850;
    wire N__40847;
    wire N__40846;
    wire N__40843;
    wire N__40842;
    wire N__40839;
    wire N__40838;
    wire N__40837;
    wire N__40834;
    wire N__40833;
    wire N__40818;
    wire N__40801;
    wire N__40794;
    wire N__40787;
    wire N__40784;
    wire N__40781;
    wire N__40778;
    wire N__40775;
    wire N__40774;
    wire N__40771;
    wire N__40768;
    wire N__40763;
    wire N__40760;
    wire N__40759;
    wire N__40756;
    wire N__40753;
    wire N__40750;
    wire N__40749;
    wire N__40744;
    wire N__40741;
    wire N__40736;
    wire N__40735;
    wire N__40732;
    wire N__40729;
    wire N__40726;
    wire N__40725;
    wire N__40722;
    wire N__40719;
    wire N__40716;
    wire N__40713;
    wire N__40710;
    wire N__40709;
    wire N__40706;
    wire N__40703;
    wire N__40700;
    wire N__40697;
    wire N__40694;
    wire N__40691;
    wire N__40688;
    wire N__40683;
    wire N__40676;
    wire N__40673;
    wire N__40670;
    wire N__40669;
    wire N__40666;
    wire N__40665;
    wire N__40662;
    wire N__40661;
    wire N__40658;
    wire N__40655;
    wire N__40652;
    wire N__40649;
    wire N__40646;
    wire N__40643;
    wire N__40640;
    wire N__40637;
    wire N__40628;
    wire N__40625;
    wire N__40622;
    wire N__40619;
    wire N__40616;
    wire N__40615;
    wire N__40614;
    wire N__40611;
    wire N__40608;
    wire N__40605;
    wire N__40604;
    wire N__40599;
    wire N__40596;
    wire N__40593;
    wire N__40590;
    wire N__40587;
    wire N__40580;
    wire N__40577;
    wire N__40574;
    wire N__40573;
    wire N__40570;
    wire N__40567;
    wire N__40564;
    wire N__40561;
    wire N__40560;
    wire N__40557;
    wire N__40554;
    wire N__40551;
    wire N__40550;
    wire N__40543;
    wire N__40540;
    wire N__40537;
    wire N__40532;
    wire N__40529;
    wire N__40528;
    wire N__40525;
    wire N__40522;
    wire N__40519;
    wire N__40516;
    wire N__40515;
    wire N__40514;
    wire N__40511;
    wire N__40508;
    wire N__40505;
    wire N__40502;
    wire N__40499;
    wire N__40494;
    wire N__40487;
    wire N__40484;
    wire N__40481;
    wire N__40478;
    wire N__40477;
    wire N__40474;
    wire N__40473;
    wire N__40470;
    wire N__40469;
    wire N__40466;
    wire N__40463;
    wire N__40460;
    wire N__40457;
    wire N__40454;
    wire N__40451;
    wire N__40448;
    wire N__40439;
    wire N__40436;
    wire N__40433;
    wire N__40430;
    wire N__40427;
    wire N__40424;
    wire N__40421;
    wire N__40420;
    wire N__40417;
    wire N__40414;
    wire N__40413;
    wire N__40412;
    wire N__40407;
    wire N__40404;
    wire N__40401;
    wire N__40396;
    wire N__40391;
    wire N__40388;
    wire N__40385;
    wire N__40384;
    wire N__40383;
    wire N__40380;
    wire N__40379;
    wire N__40376;
    wire N__40373;
    wire N__40370;
    wire N__40367;
    wire N__40362;
    wire N__40359;
    wire N__40356;
    wire N__40353;
    wire N__40346;
    wire N__40343;
    wire N__40340;
    wire N__40337;
    wire N__40334;
    wire N__40331;
    wire N__40328;
    wire N__40327;
    wire N__40324;
    wire N__40323;
    wire N__40320;
    wire N__40317;
    wire N__40314;
    wire N__40311;
    wire N__40308;
    wire N__40303;
    wire N__40302;
    wire N__40299;
    wire N__40296;
    wire N__40293;
    wire N__40290;
    wire N__40283;
    wire N__40280;
    wire N__40277;
    wire N__40274;
    wire N__40271;
    wire N__40268;
    wire N__40265;
    wire N__40262;
    wire N__40261;
    wire N__40258;
    wire N__40255;
    wire N__40254;
    wire N__40251;
    wire N__40250;
    wire N__40247;
    wire N__40244;
    wire N__40241;
    wire N__40238;
    wire N__40235;
    wire N__40232;
    wire N__40229;
    wire N__40222;
    wire N__40217;
    wire N__40214;
    wire N__40211;
    wire N__40208;
    wire N__40205;
    wire N__40202;
    wire N__40199;
    wire N__40198;
    wire N__40195;
    wire N__40194;
    wire N__40191;
    wire N__40188;
    wire N__40185;
    wire N__40182;
    wire N__40181;
    wire N__40178;
    wire N__40175;
    wire N__40172;
    wire N__40169;
    wire N__40166;
    wire N__40161;
    wire N__40158;
    wire N__40151;
    wire N__40148;
    wire N__40145;
    wire N__40142;
    wire N__40139;
    wire N__40136;
    wire N__40133;
    wire N__40130;
    wire N__40129;
    wire N__40128;
    wire N__40125;
    wire N__40122;
    wire N__40119;
    wire N__40118;
    wire N__40115;
    wire N__40112;
    wire N__40109;
    wire N__40106;
    wire N__40103;
    wire N__40098;
    wire N__40095;
    wire N__40092;
    wire N__40085;
    wire N__40082;
    wire N__40081;
    wire N__40080;
    wire N__40077;
    wire N__40074;
    wire N__40071;
    wire N__40068;
    wire N__40067;
    wire N__40064;
    wire N__40061;
    wire N__40058;
    wire N__40055;
    wire N__40050;
    wire N__40043;
    wire N__40040;
    wire N__40037;
    wire N__40034;
    wire N__40031;
    wire N__40028;
    wire N__40025;
    wire N__40022;
    wire N__40021;
    wire N__40020;
    wire N__40017;
    wire N__40016;
    wire N__40013;
    wire N__40010;
    wire N__40007;
    wire N__40004;
    wire N__40001;
    wire N__39994;
    wire N__39991;
    wire N__39986;
    wire N__39983;
    wire N__39980;
    wire N__39979;
    wire N__39976;
    wire N__39973;
    wire N__39970;
    wire N__39967;
    wire N__39966;
    wire N__39965;
    wire N__39962;
    wire N__39959;
    wire N__39956;
    wire N__39953;
    wire N__39946;
    wire N__39941;
    wire N__39938;
    wire N__39935;
    wire N__39932;
    wire N__39929;
    wire N__39926;
    wire N__39925;
    wire N__39922;
    wire N__39921;
    wire N__39920;
    wire N__39917;
    wire N__39914;
    wire N__39911;
    wire N__39908;
    wire N__39901;
    wire N__39896;
    wire N__39893;
    wire N__39892;
    wire N__39889;
    wire N__39886;
    wire N__39881;
    wire N__39878;
    wire N__39877;
    wire N__39874;
    wire N__39873;
    wire N__39870;
    wire N__39867;
    wire N__39864;
    wire N__39861;
    wire N__39858;
    wire N__39857;
    wire N__39854;
    wire N__39851;
    wire N__39848;
    wire N__39845;
    wire N__39842;
    wire N__39839;
    wire N__39836;
    wire N__39835;
    wire N__39832;
    wire N__39825;
    wire N__39822;
    wire N__39819;
    wire N__39816;
    wire N__39809;
    wire N__39806;
    wire N__39803;
    wire N__39800;
    wire N__39797;
    wire N__39796;
    wire N__39793;
    wire N__39790;
    wire N__39787;
    wire N__39786;
    wire N__39781;
    wire N__39778;
    wire N__39773;
    wire N__39770;
    wire N__39767;
    wire N__39764;
    wire N__39761;
    wire N__39758;
    wire N__39755;
    wire N__39752;
    wire N__39749;
    wire N__39748;
    wire N__39747;
    wire N__39744;
    wire N__39741;
    wire N__39738;
    wire N__39735;
    wire N__39730;
    wire N__39729;
    wire N__39726;
    wire N__39723;
    wire N__39720;
    wire N__39717;
    wire N__39710;
    wire N__39707;
    wire N__39704;
    wire N__39701;
    wire N__39698;
    wire N__39695;
    wire N__39694;
    wire N__39691;
    wire N__39690;
    wire N__39687;
    wire N__39684;
    wire N__39681;
    wire N__39678;
    wire N__39675;
    wire N__39670;
    wire N__39667;
    wire N__39666;
    wire N__39661;
    wire N__39658;
    wire N__39655;
    wire N__39650;
    wire N__39647;
    wire N__39646;
    wire N__39645;
    wire N__39642;
    wire N__39639;
    wire N__39638;
    wire N__39635;
    wire N__39632;
    wire N__39629;
    wire N__39626;
    wire N__39621;
    wire N__39618;
    wire N__39615;
    wire N__39612;
    wire N__39605;
    wire N__39602;
    wire N__39599;
    wire N__39596;
    wire N__39593;
    wire N__39590;
    wire N__39587;
    wire N__39584;
    wire N__39581;
    wire N__39580;
    wire N__39577;
    wire N__39574;
    wire N__39573;
    wire N__39570;
    wire N__39567;
    wire N__39564;
    wire N__39561;
    wire N__39558;
    wire N__39557;
    wire N__39550;
    wire N__39547;
    wire N__39542;
    wire N__39539;
    wire N__39536;
    wire N__39533;
    wire N__39530;
    wire N__39527;
    wire N__39524;
    wire N__39523;
    wire N__39520;
    wire N__39519;
    wire N__39516;
    wire N__39513;
    wire N__39512;
    wire N__39509;
    wire N__39506;
    wire N__39503;
    wire N__39500;
    wire N__39495;
    wire N__39488;
    wire N__39485;
    wire N__39482;
    wire N__39479;
    wire N__39476;
    wire N__39473;
    wire N__39472;
    wire N__39471;
    wire N__39468;
    wire N__39465;
    wire N__39462;
    wire N__39459;
    wire N__39458;
    wire N__39453;
    wire N__39450;
    wire N__39447;
    wire N__39444;
    wire N__39437;
    wire N__39434;
    wire N__39433;
    wire N__39430;
    wire N__39427;
    wire N__39422;
    wire N__39419;
    wire N__39418;
    wire N__39417;
    wire N__39414;
    wire N__39411;
    wire N__39408;
    wire N__39401;
    wire N__39398;
    wire N__39395;
    wire N__39392;
    wire N__39389;
    wire N__39388;
    wire N__39385;
    wire N__39382;
    wire N__39379;
    wire N__39376;
    wire N__39373;
    wire N__39370;
    wire N__39367;
    wire N__39362;
    wire N__39359;
    wire N__39356;
    wire N__39353;
    wire N__39352;
    wire N__39351;
    wire N__39348;
    wire N__39345;
    wire N__39342;
    wire N__39335;
    wire N__39334;
    wire N__39333;
    wire N__39332;
    wire N__39329;
    wire N__39324;
    wire N__39321;
    wire N__39318;
    wire N__39311;
    wire N__39310;
    wire N__39309;
    wire N__39308;
    wire N__39307;
    wire N__39306;
    wire N__39303;
    wire N__39300;
    wire N__39295;
    wire N__39294;
    wire N__39289;
    wire N__39282;
    wire N__39279;
    wire N__39272;
    wire N__39269;
    wire N__39266;
    wire N__39263;
    wire N__39260;
    wire N__39259;
    wire N__39256;
    wire N__39253;
    wire N__39248;
    wire N__39245;
    wire N__39244;
    wire N__39243;
    wire N__39240;
    wire N__39237;
    wire N__39234;
    wire N__39227;
    wire N__39224;
    wire N__39221;
    wire N__39220;
    wire N__39219;
    wire N__39216;
    wire N__39213;
    wire N__39210;
    wire N__39203;
    wire N__39200;
    wire N__39197;
    wire N__39196;
    wire N__39195;
    wire N__39192;
    wire N__39189;
    wire N__39186;
    wire N__39179;
    wire N__39176;
    wire N__39173;
    wire N__39172;
    wire N__39171;
    wire N__39168;
    wire N__39165;
    wire N__39162;
    wire N__39155;
    wire N__39152;
    wire N__39149;
    wire N__39148;
    wire N__39147;
    wire N__39144;
    wire N__39141;
    wire N__39138;
    wire N__39131;
    wire N__39128;
    wire N__39125;
    wire N__39124;
    wire N__39123;
    wire N__39120;
    wire N__39117;
    wire N__39114;
    wire N__39107;
    wire N__39104;
    wire N__39101;
    wire N__39100;
    wire N__39099;
    wire N__39096;
    wire N__39093;
    wire N__39090;
    wire N__39083;
    wire N__39080;
    wire N__39077;
    wire N__39076;
    wire N__39075;
    wire N__39072;
    wire N__39069;
    wire N__39066;
    wire N__39059;
    wire N__39056;
    wire N__39055;
    wire N__39054;
    wire N__39051;
    wire N__39046;
    wire N__39041;
    wire N__39040;
    wire N__39037;
    wire N__39034;
    wire N__39031;
    wire N__39026;
    wire N__39023;
    wire N__39022;
    wire N__39021;
    wire N__39018;
    wire N__39013;
    wire N__39008;
    wire N__39005;
    wire N__39002;
    wire N__39001;
    wire N__39000;
    wire N__38997;
    wire N__38994;
    wire N__38991;
    wire N__38984;
    wire N__38981;
    wire N__38980;
    wire N__38979;
    wire N__38976;
    wire N__38973;
    wire N__38970;
    wire N__38965;
    wire N__38960;
    wire N__38957;
    wire N__38954;
    wire N__38953;
    wire N__38952;
    wire N__38949;
    wire N__38946;
    wire N__38943;
    wire N__38936;
    wire N__38933;
    wire N__38930;
    wire N__38929;
    wire N__38928;
    wire N__38925;
    wire N__38922;
    wire N__38919;
    wire N__38912;
    wire N__38909;
    wire N__38906;
    wire N__38905;
    wire N__38904;
    wire N__38901;
    wire N__38898;
    wire N__38895;
    wire N__38888;
    wire N__38885;
    wire N__38882;
    wire N__38881;
    wire N__38880;
    wire N__38877;
    wire N__38874;
    wire N__38871;
    wire N__38864;
    wire N__38861;
    wire N__38858;
    wire N__38857;
    wire N__38856;
    wire N__38853;
    wire N__38850;
    wire N__38847;
    wire N__38840;
    wire N__38837;
    wire N__38834;
    wire N__38833;
    wire N__38832;
    wire N__38829;
    wire N__38826;
    wire N__38823;
    wire N__38816;
    wire N__38813;
    wire N__38810;
    wire N__38809;
    wire N__38808;
    wire N__38805;
    wire N__38802;
    wire N__38799;
    wire N__38792;
    wire N__38789;
    wire N__38786;
    wire N__38785;
    wire N__38784;
    wire N__38781;
    wire N__38778;
    wire N__38775;
    wire N__38768;
    wire N__38765;
    wire N__38762;
    wire N__38761;
    wire N__38760;
    wire N__38757;
    wire N__38754;
    wire N__38751;
    wire N__38744;
    wire N__38741;
    wire N__38738;
    wire N__38737;
    wire N__38736;
    wire N__38733;
    wire N__38730;
    wire N__38727;
    wire N__38720;
    wire N__38717;
    wire N__38714;
    wire N__38713;
    wire N__38712;
    wire N__38709;
    wire N__38706;
    wire N__38703;
    wire N__38696;
    wire N__38693;
    wire N__38690;
    wire N__38689;
    wire N__38688;
    wire N__38685;
    wire N__38682;
    wire N__38679;
    wire N__38672;
    wire N__38669;
    wire N__38666;
    wire N__38665;
    wire N__38664;
    wire N__38661;
    wire N__38658;
    wire N__38655;
    wire N__38648;
    wire N__38645;
    wire N__38642;
    wire N__38641;
    wire N__38636;
    wire N__38633;
    wire N__38630;
    wire N__38627;
    wire N__38624;
    wire N__38621;
    wire N__38618;
    wire N__38615;
    wire N__38612;
    wire N__38609;
    wire N__38606;
    wire N__38605;
    wire N__38600;
    wire N__38597;
    wire N__38594;
    wire N__38591;
    wire N__38588;
    wire N__38585;
    wire N__38584;
    wire N__38581;
    wire N__38578;
    wire N__38573;
    wire N__38570;
    wire N__38569;
    wire N__38566;
    wire N__38563;
    wire N__38562;
    wire N__38559;
    wire N__38556;
    wire N__38553;
    wire N__38546;
    wire N__38543;
    wire N__38542;
    wire N__38539;
    wire N__38536;
    wire N__38535;
    wire N__38532;
    wire N__38529;
    wire N__38526;
    wire N__38519;
    wire N__38516;
    wire N__38513;
    wire N__38510;
    wire N__38507;
    wire N__38504;
    wire N__38503;
    wire N__38502;
    wire N__38499;
    wire N__38496;
    wire N__38491;
    wire N__38486;
    wire N__38485;
    wire N__38484;
    wire N__38481;
    wire N__38478;
    wire N__38473;
    wire N__38468;
    wire N__38465;
    wire N__38462;
    wire N__38459;
    wire N__38456;
    wire N__38453;
    wire N__38452;
    wire N__38447;
    wire N__38444;
    wire N__38443;
    wire N__38438;
    wire N__38435;
    wire N__38432;
    wire N__38429;
    wire N__38426;
    wire N__38423;
    wire N__38420;
    wire N__38417;
    wire N__38414;
    wire N__38411;
    wire N__38408;
    wire N__38407;
    wire N__38406;
    wire N__38403;
    wire N__38400;
    wire N__38397;
    wire N__38390;
    wire N__38389;
    wire N__38386;
    wire N__38385;
    wire N__38382;
    wire N__38379;
    wire N__38376;
    wire N__38369;
    wire N__38366;
    wire N__38363;
    wire N__38360;
    wire N__38359;
    wire N__38354;
    wire N__38351;
    wire N__38348;
    wire N__38345;
    wire N__38342;
    wire N__38339;
    wire N__38336;
    wire N__38333;
    wire N__38330;
    wire N__38327;
    wire N__38324;
    wire N__38321;
    wire N__38320;
    wire N__38315;
    wire N__38314;
    wire N__38311;
    wire N__38308;
    wire N__38305;
    wire N__38300;
    wire N__38297;
    wire N__38296;
    wire N__38291;
    wire N__38290;
    wire N__38287;
    wire N__38284;
    wire N__38281;
    wire N__38276;
    wire N__38273;
    wire N__38270;
    wire N__38267;
    wire N__38264;
    wire N__38261;
    wire N__38260;
    wire N__38257;
    wire N__38256;
    wire N__38253;
    wire N__38250;
    wire N__38249;
    wire N__38246;
    wire N__38243;
    wire N__38240;
    wire N__38237;
    wire N__38234;
    wire N__38231;
    wire N__38228;
    wire N__38225;
    wire N__38222;
    wire N__38219;
    wire N__38216;
    wire N__38213;
    wire N__38204;
    wire N__38201;
    wire N__38200;
    wire N__38197;
    wire N__38196;
    wire N__38193;
    wire N__38190;
    wire N__38187;
    wire N__38184;
    wire N__38181;
    wire N__38176;
    wire N__38171;
    wire N__38168;
    wire N__38165;
    wire N__38162;
    wire N__38159;
    wire N__38156;
    wire N__38153;
    wire N__38150;
    wire N__38147;
    wire N__38144;
    wire N__38141;
    wire N__38138;
    wire N__38135;
    wire N__38134;
    wire N__38129;
    wire N__38128;
    wire N__38125;
    wire N__38122;
    wire N__38119;
    wire N__38114;
    wire N__38113;
    wire N__38110;
    wire N__38105;
    wire N__38102;
    wire N__38099;
    wire N__38096;
    wire N__38093;
    wire N__38092;
    wire N__38089;
    wire N__38084;
    wire N__38083;
    wire N__38080;
    wire N__38077;
    wire N__38074;
    wire N__38069;
    wire N__38066;
    wire N__38063;
    wire N__38060;
    wire N__38057;
    wire N__38054;
    wire N__38051;
    wire N__38048;
    wire N__38045;
    wire N__38042;
    wire N__38039;
    wire N__38036;
    wire N__38033;
    wire N__38030;
    wire N__38027;
    wire N__38024;
    wire N__38021;
    wire N__38018;
    wire N__38015;
    wire N__38012;
    wire N__38009;
    wire N__38006;
    wire N__38003;
    wire N__38000;
    wire N__37997;
    wire N__37994;
    wire N__37991;
    wire N__37988;
    wire N__37985;
    wire N__37982;
    wire N__37979;
    wire N__37978;
    wire N__37975;
    wire N__37972;
    wire N__37967;
    wire N__37964;
    wire N__37961;
    wire N__37958;
    wire N__37955;
    wire N__37952;
    wire N__37949;
    wire N__37948;
    wire N__37945;
    wire N__37942;
    wire N__37937;
    wire N__37934;
    wire N__37931;
    wire N__37928;
    wire N__37927;
    wire N__37924;
    wire N__37921;
    wire N__37916;
    wire N__37913;
    wire N__37910;
    wire N__37909;
    wire N__37908;
    wire N__37907;
    wire N__37906;
    wire N__37905;
    wire N__37904;
    wire N__37903;
    wire N__37902;
    wire N__37901;
    wire N__37900;
    wire N__37899;
    wire N__37898;
    wire N__37895;
    wire N__37892;
    wire N__37891;
    wire N__37890;
    wire N__37889;
    wire N__37888;
    wire N__37887;
    wire N__37886;
    wire N__37885;
    wire N__37884;
    wire N__37883;
    wire N__37882;
    wire N__37881;
    wire N__37880;
    wire N__37879;
    wire N__37878;
    wire N__37875;
    wire N__37874;
    wire N__37871;
    wire N__37870;
    wire N__37867;
    wire N__37866;
    wire N__37865;
    wire N__37862;
    wire N__37861;
    wire N__37858;
    wire N__37857;
    wire N__37854;
    wire N__37853;
    wire N__37850;
    wire N__37847;
    wire N__37846;
    wire N__37843;
    wire N__37842;
    wire N__37839;
    wire N__37838;
    wire N__37835;
    wire N__37834;
    wire N__37833;
    wire N__37832;
    wire N__37831;
    wire N__37826;
    wire N__37819;
    wire N__37810;
    wire N__37807;
    wire N__37802;
    wire N__37799;
    wire N__37798;
    wire N__37797;
    wire N__37796;
    wire N__37795;
    wire N__37794;
    wire N__37793;
    wire N__37792;
    wire N__37791;
    wire N__37790;
    wire N__37789;
    wire N__37788;
    wire N__37787;
    wire N__37786;
    wire N__37785;
    wire N__37784;
    wire N__37779;
    wire N__37764;
    wire N__37747;
    wire N__37730;
    wire N__37729;
    wire N__37726;
    wire N__37725;
    wire N__37722;
    wire N__37721;
    wire N__37718;
    wire N__37717;
    wire N__37716;
    wire N__37709;
    wire N__37702;
    wire N__37699;
    wire N__37694;
    wire N__37691;
    wire N__37688;
    wire N__37685;
    wire N__37682;
    wire N__37679;
    wire N__37672;
    wire N__37663;
    wire N__37660;
    wire N__37655;
    wire N__37652;
    wire N__37637;
    wire N__37636;
    wire N__37633;
    wire N__37632;
    wire N__37629;
    wire N__37620;
    wire N__37607;
    wire N__37604;
    wire N__37601;
    wire N__37596;
    wire N__37589;
    wire N__37586;
    wire N__37581;
    wire N__37578;
    wire N__37573;
    wire N__37570;
    wire N__37565;
    wire N__37562;
    wire N__37559;
    wire N__37556;
    wire N__37547;
    wire N__37544;
    wire N__37541;
    wire N__37538;
    wire N__37535;
    wire N__37534;
    wire N__37531;
    wire N__37528;
    wire N__37523;
    wire N__37520;
    wire N__37517;
    wire N__37514;
    wire N__37511;
    wire N__37508;
    wire N__37505;
    wire N__37502;
    wire N__37499;
    wire N__37496;
    wire N__37493;
    wire N__37490;
    wire N__37487;
    wire N__37484;
    wire N__37481;
    wire N__37478;
    wire N__37475;
    wire N__37472;
    wire N__37469;
    wire N__37468;
    wire N__37467;
    wire N__37464;
    wire N__37459;
    wire N__37454;
    wire N__37453;
    wire N__37452;
    wire N__37449;
    wire N__37444;
    wire N__37439;
    wire N__37438;
    wire N__37435;
    wire N__37434;
    wire N__37431;
    wire N__37428;
    wire N__37425;
    wire N__37418;
    wire N__37417;
    wire N__37414;
    wire N__37413;
    wire N__37410;
    wire N__37407;
    wire N__37404;
    wire N__37397;
    wire N__37394;
    wire N__37393;
    wire N__37390;
    wire N__37387;
    wire N__37382;
    wire N__37379;
    wire N__37376;
    wire N__37373;
    wire N__37370;
    wire N__37367;
    wire N__37364;
    wire N__37361;
    wire N__37358;
    wire N__37355;
    wire N__37354;
    wire N__37351;
    wire N__37348;
    wire N__37343;
    wire N__37340;
    wire N__37337;
    wire N__37334;
    wire N__37331;
    wire N__37328;
    wire N__37325;
    wire N__37322;
    wire N__37319;
    wire N__37316;
    wire N__37313;
    wire N__37310;
    wire N__37309;
    wire N__37308;
    wire N__37307;
    wire N__37306;
    wire N__37305;
    wire N__37302;
    wire N__37299;
    wire N__37298;
    wire N__37297;
    wire N__37296;
    wire N__37295;
    wire N__37292;
    wire N__37289;
    wire N__37288;
    wire N__37285;
    wire N__37284;
    wire N__37281;
    wire N__37278;
    wire N__37273;
    wire N__37268;
    wire N__37265;
    wire N__37262;
    wire N__37253;
    wire N__37246;
    wire N__37241;
    wire N__37238;
    wire N__37235;
    wire N__37230;
    wire N__37223;
    wire N__37220;
    wire N__37217;
    wire N__37214;
    wire N__37211;
    wire N__37208;
    wire N__37205;
    wire N__37202;
    wire N__37199;
    wire N__37196;
    wire N__37193;
    wire N__37190;
    wire N__37187;
    wire N__37184;
    wire N__37181;
    wire N__37178;
    wire N__37175;
    wire N__37174;
    wire N__37171;
    wire N__37170;
    wire N__37167;
    wire N__37164;
    wire N__37161;
    wire N__37154;
    wire N__37151;
    wire N__37148;
    wire N__37145;
    wire N__37142;
    wire N__37139;
    wire N__37136;
    wire N__37133;
    wire N__37130;
    wire N__37127;
    wire N__37124;
    wire N__37121;
    wire N__37118;
    wire N__37115;
    wire N__37112;
    wire N__37109;
    wire N__37106;
    wire N__37103;
    wire N__37100;
    wire N__37097;
    wire N__37094;
    wire N__37091;
    wire N__37088;
    wire N__37085;
    wire N__37082;
    wire N__37079;
    wire N__37076;
    wire N__37073;
    wire N__37070;
    wire N__37067;
    wire N__37064;
    wire N__37061;
    wire N__37058;
    wire N__37055;
    wire N__37052;
    wire N__37049;
    wire N__37046;
    wire N__37043;
    wire N__37040;
    wire N__37037;
    wire N__37034;
    wire N__37031;
    wire N__37028;
    wire N__37025;
    wire N__37022;
    wire N__37019;
    wire N__37016;
    wire N__37013;
    wire N__37010;
    wire N__37007;
    wire N__37004;
    wire N__37001;
    wire N__36998;
    wire N__36995;
    wire N__36992;
    wire N__36989;
    wire N__36986;
    wire N__36983;
    wire N__36980;
    wire N__36977;
    wire N__36974;
    wire N__36971;
    wire N__36968;
    wire N__36965;
    wire N__36962;
    wire N__36959;
    wire N__36958;
    wire N__36955;
    wire N__36954;
    wire N__36951;
    wire N__36948;
    wire N__36945;
    wire N__36938;
    wire N__36935;
    wire N__36932;
    wire N__36931;
    wire N__36928;
    wire N__36925;
    wire N__36922;
    wire N__36919;
    wire N__36916;
    wire N__36913;
    wire N__36908;
    wire N__36905;
    wire N__36902;
    wire N__36901;
    wire N__36898;
    wire N__36895;
    wire N__36892;
    wire N__36889;
    wire N__36886;
    wire N__36883;
    wire N__36880;
    wire N__36877;
    wire N__36872;
    wire N__36869;
    wire N__36868;
    wire N__36867;
    wire N__36866;
    wire N__36861;
    wire N__36858;
    wire N__36855;
    wire N__36848;
    wire N__36847;
    wire N__36846;
    wire N__36845;
    wire N__36842;
    wire N__36835;
    wire N__36830;
    wire N__36829;
    wire N__36826;
    wire N__36823;
    wire N__36820;
    wire N__36817;
    wire N__36814;
    wire N__36811;
    wire N__36808;
    wire N__36803;
    wire N__36800;
    wire N__36797;
    wire N__36794;
    wire N__36791;
    wire N__36788;
    wire N__36785;
    wire N__36782;
    wire N__36779;
    wire N__36776;
    wire N__36773;
    wire N__36770;
    wire N__36767;
    wire N__36764;
    wire N__36761;
    wire N__36758;
    wire N__36755;
    wire N__36752;
    wire N__36749;
    wire N__36746;
    wire N__36743;
    wire N__36740;
    wire N__36737;
    wire N__36734;
    wire N__36731;
    wire N__36728;
    wire N__36727;
    wire N__36726;
    wire N__36725;
    wire N__36724;
    wire N__36723;
    wire N__36722;
    wire N__36721;
    wire N__36720;
    wire N__36719;
    wire N__36718;
    wire N__36717;
    wire N__36716;
    wire N__36715;
    wire N__36714;
    wire N__36713;
    wire N__36712;
    wire N__36711;
    wire N__36710;
    wire N__36709;
    wire N__36708;
    wire N__36707;
    wire N__36706;
    wire N__36705;
    wire N__36704;
    wire N__36703;
    wire N__36702;
    wire N__36701;
    wire N__36700;
    wire N__36699;
    wire N__36690;
    wire N__36681;
    wire N__36672;
    wire N__36663;
    wire N__36654;
    wire N__36649;
    wire N__36640;
    wire N__36631;
    wire N__36626;
    wire N__36619;
    wire N__36608;
    wire N__36607;
    wire N__36606;
    wire N__36605;
    wire N__36602;
    wire N__36601;
    wire N__36598;
    wire N__36597;
    wire N__36596;
    wire N__36595;
    wire N__36594;
    wire N__36593;
    wire N__36590;
    wire N__36587;
    wire N__36584;
    wire N__36581;
    wire N__36580;
    wire N__36579;
    wire N__36578;
    wire N__36577;
    wire N__36576;
    wire N__36575;
    wire N__36574;
    wire N__36573;
    wire N__36572;
    wire N__36571;
    wire N__36570;
    wire N__36569;
    wire N__36568;
    wire N__36567;
    wire N__36566;
    wire N__36565;
    wire N__36564;
    wire N__36563;
    wire N__36562;
    wire N__36561;
    wire N__36560;
    wire N__36559;
    wire N__36558;
    wire N__36555;
    wire N__36552;
    wire N__36549;
    wire N__36548;
    wire N__36547;
    wire N__36546;
    wire N__36545;
    wire N__36544;
    wire N__36543;
    wire N__36542;
    wire N__36539;
    wire N__36538;
    wire N__36535;
    wire N__36532;
    wire N__36531;
    wire N__36522;
    wire N__36513;
    wire N__36506;
    wire N__36497;
    wire N__36488;
    wire N__36479;
    wire N__36470;
    wire N__36469;
    wire N__36464;
    wire N__36461;
    wire N__36454;
    wire N__36445;
    wire N__36444;
    wire N__36441;
    wire N__36438;
    wire N__36435;
    wire N__36432;
    wire N__36429;
    wire N__36426;
    wire N__36417;
    wire N__36412;
    wire N__36409;
    wire N__36404;
    wire N__36399;
    wire N__36396;
    wire N__36393;
    wire N__36386;
    wire N__36383;
    wire N__36380;
    wire N__36375;
    wire N__36372;
    wire N__36367;
    wire N__36364;
    wire N__36357;
    wire N__36354;
    wire N__36351;
    wire N__36346;
    wire N__36341;
    wire N__36338;
    wire N__36335;
    wire N__36332;
    wire N__36323;
    wire N__36320;
    wire N__36317;
    wire N__36316;
    wire N__36313;
    wire N__36310;
    wire N__36307;
    wire N__36304;
    wire N__36301;
    wire N__36298;
    wire N__36293;
    wire N__36290;
    wire N__36287;
    wire N__36284;
    wire N__36283;
    wire N__36280;
    wire N__36277;
    wire N__36274;
    wire N__36269;
    wire N__36266;
    wire N__36263;
    wire N__36260;
    wire N__36257;
    wire N__36254;
    wire N__36251;
    wire N__36248;
    wire N__36245;
    wire N__36242;
    wire N__36239;
    wire N__36236;
    wire N__36233;
    wire N__36230;
    wire N__36227;
    wire N__36224;
    wire N__36221;
    wire N__36218;
    wire N__36215;
    wire N__36214;
    wire N__36213;
    wire N__36212;
    wire N__36209;
    wire N__36202;
    wire N__36197;
    wire N__36194;
    wire N__36193;
    wire N__36192;
    wire N__36191;
    wire N__36190;
    wire N__36189;
    wire N__36188;
    wire N__36187;
    wire N__36186;
    wire N__36185;
    wire N__36184;
    wire N__36183;
    wire N__36182;
    wire N__36181;
    wire N__36180;
    wire N__36179;
    wire N__36178;
    wire N__36177;
    wire N__36176;
    wire N__36175;
    wire N__36174;
    wire N__36173;
    wire N__36172;
    wire N__36171;
    wire N__36170;
    wire N__36169;
    wire N__36160;
    wire N__36151;
    wire N__36142;
    wire N__36135;
    wire N__36126;
    wire N__36125;
    wire N__36124;
    wire N__36123;
    wire N__36122;
    wire N__36121;
    wire N__36120;
    wire N__36113;
    wire N__36104;
    wire N__36093;
    wire N__36090;
    wire N__36081;
    wire N__36078;
    wire N__36071;
    wire N__36068;
    wire N__36065;
    wire N__36060;
    wire N__36057;
    wire N__36050;
    wire N__36047;
    wire N__36046;
    wire N__36045;
    wire N__36042;
    wire N__36041;
    wire N__36038;
    wire N__36035;
    wire N__36028;
    wire N__36023;
    wire N__36020;
    wire N__36017;
    wire N__36014;
    wire N__36011;
    wire N__36008;
    wire N__36005;
    wire N__36002;
    wire N__35999;
    wire N__35996;
    wire N__35993;
    wire N__35990;
    wire N__35987;
    wire N__35984;
    wire N__35983;
    wire N__35982;
    wire N__35979;
    wire N__35976;
    wire N__35971;
    wire N__35966;
    wire N__35963;
    wire N__35962;
    wire N__35959;
    wire N__35958;
    wire N__35955;
    wire N__35952;
    wire N__35949;
    wire N__35942;
    wire N__35939;
    wire N__35938;
    wire N__35935;
    wire N__35932;
    wire N__35929;
    wire N__35924;
    wire N__35921;
    wire N__35920;
    wire N__35917;
    wire N__35914;
    wire N__35911;
    wire N__35906;
    wire N__35903;
    wire N__35902;
    wire N__35899;
    wire N__35896;
    wire N__35893;
    wire N__35888;
    wire N__35885;
    wire N__35884;
    wire N__35883;
    wire N__35880;
    wire N__35877;
    wire N__35872;
    wire N__35867;
    wire N__35864;
    wire N__35863;
    wire N__35862;
    wire N__35859;
    wire N__35856;
    wire N__35853;
    wire N__35846;
    wire N__35843;
    wire N__35840;
    wire N__35837;
    wire N__35834;
    wire N__35831;
    wire N__35828;
    wire N__35825;
    wire N__35824;
    wire N__35821;
    wire N__35818;
    wire N__35815;
    wire N__35810;
    wire N__35807;
    wire N__35806;
    wire N__35803;
    wire N__35800;
    wire N__35797;
    wire N__35792;
    wire N__35789;
    wire N__35788;
    wire N__35785;
    wire N__35782;
    wire N__35779;
    wire N__35774;
    wire N__35771;
    wire N__35770;
    wire N__35767;
    wire N__35764;
    wire N__35761;
    wire N__35756;
    wire N__35753;
    wire N__35752;
    wire N__35749;
    wire N__35746;
    wire N__35743;
    wire N__35738;
    wire N__35735;
    wire N__35734;
    wire N__35731;
    wire N__35728;
    wire N__35725;
    wire N__35720;
    wire N__35717;
    wire N__35716;
    wire N__35713;
    wire N__35710;
    wire N__35707;
    wire N__35702;
    wire N__35699;
    wire N__35698;
    wire N__35695;
    wire N__35692;
    wire N__35689;
    wire N__35684;
    wire N__35681;
    wire N__35678;
    wire N__35675;
    wire N__35672;
    wire N__35669;
    wire N__35666;
    wire N__35663;
    wire N__35660;
    wire N__35657;
    wire N__35654;
    wire N__35651;
    wire N__35648;
    wire N__35645;
    wire N__35642;
    wire N__35639;
    wire N__35638;
    wire N__35635;
    wire N__35632;
    wire N__35629;
    wire N__35626;
    wire N__35623;
    wire N__35620;
    wire N__35615;
    wire N__35612;
    wire N__35609;
    wire N__35606;
    wire N__35603;
    wire N__35600;
    wire N__35599;
    wire N__35596;
    wire N__35593;
    wire N__35590;
    wire N__35585;
    wire N__35582;
    wire N__35579;
    wire N__35578;
    wire N__35575;
    wire N__35572;
    wire N__35569;
    wire N__35568;
    wire N__35565;
    wire N__35562;
    wire N__35559;
    wire N__35552;
    wire N__35551;
    wire N__35548;
    wire N__35545;
    wire N__35542;
    wire N__35537;
    wire N__35534;
    wire N__35531;
    wire N__35528;
    wire N__35525;
    wire N__35524;
    wire N__35521;
    wire N__35518;
    wire N__35515;
    wire N__35510;
    wire N__35507;
    wire N__35506;
    wire N__35503;
    wire N__35500;
    wire N__35497;
    wire N__35492;
    wire N__35489;
    wire N__35486;
    wire N__35483;
    wire N__35480;
    wire N__35477;
    wire N__35474;
    wire N__35471;
    wire N__35468;
    wire N__35465;
    wire N__35462;
    wire N__35459;
    wire N__35456;
    wire N__35453;
    wire N__35450;
    wire N__35447;
    wire N__35444;
    wire N__35441;
    wire N__35438;
    wire N__35435;
    wire N__35432;
    wire N__35429;
    wire N__35426;
    wire N__35423;
    wire N__35420;
    wire N__35417;
    wire N__35414;
    wire N__35411;
    wire N__35408;
    wire N__35405;
    wire N__35402;
    wire N__35399;
    wire N__35396;
    wire N__35393;
    wire N__35390;
    wire N__35387;
    wire N__35384;
    wire N__35381;
    wire N__35378;
    wire N__35375;
    wire N__35372;
    wire N__35369;
    wire N__35366;
    wire N__35363;
    wire N__35360;
    wire N__35357;
    wire N__35354;
    wire N__35351;
    wire N__35348;
    wire N__35345;
    wire N__35342;
    wire N__35339;
    wire N__35336;
    wire N__35333;
    wire N__35330;
    wire N__35327;
    wire N__35324;
    wire N__35323;
    wire N__35322;
    wire N__35321;
    wire N__35320;
    wire N__35319;
    wire N__35316;
    wire N__35315;
    wire N__35312;
    wire N__35311;
    wire N__35308;
    wire N__35303;
    wire N__35290;
    wire N__35287;
    wire N__35284;
    wire N__35279;
    wire N__35276;
    wire N__35273;
    wire N__35270;
    wire N__35267;
    wire N__35264;
    wire N__35261;
    wire N__35258;
    wire N__35255;
    wire N__35252;
    wire N__35249;
    wire N__35246;
    wire N__35243;
    wire N__35240;
    wire N__35237;
    wire N__35236;
    wire N__35233;
    wire N__35230;
    wire N__35227;
    wire N__35224;
    wire N__35219;
    wire N__35218;
    wire N__35217;
    wire N__35216;
    wire N__35213;
    wire N__35206;
    wire N__35201;
    wire N__35198;
    wire N__35195;
    wire N__35192;
    wire N__35191;
    wire N__35190;
    wire N__35189;
    wire N__35186;
    wire N__35179;
    wire N__35174;
    wire N__35173;
    wire N__35172;
    wire N__35169;
    wire N__35166;
    wire N__35163;
    wire N__35158;
    wire N__35157;
    wire N__35156;
    wire N__35153;
    wire N__35150;
    wire N__35145;
    wire N__35138;
    wire N__35135;
    wire N__35132;
    wire N__35131;
    wire N__35128;
    wire N__35125;
    wire N__35120;
    wire N__35117;
    wire N__35116;
    wire N__35113;
    wire N__35110;
    wire N__35107;
    wire N__35104;
    wire N__35101;
    wire N__35098;
    wire N__35093;
    wire N__35092;
    wire N__35089;
    wire N__35086;
    wire N__35083;
    wire N__35080;
    wire N__35077;
    wire N__35076;
    wire N__35075;
    wire N__35074;
    wire N__35071;
    wire N__35068;
    wire N__35063;
    wire N__35060;
    wire N__35057;
    wire N__35052;
    wire N__35045;
    wire N__35042;
    wire N__35041;
    wire N__35038;
    wire N__35035;
    wire N__35030;
    wire N__35027;
    wire N__35024;
    wire N__35021;
    wire N__35018;
    wire N__35015;
    wire N__35012;
    wire N__35009;
    wire N__35006;
    wire N__35003;
    wire N__35000;
    wire N__34997;
    wire N__34994;
    wire N__34991;
    wire N__34988;
    wire N__34985;
    wire N__34982;
    wire N__34979;
    wire N__34976;
    wire N__34973;
    wire N__34970;
    wire N__34967;
    wire N__34964;
    wire N__34961;
    wire N__34958;
    wire N__34955;
    wire N__34952;
    wire N__34949;
    wire N__34946;
    wire N__34943;
    wire N__34940;
    wire N__34937;
    wire N__34934;
    wire N__34931;
    wire N__34928;
    wire N__34925;
    wire N__34922;
    wire N__34919;
    wire N__34916;
    wire N__34913;
    wire N__34910;
    wire N__34907;
    wire N__34904;
    wire N__34901;
    wire N__34898;
    wire N__34895;
    wire N__34892;
    wire N__34889;
    wire N__34886;
    wire N__34883;
    wire N__34880;
    wire N__34877;
    wire N__34874;
    wire N__34871;
    wire N__34868;
    wire N__34865;
    wire N__34862;
    wire N__34859;
    wire N__34856;
    wire N__34853;
    wire N__34850;
    wire N__34847;
    wire N__34844;
    wire N__34841;
    wire N__34838;
    wire N__34835;
    wire N__34832;
    wire N__34829;
    wire N__34826;
    wire N__34823;
    wire N__34820;
    wire N__34817;
    wire N__34814;
    wire N__34811;
    wire N__34808;
    wire N__34805;
    wire N__34802;
    wire N__34799;
    wire N__34796;
    wire N__34793;
    wire N__34790;
    wire N__34787;
    wire N__34784;
    wire N__34781;
    wire N__34778;
    wire N__34775;
    wire N__34772;
    wire N__34769;
    wire N__34766;
    wire N__34763;
    wire N__34760;
    wire N__34757;
    wire N__34754;
    wire N__34751;
    wire N__34748;
    wire N__34745;
    wire N__34742;
    wire N__34739;
    wire N__34736;
    wire N__34733;
    wire N__34730;
    wire N__34727;
    wire N__34724;
    wire N__34721;
    wire N__34718;
    wire N__34715;
    wire N__34712;
    wire N__34709;
    wire N__34706;
    wire N__34703;
    wire N__34700;
    wire N__34697;
    wire N__34694;
    wire N__34691;
    wire N__34688;
    wire N__34685;
    wire N__34682;
    wire N__34679;
    wire N__34676;
    wire N__34673;
    wire N__34670;
    wire N__34667;
    wire N__34664;
    wire N__34661;
    wire N__34658;
    wire N__34655;
    wire N__34652;
    wire N__34649;
    wire N__34646;
    wire N__34643;
    wire N__34640;
    wire N__34637;
    wire N__34634;
    wire N__34631;
    wire N__34628;
    wire N__34625;
    wire N__34622;
    wire N__34619;
    wire N__34616;
    wire N__34613;
    wire N__34610;
    wire N__34607;
    wire N__34604;
    wire N__34601;
    wire N__34598;
    wire N__34595;
    wire N__34592;
    wire N__34589;
    wire N__34586;
    wire N__34583;
    wire N__34580;
    wire N__34577;
    wire N__34574;
    wire N__34571;
    wire N__34568;
    wire N__34565;
    wire N__34562;
    wire N__34559;
    wire N__34556;
    wire N__34553;
    wire N__34550;
    wire N__34547;
    wire N__34544;
    wire N__34541;
    wire N__34538;
    wire N__34535;
    wire N__34532;
    wire N__34529;
    wire N__34526;
    wire N__34523;
    wire N__34520;
    wire N__34517;
    wire N__34514;
    wire N__34511;
    wire N__34508;
    wire N__34505;
    wire N__34502;
    wire N__34499;
    wire N__34496;
    wire N__34493;
    wire N__34490;
    wire N__34487;
    wire N__34484;
    wire N__34481;
    wire N__34478;
    wire N__34475;
    wire N__34472;
    wire N__34469;
    wire N__34466;
    wire N__34463;
    wire N__34460;
    wire N__34457;
    wire N__34454;
    wire N__34451;
    wire N__34448;
    wire N__34445;
    wire N__34442;
    wire N__34439;
    wire N__34436;
    wire N__34433;
    wire N__34430;
    wire N__34427;
    wire N__34424;
    wire N__34421;
    wire N__34418;
    wire N__34415;
    wire N__34412;
    wire N__34409;
    wire N__34406;
    wire N__34403;
    wire N__34400;
    wire N__34397;
    wire N__34394;
    wire N__34391;
    wire N__34388;
    wire N__34385;
    wire N__34382;
    wire N__34379;
    wire N__34376;
    wire N__34373;
    wire N__34370;
    wire N__34367;
    wire N__34364;
    wire N__34361;
    wire N__34358;
    wire N__34355;
    wire N__34352;
    wire N__34349;
    wire N__34346;
    wire N__34343;
    wire N__34340;
    wire N__34337;
    wire N__34334;
    wire N__34333;
    wire N__34332;
    wire N__34329;
    wire N__34326;
    wire N__34323;
    wire N__34320;
    wire N__34313;
    wire N__34312;
    wire N__34309;
    wire N__34308;
    wire N__34305;
    wire N__34302;
    wire N__34299;
    wire N__34292;
    wire N__34291;
    wire N__34290;
    wire N__34287;
    wire N__34284;
    wire N__34281;
    wire N__34278;
    wire N__34271;
    wire N__34270;
    wire N__34269;
    wire N__34266;
    wire N__34263;
    wire N__34260;
    wire N__34257;
    wire N__34250;
    wire N__34247;
    wire N__34246;
    wire N__34245;
    wire N__34242;
    wire N__34239;
    wire N__34236;
    wire N__34233;
    wire N__34226;
    wire N__34225;
    wire N__34224;
    wire N__34223;
    wire N__34222;
    wire N__34221;
    wire N__34220;
    wire N__34219;
    wire N__34210;
    wire N__34209;
    wire N__34208;
    wire N__34207;
    wire N__34206;
    wire N__34205;
    wire N__34204;
    wire N__34195;
    wire N__34194;
    wire N__34193;
    wire N__34192;
    wire N__34191;
    wire N__34188;
    wire N__34183;
    wire N__34174;
    wire N__34171;
    wire N__34162;
    wire N__34161;
    wire N__34160;
    wire N__34159;
    wire N__34158;
    wire N__34157;
    wire N__34156;
    wire N__34155;
    wire N__34154;
    wire N__34143;
    wire N__34134;
    wire N__34125;
    wire N__34124;
    wire N__34123;
    wire N__34122;
    wire N__34121;
    wire N__34116;
    wire N__34113;
    wire N__34104;
    wire N__34099;
    wire N__34096;
    wire N__34093;
    wire N__34088;
    wire N__34087;
    wire N__34086;
    wire N__34083;
    wire N__34080;
    wire N__34077;
    wire N__34074;
    wire N__34067;
    wire N__34066;
    wire N__34063;
    wire N__34062;
    wire N__34059;
    wire N__34056;
    wire N__34053;
    wire N__34046;
    wire N__34045;
    wire N__34044;
    wire N__34041;
    wire N__34038;
    wire N__34035;
    wire N__34032;
    wire N__34025;
    wire N__34024;
    wire N__34023;
    wire N__34020;
    wire N__34017;
    wire N__34014;
    wire N__34011;
    wire N__34004;
    wire N__34003;
    wire N__34002;
    wire N__33999;
    wire N__33996;
    wire N__33993;
    wire N__33990;
    wire N__33983;
    wire N__33980;
    wire N__33977;
    wire N__33974;
    wire N__33973;
    wire N__33972;
    wire N__33971;
    wire N__33970;
    wire N__33969;
    wire N__33968;
    wire N__33967;
    wire N__33966;
    wire N__33965;
    wire N__33956;
    wire N__33951;
    wire N__33942;
    wire N__33935;
    wire N__33932;
    wire N__33931;
    wire N__33928;
    wire N__33925;
    wire N__33922;
    wire N__33919;
    wire N__33916;
    wire N__33913;
    wire N__33910;
    wire N__33907;
    wire N__33902;
    wire N__33899;
    wire N__33898;
    wire N__33895;
    wire N__33892;
    wire N__33889;
    wire N__33886;
    wire N__33883;
    wire N__33880;
    wire N__33877;
    wire N__33874;
    wire N__33869;
    wire N__33866;
    wire N__33863;
    wire N__33860;
    wire N__33859;
    wire N__33856;
    wire N__33853;
    wire N__33850;
    wire N__33849;
    wire N__33848;
    wire N__33845;
    wire N__33842;
    wire N__33839;
    wire N__33836;
    wire N__33833;
    wire N__33826;
    wire N__33823;
    wire N__33820;
    wire N__33815;
    wire N__33812;
    wire N__33811;
    wire N__33810;
    wire N__33807;
    wire N__33804;
    wire N__33801;
    wire N__33798;
    wire N__33795;
    wire N__33788;
    wire N__33785;
    wire N__33782;
    wire N__33779;
    wire N__33776;
    wire N__33773;
    wire N__33772;
    wire N__33771;
    wire N__33768;
    wire N__33765;
    wire N__33762;
    wire N__33759;
    wire N__33754;
    wire N__33751;
    wire N__33748;
    wire N__33743;
    wire N__33742;
    wire N__33741;
    wire N__33740;
    wire N__33739;
    wire N__33738;
    wire N__33737;
    wire N__33736;
    wire N__33719;
    wire N__33716;
    wire N__33713;
    wire N__33712;
    wire N__33709;
    wire N__33708;
    wire N__33705;
    wire N__33702;
    wire N__33699;
    wire N__33696;
    wire N__33695;
    wire N__33688;
    wire N__33685;
    wire N__33682;
    wire N__33677;
    wire N__33674;
    wire N__33671;
    wire N__33668;
    wire N__33667;
    wire N__33664;
    wire N__33661;
    wire N__33658;
    wire N__33655;
    wire N__33650;
    wire N__33649;
    wire N__33648;
    wire N__33645;
    wire N__33642;
    wire N__33639;
    wire N__33632;
    wire N__33629;
    wire N__33626;
    wire N__33623;
    wire N__33620;
    wire N__33617;
    wire N__33616;
    wire N__33615;
    wire N__33612;
    wire N__33611;
    wire N__33610;
    wire N__33609;
    wire N__33608;
    wire N__33607;
    wire N__33606;
    wire N__33605;
    wire N__33604;
    wire N__33603;
    wire N__33602;
    wire N__33601;
    wire N__33600;
    wire N__33597;
    wire N__33596;
    wire N__33595;
    wire N__33594;
    wire N__33593;
    wire N__33592;
    wire N__33591;
    wire N__33590;
    wire N__33589;
    wire N__33582;
    wire N__33573;
    wire N__33572;
    wire N__33571;
    wire N__33570;
    wire N__33569;
    wire N__33568;
    wire N__33567;
    wire N__33562;
    wire N__33561;
    wire N__33560;
    wire N__33559;
    wire N__33558;
    wire N__33557;
    wire N__33556;
    wire N__33555;
    wire N__33554;
    wire N__33553;
    wire N__33552;
    wire N__33551;
    wire N__33550;
    wire N__33549;
    wire N__33548;
    wire N__33547;
    wire N__33542;
    wire N__33529;
    wire N__33518;
    wire N__33517;
    wire N__33516;
    wire N__33515;
    wire N__33512;
    wire N__33509;
    wire N__33506;
    wire N__33493;
    wire N__33492;
    wire N__33489;
    wire N__33486;
    wire N__33471;
    wire N__33470;
    wire N__33469;
    wire N__33468;
    wire N__33467;
    wire N__33466;
    wire N__33455;
    wire N__33454;
    wire N__33453;
    wire N__33452;
    wire N__33451;
    wire N__33450;
    wire N__33447;
    wire N__33444;
    wire N__33441;
    wire N__33436;
    wire N__33435;
    wire N__33434;
    wire N__33433;
    wire N__33426;
    wire N__33417;
    wire N__33414;
    wire N__33407;
    wire N__33406;
    wire N__33405;
    wire N__33404;
    wire N__33403;
    wire N__33402;
    wire N__33401;
    wire N__33400;
    wire N__33389;
    wire N__33386;
    wire N__33385;
    wire N__33384;
    wire N__33383;
    wire N__33372;
    wire N__33367;
    wire N__33364;
    wire N__33361;
    wire N__33354;
    wire N__33349;
    wire N__33344;
    wire N__33329;
    wire N__33324;
    wire N__33317;
    wire N__33310;
    wire N__33293;
    wire N__33292;
    wire N__33291;
    wire N__33290;
    wire N__33289;
    wire N__33288;
    wire N__33287;
    wire N__33286;
    wire N__33285;
    wire N__33282;
    wire N__33281;
    wire N__33280;
    wire N__33279;
    wire N__33278;
    wire N__33277;
    wire N__33276;
    wire N__33275;
    wire N__33274;
    wire N__33273;
    wire N__33272;
    wire N__33271;
    wire N__33270;
    wire N__33269;
    wire N__33268;
    wire N__33267;
    wire N__33266;
    wire N__33265;
    wire N__33264;
    wire N__33263;
    wire N__33262;
    wire N__33261;
    wire N__33260;
    wire N__33259;
    wire N__33258;
    wire N__33255;
    wire N__33242;
    wire N__33235;
    wire N__33234;
    wire N__33231;
    wire N__33230;
    wire N__33229;
    wire N__33228;
    wire N__33225;
    wire N__33224;
    wire N__33223;
    wire N__33222;
    wire N__33221;
    wire N__33220;
    wire N__33219;
    wire N__33218;
    wire N__33215;
    wire N__33212;
    wire N__33211;
    wire N__33210;
    wire N__33209;
    wire N__33208;
    wire N__33205;
    wire N__33202;
    wire N__33199;
    wire N__33194;
    wire N__33193;
    wire N__33192;
    wire N__33191;
    wire N__33188;
    wire N__33187;
    wire N__33186;
    wire N__33185;
    wire N__33184;
    wire N__33181;
    wire N__33180;
    wire N__33179;
    wire N__33176;
    wire N__33173;
    wire N__33170;
    wire N__33169;
    wire N__33168;
    wire N__33167;
    wire N__33166;
    wire N__33165;
    wire N__33162;
    wire N__33161;
    wire N__33160;
    wire N__33157;
    wire N__33156;
    wire N__33153;
    wire N__33152;
    wire N__33149;
    wire N__33148;
    wire N__33147;
    wire N__33144;
    wire N__33143;
    wire N__33140;
    wire N__33139;
    wire N__33136;
    wire N__33135;
    wire N__33132;
    wire N__33131;
    wire N__33130;
    wire N__33129;
    wire N__33128;
    wire N__33127;
    wire N__33126;
    wire N__33125;
    wire N__33124;
    wire N__33123;
    wire N__33122;
    wire N__33121;
    wire N__33120;
    wire N__33119;
    wire N__33118;
    wire N__33115;
    wire N__33114;
    wire N__33111;
    wire N__33106;
    wire N__33103;
    wire N__33092;
    wire N__33087;
    wire N__33086;
    wire N__33083;
    wire N__33080;
    wire N__33079;
    wire N__33076;
    wire N__33075;
    wire N__33072;
    wire N__33069;
    wire N__33068;
    wire N__33067;
    wire N__33066;
    wire N__33065;
    wire N__33060;
    wire N__33045;
    wire N__33042;
    wire N__33041;
    wire N__33038;
    wire N__33037;
    wire N__33034;
    wire N__33033;
    wire N__33030;
    wire N__33029;
    wire N__33024;
    wire N__33011;
    wire N__33004;
    wire N__32991;
    wire N__32974;
    wire N__32957;
    wire N__32954;
    wire N__32953;
    wire N__32950;
    wire N__32949;
    wire N__32946;
    wire N__32945;
    wire N__32942;
    wire N__32941;
    wire N__32940;
    wire N__32937;
    wire N__32936;
    wire N__32933;
    wire N__32932;
    wire N__32929;
    wire N__32928;
    wire N__32925;
    wire N__32924;
    wire N__32921;
    wire N__32920;
    wire N__32917;
    wire N__32916;
    wire N__32913;
    wire N__32912;
    wire N__32911;
    wire N__32910;
    wire N__32899;
    wire N__32892;
    wire N__32889;
    wire N__32886;
    wire N__32883;
    wire N__32878;
    wire N__32867;
    wire N__32864;
    wire N__32863;
    wire N__32860;
    wire N__32859;
    wire N__32856;
    wire N__32855;
    wire N__32852;
    wire N__32851;
    wire N__32848;
    wire N__32843;
    wire N__32828;
    wire N__32815;
    wire N__32798;
    wire N__32781;
    wire N__32768;
    wire N__32765;
    wire N__32764;
    wire N__32761;
    wire N__32760;
    wire N__32757;
    wire N__32756;
    wire N__32753;
    wire N__32750;
    wire N__32747;
    wire N__32738;
    wire N__32721;
    wire N__32706;
    wire N__32693;
    wire N__32678;
    wire N__32675;
    wire N__32674;
    wire N__32671;
    wire N__32668;
    wire N__32667;
    wire N__32662;
    wire N__32659;
    wire N__32656;
    wire N__32653;
    wire N__32652;
    wire N__32649;
    wire N__32646;
    wire N__32643;
    wire N__32636;
    wire N__32633;
    wire N__32632;
    wire N__32629;
    wire N__32626;
    wire N__32625;
    wire N__32620;
    wire N__32617;
    wire N__32612;
    wire N__32609;
    wire N__32606;
    wire N__32603;
    wire N__32600;
    wire N__32597;
    wire N__32594;
    wire N__32591;
    wire N__32588;
    wire N__32585;
    wire N__32584;
    wire N__32583;
    wire N__32582;
    wire N__32579;
    wire N__32576;
    wire N__32573;
    wire N__32570;
    wire N__32565;
    wire N__32562;
    wire N__32559;
    wire N__32556;
    wire N__32551;
    wire N__32548;
    wire N__32545;
    wire N__32540;
    wire N__32537;
    wire N__32534;
    wire N__32531;
    wire N__32528;
    wire N__32525;
    wire N__32522;
    wire N__32519;
    wire N__32516;
    wire N__32515;
    wire N__32512;
    wire N__32509;
    wire N__32506;
    wire N__32503;
    wire N__32500;
    wire N__32499;
    wire N__32496;
    wire N__32493;
    wire N__32490;
    wire N__32483;
    wire N__32482;
    wire N__32479;
    wire N__32476;
    wire N__32473;
    wire N__32470;
    wire N__32467;
    wire N__32464;
    wire N__32461;
    wire N__32460;
    wire N__32459;
    wire N__32456;
    wire N__32453;
    wire N__32450;
    wire N__32447;
    wire N__32444;
    wire N__32437;
    wire N__32432;
    wire N__32429;
    wire N__32426;
    wire N__32423;
    wire N__32422;
    wire N__32419;
    wire N__32418;
    wire N__32415;
    wire N__32412;
    wire N__32409;
    wire N__32406;
    wire N__32401;
    wire N__32400;
    wire N__32397;
    wire N__32394;
    wire N__32391;
    wire N__32384;
    wire N__32381;
    wire N__32378;
    wire N__32375;
    wire N__32374;
    wire N__32371;
    wire N__32368;
    wire N__32363;
    wire N__32362;
    wire N__32359;
    wire N__32356;
    wire N__32351;
    wire N__32348;
    wire N__32345;
    wire N__32342;
    wire N__32339;
    wire N__32338;
    wire N__32335;
    wire N__32332;
    wire N__32329;
    wire N__32328;
    wire N__32325;
    wire N__32322;
    wire N__32319;
    wire N__32318;
    wire N__32315;
    wire N__32310;
    wire N__32307;
    wire N__32302;
    wire N__32299;
    wire N__32294;
    wire N__32291;
    wire N__32290;
    wire N__32287;
    wire N__32284;
    wire N__32283;
    wire N__32280;
    wire N__32277;
    wire N__32274;
    wire N__32267;
    wire N__32264;
    wire N__32261;
    wire N__32258;
    wire N__32255;
    wire N__32252;
    wire N__32249;
    wire N__32248;
    wire N__32245;
    wire N__32242;
    wire N__32239;
    wire N__32238;
    wire N__32235;
    wire N__32234;
    wire N__32231;
    wire N__32228;
    wire N__32225;
    wire N__32222;
    wire N__32219;
    wire N__32216;
    wire N__32211;
    wire N__32208;
    wire N__32205;
    wire N__32202;
    wire N__32195;
    wire N__32194;
    wire N__32191;
    wire N__32188;
    wire N__32187;
    wire N__32184;
    wire N__32181;
    wire N__32178;
    wire N__32175;
    wire N__32170;
    wire N__32165;
    wire N__32162;
    wire N__32159;
    wire N__32156;
    wire N__32155;
    wire N__32152;
    wire N__32149;
    wire N__32144;
    wire N__32143;
    wire N__32140;
    wire N__32139;
    wire N__32136;
    wire N__32133;
    wire N__32130;
    wire N__32127;
    wire N__32122;
    wire N__32117;
    wire N__32114;
    wire N__32113;
    wire N__32112;
    wire N__32109;
    wire N__32106;
    wire N__32103;
    wire N__32098;
    wire N__32095;
    wire N__32092;
    wire N__32089;
    wire N__32084;
    wire N__32081;
    wire N__32078;
    wire N__32075;
    wire N__32072;
    wire N__32069;
    wire N__32066;
    wire N__32063;
    wire N__32060;
    wire N__32057;
    wire N__32054;
    wire N__32053;
    wire N__32050;
    wire N__32047;
    wire N__32042;
    wire N__32041;
    wire N__32036;
    wire N__32033;
    wire N__32030;
    wire N__32027;
    wire N__32024;
    wire N__32023;
    wire N__32022;
    wire N__32015;
    wire N__32012;
    wire N__32009;
    wire N__32006;
    wire N__32003;
    wire N__32000;
    wire N__31999;
    wire N__31996;
    wire N__31993;
    wire N__31988;
    wire N__31985;
    wire N__31984;
    wire N__31983;
    wire N__31982;
    wire N__31979;
    wire N__31974;
    wire N__31971;
    wire N__31968;
    wire N__31965;
    wire N__31962;
    wire N__31959;
    wire N__31958;
    wire N__31955;
    wire N__31952;
    wire N__31949;
    wire N__31946;
    wire N__31943;
    wire N__31934;
    wire N__31933;
    wire N__31928;
    wire N__31925;
    wire N__31922;
    wire N__31921;
    wire N__31918;
    wire N__31915;
    wire N__31910;
    wire N__31907;
    wire N__31906;
    wire N__31903;
    wire N__31900;
    wire N__31895;
    wire N__31892;
    wire N__31891;
    wire N__31890;
    wire N__31885;
    wire N__31882;
    wire N__31879;
    wire N__31878;
    wire N__31873;
    wire N__31870;
    wire N__31865;
    wire N__31862;
    wire N__31859;
    wire N__31856;
    wire N__31853;
    wire N__31852;
    wire N__31849;
    wire N__31846;
    wire N__31841;
    wire N__31838;
    wire N__31837;
    wire N__31834;
    wire N__31831;
    wire N__31830;
    wire N__31825;
    wire N__31822;
    wire N__31819;
    wire N__31816;
    wire N__31813;
    wire N__31808;
    wire N__31805;
    wire N__31802;
    wire N__31801;
    wire N__31800;
    wire N__31799;
    wire N__31796;
    wire N__31793;
    wire N__31790;
    wire N__31787;
    wire N__31784;
    wire N__31781;
    wire N__31772;
    wire N__31769;
    wire N__31768;
    wire N__31765;
    wire N__31762;
    wire N__31761;
    wire N__31758;
    wire N__31755;
    wire N__31752;
    wire N__31749;
    wire N__31746;
    wire N__31743;
    wire N__31738;
    wire N__31733;
    wire N__31732;
    wire N__31731;
    wire N__31728;
    wire N__31725;
    wire N__31722;
    wire N__31719;
    wire N__31716;
    wire N__31715;
    wire N__31712;
    wire N__31709;
    wire N__31706;
    wire N__31703;
    wire N__31698;
    wire N__31695;
    wire N__31690;
    wire N__31685;
    wire N__31682;
    wire N__31679;
    wire N__31676;
    wire N__31673;
    wire N__31672;
    wire N__31667;
    wire N__31664;
    wire N__31661;
    wire N__31660;
    wire N__31659;
    wire N__31656;
    wire N__31653;
    wire N__31648;
    wire N__31643;
    wire N__31642;
    wire N__31641;
    wire N__31638;
    wire N__31635;
    wire N__31630;
    wire N__31625;
    wire N__31622;
    wire N__31619;
    wire N__31616;
    wire N__31613;
    wire N__31612;
    wire N__31609;
    wire N__31608;
    wire N__31605;
    wire N__31602;
    wire N__31599;
    wire N__31592;
    wire N__31589;
    wire N__31586;
    wire N__31585;
    wire N__31584;
    wire N__31581;
    wire N__31578;
    wire N__31575;
    wire N__31574;
    wire N__31571;
    wire N__31568;
    wire N__31565;
    wire N__31562;
    wire N__31555;
    wire N__31550;
    wire N__31549;
    wire N__31544;
    wire N__31541;
    wire N__31538;
    wire N__31535;
    wire N__31534;
    wire N__31533;
    wire N__31530;
    wire N__31527;
    wire N__31524;
    wire N__31521;
    wire N__31518;
    wire N__31511;
    wire N__31510;
    wire N__31507;
    wire N__31504;
    wire N__31503;
    wire N__31502;
    wire N__31499;
    wire N__31496;
    wire N__31493;
    wire N__31490;
    wire N__31487;
    wire N__31482;
    wire N__31479;
    wire N__31476;
    wire N__31471;
    wire N__31466;
    wire N__31465;
    wire N__31460;
    wire N__31457;
    wire N__31454;
    wire N__31451;
    wire N__31448;
    wire N__31445;
    wire N__31444;
    wire N__31443;
    wire N__31440;
    wire N__31435;
    wire N__31430;
    wire N__31427;
    wire N__31426;
    wire N__31425;
    wire N__31420;
    wire N__31417;
    wire N__31414;
    wire N__31409;
    wire N__31406;
    wire N__31403;
    wire N__31400;
    wire N__31397;
    wire N__31394;
    wire N__31391;
    wire N__31390;
    wire N__31385;
    wire N__31382;
    wire N__31379;
    wire N__31378;
    wire N__31375;
    wire N__31374;
    wire N__31371;
    wire N__31368;
    wire N__31365;
    wire N__31358;
    wire N__31357;
    wire N__31356;
    wire N__31353;
    wire N__31350;
    wire N__31347;
    wire N__31346;
    wire N__31343;
    wire N__31338;
    wire N__31335;
    wire N__31332;
    wire N__31329;
    wire N__31326;
    wire N__31319;
    wire N__31316;
    wire N__31313;
    wire N__31312;
    wire N__31307;
    wire N__31304;
    wire N__31303;
    wire N__31302;
    wire N__31299;
    wire N__31296;
    wire N__31293;
    wire N__31286;
    wire N__31285;
    wire N__31282;
    wire N__31279;
    wire N__31276;
    wire N__31273;
    wire N__31270;
    wire N__31265;
    wire N__31264;
    wire N__31263;
    wire N__31260;
    wire N__31257;
    wire N__31254;
    wire N__31247;
    wire N__31244;
    wire N__31241;
    wire N__31238;
    wire N__31235;
    wire N__31234;
    wire N__31231;
    wire N__31228;
    wire N__31223;
    wire N__31222;
    wire N__31219;
    wire N__31218;
    wire N__31215;
    wire N__31212;
    wire N__31209;
    wire N__31206;
    wire N__31203;
    wire N__31196;
    wire N__31195;
    wire N__31192;
    wire N__31189;
    wire N__31186;
    wire N__31183;
    wire N__31180;
    wire N__31177;
    wire N__31174;
    wire N__31169;
    wire N__31168;
    wire N__31165;
    wire N__31164;
    wire N__31161;
    wire N__31158;
    wire N__31155;
    wire N__31152;
    wire N__31149;
    wire N__31142;
    wire N__31139;
    wire N__31136;
    wire N__31133;
    wire N__31130;
    wire N__31127;
    wire N__31126;
    wire N__31125;
    wire N__31118;
    wire N__31115;
    wire N__31112;
    wire N__31111;
    wire N__31108;
    wire N__31105;
    wire N__31100;
    wire N__31097;
    wire N__31094;
    wire N__31091;
    wire N__31088;
    wire N__31085;
    wire N__31082;
    wire N__31079;
    wire N__31076;
    wire N__31073;
    wire N__31070;
    wire N__31069;
    wire N__31068;
    wire N__31067;
    wire N__31064;
    wire N__31057;
    wire N__31052;
    wire N__31051;
    wire N__31050;
    wire N__31043;
    wire N__31040;
    wire N__31037;
    wire N__31034;
    wire N__31031;
    wire N__31028;
    wire N__31025;
    wire N__31022;
    wire N__31019;
    wire N__31016;
    wire N__31013;
    wire N__31010;
    wire N__31007;
    wire N__31004;
    wire N__31001;
    wire N__30998;
    wire N__30995;
    wire N__30992;
    wire N__30989;
    wire N__30986;
    wire N__30983;
    wire N__30980;
    wire N__30977;
    wire N__30974;
    wire N__30971;
    wire N__30970;
    wire N__30969;
    wire N__30968;
    wire N__30967;
    wire N__30966;
    wire N__30965;
    wire N__30964;
    wire N__30963;
    wire N__30962;
    wire N__30961;
    wire N__30960;
    wire N__30959;
    wire N__30958;
    wire N__30957;
    wire N__30956;
    wire N__30955;
    wire N__30954;
    wire N__30953;
    wire N__30952;
    wire N__30947;
    wire N__30940;
    wire N__30939;
    wire N__30922;
    wire N__30907;
    wire N__30904;
    wire N__30901;
    wire N__30900;
    wire N__30899;
    wire N__30898;
    wire N__30897;
    wire N__30896;
    wire N__30895;
    wire N__30892;
    wire N__30891;
    wire N__30886;
    wire N__30881;
    wire N__30878;
    wire N__30877;
    wire N__30874;
    wire N__30871;
    wire N__30870;
    wire N__30869;
    wire N__30866;
    wire N__30863;
    wire N__30860;
    wire N__30859;
    wire N__30854;
    wire N__30851;
    wire N__30848;
    wire N__30845;
    wire N__30832;
    wire N__30825;
    wire N__30820;
    wire N__30817;
    wire N__30806;
    wire N__30803;
    wire N__30800;
    wire N__30797;
    wire N__30794;
    wire N__30791;
    wire N__30788;
    wire N__30785;
    wire N__30782;
    wire N__30779;
    wire N__30776;
    wire N__30773;
    wire N__30770;
    wire N__30769;
    wire N__30768;
    wire N__30767;
    wire N__30764;
    wire N__30761;
    wire N__30758;
    wire N__30755;
    wire N__30752;
    wire N__30749;
    wire N__30746;
    wire N__30741;
    wire N__30738;
    wire N__30735;
    wire N__30730;
    wire N__30725;
    wire N__30722;
    wire N__30719;
    wire N__30718;
    wire N__30715;
    wire N__30714;
    wire N__30711;
    wire N__30708;
    wire N__30705;
    wire N__30698;
    wire N__30695;
    wire N__30692;
    wire N__30689;
    wire N__30686;
    wire N__30683;
    wire N__30680;
    wire N__30679;
    wire N__30676;
    wire N__30673;
    wire N__30668;
    wire N__30665;
    wire N__30662;
    wire N__30659;
    wire N__30656;
    wire N__30653;
    wire N__30650;
    wire N__30647;
    wire N__30644;
    wire N__30641;
    wire N__30638;
    wire N__30635;
    wire N__30632;
    wire N__30629;
    wire N__30626;
    wire N__30623;
    wire N__30620;
    wire N__30617;
    wire N__30614;
    wire N__30611;
    wire N__30608;
    wire N__30605;
    wire N__30602;
    wire N__30599;
    wire N__30596;
    wire N__30593;
    wire N__30590;
    wire N__30587;
    wire N__30584;
    wire N__30581;
    wire N__30580;
    wire N__30577;
    wire N__30574;
    wire N__30573;
    wire N__30570;
    wire N__30567;
    wire N__30564;
    wire N__30561;
    wire N__30556;
    wire N__30555;
    wire N__30552;
    wire N__30549;
    wire N__30546;
    wire N__30539;
    wire N__30538;
    wire N__30535;
    wire N__30532;
    wire N__30529;
    wire N__30526;
    wire N__30525;
    wire N__30522;
    wire N__30519;
    wire N__30516;
    wire N__30509;
    wire N__30506;
    wire N__30503;
    wire N__30500;
    wire N__30499;
    wire N__30496;
    wire N__30495;
    wire N__30492;
    wire N__30491;
    wire N__30488;
    wire N__30485;
    wire N__30482;
    wire N__30479;
    wire N__30476;
    wire N__30473;
    wire N__30468;
    wire N__30465;
    wire N__30462;
    wire N__30459;
    wire N__30452;
    wire N__30451;
    wire N__30450;
    wire N__30447;
    wire N__30444;
    wire N__30441;
    wire N__30438;
    wire N__30435;
    wire N__30432;
    wire N__30425;
    wire N__30422;
    wire N__30419;
    wire N__30416;
    wire N__30413;
    wire N__30412;
    wire N__30409;
    wire N__30406;
    wire N__30405;
    wire N__30400;
    wire N__30397;
    wire N__30396;
    wire N__30393;
    wire N__30390;
    wire N__30387;
    wire N__30384;
    wire N__30379;
    wire N__30374;
    wire N__30371;
    wire N__30370;
    wire N__30369;
    wire N__30366;
    wire N__30363;
    wire N__30360;
    wire N__30353;
    wire N__30350;
    wire N__30347;
    wire N__30344;
    wire N__30341;
    wire N__30338;
    wire N__30337;
    wire N__30334;
    wire N__30331;
    wire N__30328;
    wire N__30327;
    wire N__30324;
    wire N__30321;
    wire N__30318;
    wire N__30311;
    wire N__30310;
    wire N__30307;
    wire N__30304;
    wire N__30303;
    wire N__30300;
    wire N__30297;
    wire N__30294;
    wire N__30287;
    wire N__30286;
    wire N__30283;
    wire N__30280;
    wire N__30275;
    wire N__30272;
    wire N__30269;
    wire N__30266;
    wire N__30263;
    wire N__30260;
    wire N__30259;
    wire N__30256;
    wire N__30253;
    wire N__30250;
    wire N__30249;
    wire N__30246;
    wire N__30243;
    wire N__30240;
    wire N__30237;
    wire N__30236;
    wire N__30231;
    wire N__30228;
    wire N__30225;
    wire N__30222;
    wire N__30217;
    wire N__30212;
    wire N__30209;
    wire N__30206;
    wire N__30203;
    wire N__30202;
    wire N__30199;
    wire N__30196;
    wire N__30195;
    wire N__30190;
    wire N__30187;
    wire N__30182;
    wire N__30179;
    wire N__30176;
    wire N__30173;
    wire N__30170;
    wire N__30169;
    wire N__30168;
    wire N__30165;
    wire N__30160;
    wire N__30159;
    wire N__30156;
    wire N__30153;
    wire N__30150;
    wire N__30147;
    wire N__30142;
    wire N__30139;
    wire N__30136;
    wire N__30131;
    wire N__30130;
    wire N__30127;
    wire N__30126;
    wire N__30123;
    wire N__30120;
    wire N__30117;
    wire N__30110;
    wire N__30107;
    wire N__30104;
    wire N__30101;
    wire N__30098;
    wire N__30095;
    wire N__30094;
    wire N__30091;
    wire N__30090;
    wire N__30087;
    wire N__30084;
    wire N__30081;
    wire N__30074;
    wire N__30073;
    wire N__30070;
    wire N__30069;
    wire N__30066;
    wire N__30063;
    wire N__30060;
    wire N__30057;
    wire N__30056;
    wire N__30053;
    wire N__30050;
    wire N__30047;
    wire N__30044;
    wire N__30041;
    wire N__30038;
    wire N__30033;
    wire N__30026;
    wire N__30023;
    wire N__30020;
    wire N__30017;
    wire N__30014;
    wire N__30011;
    wire N__30008;
    wire N__30007;
    wire N__30006;
    wire N__30005;
    wire N__30002;
    wire N__29999;
    wire N__29996;
    wire N__29993;
    wire N__29990;
    wire N__29987;
    wire N__29982;
    wire N__29977;
    wire N__29974;
    wire N__29969;
    wire N__29966;
    wire N__29965;
    wire N__29964;
    wire N__29961;
    wire N__29958;
    wire N__29955;
    wire N__29948;
    wire N__29945;
    wire N__29942;
    wire N__29939;
    wire N__29936;
    wire N__29933;
    wire N__29930;
    wire N__29929;
    wire N__29928;
    wire N__29927;
    wire N__29918;
    wire N__29915;
    wire N__29914;
    wire N__29911;
    wire N__29910;
    wire N__29903;
    wire N__29900;
    wire N__29897;
    wire N__29894;
    wire N__29891;
    wire N__29888;
    wire N__29887;
    wire N__29886;
    wire N__29883;
    wire N__29882;
    wire N__29879;
    wire N__29876;
    wire N__29875;
    wire N__29872;
    wire N__29869;
    wire N__29866;
    wire N__29863;
    wire N__29860;
    wire N__29857;
    wire N__29854;
    wire N__29847;
    wire N__29844;
    wire N__29841;
    wire N__29838;
    wire N__29835;
    wire N__29830;
    wire N__29825;
    wire N__29822;
    wire N__29819;
    wire N__29816;
    wire N__29815;
    wire N__29812;
    wire N__29809;
    wire N__29806;
    wire N__29803;
    wire N__29802;
    wire N__29799;
    wire N__29796;
    wire N__29793;
    wire N__29788;
    wire N__29785;
    wire N__29784;
    wire N__29781;
    wire N__29778;
    wire N__29775;
    wire N__29768;
    wire N__29767;
    wire N__29764;
    wire N__29761;
    wire N__29760;
    wire N__29757;
    wire N__29754;
    wire N__29751;
    wire N__29744;
    wire N__29741;
    wire N__29738;
    wire N__29735;
    wire N__29732;
    wire N__29729;
    wire N__29726;
    wire N__29723;
    wire N__29720;
    wire N__29719;
    wire N__29716;
    wire N__29713;
    wire N__29710;
    wire N__29709;
    wire N__29706;
    wire N__29703;
    wire N__29700;
    wire N__29693;
    wire N__29692;
    wire N__29691;
    wire N__29688;
    wire N__29685;
    wire N__29682;
    wire N__29679;
    wire N__29676;
    wire N__29675;
    wire N__29672;
    wire N__29669;
    wire N__29666;
    wire N__29663;
    wire N__29660;
    wire N__29653;
    wire N__29648;
    wire N__29645;
    wire N__29642;
    wire N__29639;
    wire N__29636;
    wire N__29635;
    wire N__29632;
    wire N__29629;
    wire N__29628;
    wire N__29625;
    wire N__29622;
    wire N__29619;
    wire N__29616;
    wire N__29613;
    wire N__29610;
    wire N__29607;
    wire N__29604;
    wire N__29601;
    wire N__29600;
    wire N__29595;
    wire N__29592;
    wire N__29589;
    wire N__29582;
    wire N__29579;
    wire N__29576;
    wire N__29575;
    wire N__29574;
    wire N__29571;
    wire N__29568;
    wire N__29565;
    wire N__29560;
    wire N__29557;
    wire N__29552;
    wire N__29549;
    wire N__29546;
    wire N__29543;
    wire N__29540;
    wire N__29537;
    wire N__29534;
    wire N__29533;
    wire N__29532;
    wire N__29529;
    wire N__29526;
    wire N__29523;
    wire N__29520;
    wire N__29519;
    wire N__29516;
    wire N__29513;
    wire N__29510;
    wire N__29507;
    wire N__29504;
    wire N__29501;
    wire N__29496;
    wire N__29489;
    wire N__29488;
    wire N__29485;
    wire N__29482;
    wire N__29479;
    wire N__29478;
    wire N__29475;
    wire N__29472;
    wire N__29469;
    wire N__29462;
    wire N__29459;
    wire N__29456;
    wire N__29453;
    wire N__29450;
    wire N__29447;
    wire N__29446;
    wire N__29443;
    wire N__29440;
    wire N__29437;
    wire N__29434;
    wire N__29431;
    wire N__29428;
    wire N__29425;
    wire N__29420;
    wire N__29417;
    wire N__29414;
    wire N__29411;
    wire N__29408;
    wire N__29405;
    wire N__29402;
    wire N__29399;
    wire N__29396;
    wire N__29393;
    wire N__29390;
    wire N__29387;
    wire N__29384;
    wire N__29381;
    wire N__29378;
    wire N__29375;
    wire N__29372;
    wire N__29369;
    wire N__29366;
    wire N__29363;
    wire N__29360;
    wire N__29357;
    wire N__29354;
    wire N__29351;
    wire N__29348;
    wire N__29345;
    wire N__29342;
    wire N__29339;
    wire N__29336;
    wire N__29333;
    wire N__29330;
    wire N__29327;
    wire N__29324;
    wire N__29321;
    wire N__29318;
    wire N__29315;
    wire N__29314;
    wire N__29313;
    wire N__29312;
    wire N__29311;
    wire N__29310;
    wire N__29309;
    wire N__29308;
    wire N__29307;
    wire N__29306;
    wire N__29305;
    wire N__29304;
    wire N__29303;
    wire N__29302;
    wire N__29301;
    wire N__29298;
    wire N__29291;
    wire N__29278;
    wire N__29271;
    wire N__29266;
    wire N__29263;
    wire N__29260;
    wire N__29257;
    wire N__29252;
    wire N__29249;
    wire N__29246;
    wire N__29243;
    wire N__29240;
    wire N__29231;
    wire N__29228;
    wire N__29225;
    wire N__29222;
    wire N__29219;
    wire N__29218;
    wire N__29217;
    wire N__29214;
    wire N__29211;
    wire N__29210;
    wire N__29207;
    wire N__29204;
    wire N__29201;
    wire N__29198;
    wire N__29195;
    wire N__29192;
    wire N__29189;
    wire N__29186;
    wire N__29183;
    wire N__29180;
    wire N__29177;
    wire N__29174;
    wire N__29171;
    wire N__29164;
    wire N__29159;
    wire N__29158;
    wire N__29153;
    wire N__29150;
    wire N__29147;
    wire N__29144;
    wire N__29143;
    wire N__29142;
    wire N__29139;
    wire N__29136;
    wire N__29133;
    wire N__29130;
    wire N__29123;
    wire N__29122;
    wire N__29121;
    wire N__29120;
    wire N__29119;
    wire N__29118;
    wire N__29117;
    wire N__29116;
    wire N__29115;
    wire N__29114;
    wire N__29113;
    wire N__29112;
    wire N__29111;
    wire N__29110;
    wire N__29109;
    wire N__29108;
    wire N__29107;
    wire N__29106;
    wire N__29105;
    wire N__29104;
    wire N__29103;
    wire N__29102;
    wire N__29101;
    wire N__29100;
    wire N__29091;
    wire N__29082;
    wire N__29073;
    wire N__29064;
    wire N__29063;
    wire N__29062;
    wire N__29061;
    wire N__29060;
    wire N__29059;
    wire N__29058;
    wire N__29049;
    wire N__29040;
    wire N__29031;
    wire N__29026;
    wire N__29017;
    wire N__29010;
    wire N__29005;
    wire N__29002;
    wire N__28999;
    wire N__28996;
    wire N__28991;
    wire N__28988;
    wire N__28985;
    wire N__28982;
    wire N__28979;
    wire N__28976;
    wire N__28973;
    wire N__28970;
    wire N__28967;
    wire N__28964;
    wire N__28961;
    wire N__28958;
    wire N__28955;
    wire N__28952;
    wire N__28949;
    wire N__28946;
    wire N__28943;
    wire N__28940;
    wire N__28937;
    wire N__28934;
    wire N__28931;
    wire N__28928;
    wire N__28925;
    wire N__28922;
    wire N__28919;
    wire N__28916;
    wire N__28913;
    wire N__28910;
    wire N__28907;
    wire N__28904;
    wire N__28901;
    wire N__28898;
    wire N__28895;
    wire N__28892;
    wire N__28889;
    wire N__28886;
    wire N__28883;
    wire N__28880;
    wire N__28877;
    wire N__28874;
    wire N__28871;
    wire N__28868;
    wire N__28865;
    wire N__28862;
    wire N__28859;
    wire N__28856;
    wire N__28853;
    wire N__28850;
    wire N__28847;
    wire N__28844;
    wire N__28841;
    wire N__28838;
    wire N__28835;
    wire N__28832;
    wire N__28829;
    wire N__28826;
    wire N__28823;
    wire N__28820;
    wire N__28817;
    wire N__28814;
    wire N__28811;
    wire N__28808;
    wire N__28805;
    wire N__28802;
    wire N__28799;
    wire N__28796;
    wire N__28793;
    wire N__28790;
    wire N__28787;
    wire N__28784;
    wire N__28781;
    wire N__28778;
    wire N__28775;
    wire N__28772;
    wire N__28769;
    wire N__28766;
    wire N__28763;
    wire N__28760;
    wire N__28757;
    wire N__28754;
    wire N__28751;
    wire N__28748;
    wire N__28745;
    wire N__28744;
    wire N__28743;
    wire N__28740;
    wire N__28739;
    wire N__28736;
    wire N__28733;
    wire N__28730;
    wire N__28727;
    wire N__28724;
    wire N__28721;
    wire N__28718;
    wire N__28715;
    wire N__28706;
    wire N__28705;
    wire N__28702;
    wire N__28701;
    wire N__28698;
    wire N__28695;
    wire N__28692;
    wire N__28689;
    wire N__28686;
    wire N__28679;
    wire N__28676;
    wire N__28673;
    wire N__28670;
    wire N__28667;
    wire N__28666;
    wire N__28663;
    wire N__28662;
    wire N__28659;
    wire N__28656;
    wire N__28653;
    wire N__28646;
    wire N__28645;
    wire N__28642;
    wire N__28641;
    wire N__28640;
    wire N__28637;
    wire N__28634;
    wire N__28631;
    wire N__28628;
    wire N__28625;
    wire N__28620;
    wire N__28617;
    wire N__28614;
    wire N__28609;
    wire N__28604;
    wire N__28601;
    wire N__28600;
    wire N__28595;
    wire N__28592;
    wire N__28591;
    wire N__28588;
    wire N__28585;
    wire N__28584;
    wire N__28581;
    wire N__28578;
    wire N__28577;
    wire N__28574;
    wire N__28571;
    wire N__28568;
    wire N__28565;
    wire N__28562;
    wire N__28559;
    wire N__28554;
    wire N__28551;
    wire N__28548;
    wire N__28545;
    wire N__28538;
    wire N__28535;
    wire N__28534;
    wire N__28531;
    wire N__28530;
    wire N__28527;
    wire N__28524;
    wire N__28521;
    wire N__28514;
    wire N__28513;
    wire N__28512;
    wire N__28511;
    wire N__28510;
    wire N__28509;
    wire N__28508;
    wire N__28507;
    wire N__28506;
    wire N__28505;
    wire N__28504;
    wire N__28503;
    wire N__28502;
    wire N__28475;
    wire N__28472;
    wire N__28469;
    wire N__28466;
    wire N__28463;
    wire N__28462;
    wire N__28459;
    wire N__28456;
    wire N__28451;
    wire N__28450;
    wire N__28449;
    wire N__28446;
    wire N__28443;
    wire N__28440;
    wire N__28437;
    wire N__28430;
    wire N__28427;
    wire N__28426;
    wire N__28423;
    wire N__28422;
    wire N__28419;
    wire N__28416;
    wire N__28413;
    wire N__28410;
    wire N__28407;
    wire N__28400;
    wire N__28397;
    wire N__28394;
    wire N__28393;
    wire N__28390;
    wire N__28387;
    wire N__28382;
    wire N__28379;
    wire N__28376;
    wire N__28373;
    wire N__28370;
    wire N__28367;
    wire N__28366;
    wire N__28363;
    wire N__28360;
    wire N__28357;
    wire N__28354;
    wire N__28351;
    wire N__28348;
    wire N__28343;
    wire N__28340;
    wire N__28337;
    wire N__28334;
    wire N__28331;
    wire N__28330;
    wire N__28327;
    wire N__28326;
    wire N__28321;
    wire N__28318;
    wire N__28317;
    wire N__28314;
    wire N__28311;
    wire N__28308;
    wire N__28301;
    wire N__28298;
    wire N__28297;
    wire N__28294;
    wire N__28291;
    wire N__28288;
    wire N__28283;
    wire N__28280;
    wire N__28279;
    wire N__28278;
    wire N__28277;
    wire N__28274;
    wire N__28267;
    wire N__28262;
    wire N__28261;
    wire N__28258;
    wire N__28257;
    wire N__28256;
    wire N__28247;
    wire N__28244;
    wire N__28241;
    wire N__28238;
    wire N__28237;
    wire N__28234;
    wire N__28231;
    wire N__28228;
    wire N__28225;
    wire N__28222;
    wire N__28219;
    wire N__28214;
    wire N__28211;
    wire N__28210;
    wire N__28209;
    wire N__28204;
    wire N__28201;
    wire N__28198;
    wire N__28197;
    wire N__28196;
    wire N__28193;
    wire N__28190;
    wire N__28185;
    wire N__28178;
    wire N__28175;
    wire N__28174;
    wire N__28173;
    wire N__28170;
    wire N__28167;
    wire N__28166;
    wire N__28163;
    wire N__28158;
    wire N__28155;
    wire N__28152;
    wire N__28149;
    wire N__28146;
    wire N__28143;
    wire N__28140;
    wire N__28137;
    wire N__28130;
    wire N__28127;
    wire N__28126;
    wire N__28125;
    wire N__28122;
    wire N__28119;
    wire N__28116;
    wire N__28113;
    wire N__28110;
    wire N__28103;
    wire N__28100;
    wire N__28097;
    wire N__28094;
    wire N__28091;
    wire N__28090;
    wire N__28089;
    wire N__28084;
    wire N__28081;
    wire N__28078;
    wire N__28073;
    wire N__28070;
    wire N__28069;
    wire N__28064;
    wire N__28061;
    wire N__28058;
    wire N__28055;
    wire N__28052;
    wire N__28051;
    wire N__28048;
    wire N__28043;
    wire N__28042;
    wire N__28039;
    wire N__28036;
    wire N__28033;
    wire N__28028;
    wire N__28027;
    wire N__28022;
    wire N__28019;
    wire N__28016;
    wire N__28013;
    wire N__28010;
    wire N__28007;
    wire N__28004;
    wire N__28001;
    wire N__27998;
    wire N__27995;
    wire N__27992;
    wire N__27989;
    wire N__27988;
    wire N__27987;
    wire N__27984;
    wire N__27979;
    wire N__27974;
    wire N__27971;
    wire N__27970;
    wire N__27969;
    wire N__27964;
    wire N__27961;
    wire N__27958;
    wire N__27953;
    wire N__27950;
    wire N__27947;
    wire N__27944;
    wire N__27941;
    wire N__27940;
    wire N__27935;
    wire N__27932;
    wire N__27931;
    wire N__27928;
    wire N__27923;
    wire N__27922;
    wire N__27919;
    wire N__27916;
    wire N__27913;
    wire N__27908;
    wire N__27905;
    wire N__27902;
    wire N__27899;
    wire N__27898;
    wire N__27897;
    wire N__27896;
    wire N__27889;
    wire N__27886;
    wire N__27883;
    wire N__27878;
    wire N__27875;
    wire N__27872;
    wire N__27871;
    wire N__27870;
    wire N__27867;
    wire N__27864;
    wire N__27857;
    wire N__27856;
    wire N__27853;
    wire N__27850;
    wire N__27847;
    wire N__27842;
    wire N__27839;
    wire N__27836;
    wire N__27835;
    wire N__27834;
    wire N__27831;
    wire N__27828;
    wire N__27825;
    wire N__27818;
    wire N__27815;
    wire N__27814;
    wire N__27813;
    wire N__27810;
    wire N__27807;
    wire N__27804;
    wire N__27799;
    wire N__27794;
    wire N__27793;
    wire N__27790;
    wire N__27787;
    wire N__27784;
    wire N__27781;
    wire N__27776;
    wire N__27775;
    wire N__27774;
    wire N__27769;
    wire N__27766;
    wire N__27763;
    wire N__27758;
    wire N__27755;
    wire N__27752;
    wire N__27749;
    wire N__27746;
    wire N__27743;
    wire N__27740;
    wire N__27739;
    wire N__27736;
    wire N__27735;
    wire N__27732;
    wire N__27729;
    wire N__27726;
    wire N__27723;
    wire N__27720;
    wire N__27713;
    wire N__27710;
    wire N__27709;
    wire N__27706;
    wire N__27703;
    wire N__27702;
    wire N__27699;
    wire N__27696;
    wire N__27693;
    wire N__27690;
    wire N__27687;
    wire N__27680;
    wire N__27677;
    wire N__27676;
    wire N__27673;
    wire N__27668;
    wire N__27667;
    wire N__27664;
    wire N__27661;
    wire N__27658;
    wire N__27653;
    wire N__27650;
    wire N__27649;
    wire N__27646;
    wire N__27643;
    wire N__27638;
    wire N__27635;
    wire N__27634;
    wire N__27631;
    wire N__27628;
    wire N__27623;
    wire N__27620;
    wire N__27619;
    wire N__27616;
    wire N__27613;
    wire N__27608;
    wire N__27605;
    wire N__27604;
    wire N__27601;
    wire N__27598;
    wire N__27593;
    wire N__27590;
    wire N__27589;
    wire N__27586;
    wire N__27583;
    wire N__27578;
    wire N__27575;
    wire N__27574;
    wire N__27571;
    wire N__27568;
    wire N__27563;
    wire N__27560;
    wire N__27557;
    wire N__27554;
    wire N__27553;
    wire N__27550;
    wire N__27549;
    wire N__27544;
    wire N__27541;
    wire N__27538;
    wire N__27533;
    wire N__27530;
    wire N__27529;
    wire N__27526;
    wire N__27523;
    wire N__27518;
    wire N__27515;
    wire N__27512;
    wire N__27509;
    wire N__27506;
    wire N__27503;
    wire N__27502;
    wire N__27499;
    wire N__27496;
    wire N__27491;
    wire N__27488;
    wire N__27487;
    wire N__27484;
    wire N__27481;
    wire N__27476;
    wire N__27473;
    wire N__27472;
    wire N__27469;
    wire N__27466;
    wire N__27461;
    wire N__27458;
    wire N__27457;
    wire N__27454;
    wire N__27451;
    wire N__27446;
    wire N__27443;
    wire N__27442;
    wire N__27439;
    wire N__27436;
    wire N__27431;
    wire N__27428;
    wire N__27427;
    wire N__27424;
    wire N__27421;
    wire N__27416;
    wire N__27413;
    wire N__27412;
    wire N__27409;
    wire N__27406;
    wire N__27401;
    wire N__27398;
    wire N__27395;
    wire N__27392;
    wire N__27389;
    wire N__27386;
    wire N__27383;
    wire N__27380;
    wire N__27377;
    wire N__27374;
    wire N__27371;
    wire N__27368;
    wire N__27365;
    wire N__27362;
    wire N__27359;
    wire N__27356;
    wire N__27353;
    wire N__27350;
    wire N__27347;
    wire N__27344;
    wire N__27341;
    wire N__27340;
    wire N__27335;
    wire N__27332;
    wire N__27329;
    wire N__27328;
    wire N__27327;
    wire N__27324;
    wire N__27321;
    wire N__27318;
    wire N__27315;
    wire N__27312;
    wire N__27305;
    wire N__27302;
    wire N__27301;
    wire N__27298;
    wire N__27297;
    wire N__27296;
    wire N__27293;
    wire N__27290;
    wire N__27285;
    wire N__27282;
    wire N__27277;
    wire N__27274;
    wire N__27271;
    wire N__27266;
    wire N__27263;
    wire N__27260;
    wire N__27257;
    wire N__27254;
    wire N__27251;
    wire N__27248;
    wire N__27245;
    wire N__27242;
    wire N__27239;
    wire N__27236;
    wire N__27233;
    wire N__27230;
    wire N__27227;
    wire N__27224;
    wire N__27221;
    wire N__27218;
    wire N__27215;
    wire N__27212;
    wire N__27209;
    wire N__27206;
    wire N__27203;
    wire N__27200;
    wire N__27197;
    wire N__27194;
    wire N__27191;
    wire N__27190;
    wire N__27189;
    wire N__27184;
    wire N__27181;
    wire N__27180;
    wire N__27177;
    wire N__27174;
    wire N__27171;
    wire N__27168;
    wire N__27163;
    wire N__27158;
    wire N__27155;
    wire N__27154;
    wire N__27149;
    wire N__27148;
    wire N__27145;
    wire N__27142;
    wire N__27137;
    wire N__27134;
    wire N__27131;
    wire N__27128;
    wire N__27127;
    wire N__27126;
    wire N__27123;
    wire N__27120;
    wire N__27119;
    wire N__27116;
    wire N__27113;
    wire N__27110;
    wire N__27107;
    wire N__27104;
    wire N__27097;
    wire N__27094;
    wire N__27091;
    wire N__27086;
    wire N__27085;
    wire N__27084;
    wire N__27081;
    wire N__27078;
    wire N__27075;
    wire N__27072;
    wire N__27069;
    wire N__27066;
    wire N__27063;
    wire N__27056;
    wire N__27055;
    wire N__27052;
    wire N__27051;
    wire N__27048;
    wire N__27045;
    wire N__27044;
    wire N__27041;
    wire N__27038;
    wire N__27035;
    wire N__27032;
    wire N__27029;
    wire N__27022;
    wire N__27019;
    wire N__27016;
    wire N__27011;
    wire N__27010;
    wire N__27009;
    wire N__27006;
    wire N__27003;
    wire N__27000;
    wire N__26993;
    wire N__26992;
    wire N__26989;
    wire N__26988;
    wire N__26987;
    wire N__26986;
    wire N__26985;
    wire N__26984;
    wire N__26983;
    wire N__26982;
    wire N__26981;
    wire N__26978;
    wire N__26977;
    wire N__26976;
    wire N__26973;
    wire N__26966;
    wire N__26965;
    wire N__26964;
    wire N__26961;
    wire N__26958;
    wire N__26951;
    wire N__26948;
    wire N__26943;
    wire N__26942;
    wire N__26941;
    wire N__26940;
    wire N__26939;
    wire N__26938;
    wire N__26937;
    wire N__26936;
    wire N__26931;
    wire N__26926;
    wire N__26923;
    wire N__26922;
    wire N__26921;
    wire N__26912;
    wire N__26911;
    wire N__26910;
    wire N__26895;
    wire N__26890;
    wire N__26887;
    wire N__26884;
    wire N__26881;
    wire N__26878;
    wire N__26873;
    wire N__26866;
    wire N__26855;
    wire N__26852;
    wire N__26849;
    wire N__26846;
    wire N__26843;
    wire N__26840;
    wire N__26837;
    wire N__26834;
    wire N__26833;
    wire N__26832;
    wire N__26831;
    wire N__26830;
    wire N__26829;
    wire N__26828;
    wire N__26827;
    wire N__26826;
    wire N__26825;
    wire N__26824;
    wire N__26823;
    wire N__26822;
    wire N__26821;
    wire N__26820;
    wire N__26819;
    wire N__26818;
    wire N__26801;
    wire N__26784;
    wire N__26781;
    wire N__26780;
    wire N__26775;
    wire N__26772;
    wire N__26769;
    wire N__26766;
    wire N__26763;
    wire N__26760;
    wire N__26757;
    wire N__26754;
    wire N__26751;
    wire N__26748;
    wire N__26743;
    wire N__26738;
    wire N__26735;
    wire N__26732;
    wire N__26729;
    wire N__26726;
    wire N__26723;
    wire N__26720;
    wire N__26717;
    wire N__26714;
    wire N__26711;
    wire N__26708;
    wire N__26705;
    wire N__26702;
    wire N__26699;
    wire N__26696;
    wire N__26693;
    wire N__26690;
    wire N__26687;
    wire N__26684;
    wire N__26681;
    wire N__26678;
    wire N__26675;
    wire N__26672;
    wire N__26669;
    wire N__26666;
    wire N__26663;
    wire N__26660;
    wire N__26657;
    wire N__26654;
    wire N__26651;
    wire N__26648;
    wire N__26647;
    wire N__26644;
    wire N__26643;
    wire N__26642;
    wire N__26639;
    wire N__26636;
    wire N__26633;
    wire N__26630;
    wire N__26625;
    wire N__26620;
    wire N__26617;
    wire N__26614;
    wire N__26609;
    wire N__26606;
    wire N__26605;
    wire N__26604;
    wire N__26599;
    wire N__26596;
    wire N__26591;
    wire N__26588;
    wire N__26585;
    wire N__26582;
    wire N__26579;
    wire N__26576;
    wire N__26573;
    wire N__26570;
    wire N__26567;
    wire N__26566;
    wire N__26563;
    wire N__26560;
    wire N__26557;
    wire N__26554;
    wire N__26551;
    wire N__26550;
    wire N__26549;
    wire N__26546;
    wire N__26543;
    wire N__26538;
    wire N__26531;
    wire N__26528;
    wire N__26527;
    wire N__26526;
    wire N__26523;
    wire N__26520;
    wire N__26517;
    wire N__26514;
    wire N__26507;
    wire N__26504;
    wire N__26501;
    wire N__26498;
    wire N__26495;
    wire N__26492;
    wire N__26489;
    wire N__26486;
    wire N__26483;
    wire N__26480;
    wire N__26477;
    wire N__26474;
    wire N__26471;
    wire N__26468;
    wire N__26465;
    wire N__26462;
    wire N__26459;
    wire N__26456;
    wire N__26453;
    wire N__26450;
    wire N__26447;
    wire N__26444;
    wire N__26441;
    wire N__26438;
    wire N__26435;
    wire N__26432;
    wire N__26429;
    wire N__26426;
    wire N__26423;
    wire N__26420;
    wire N__26417;
    wire N__26414;
    wire N__26411;
    wire N__26408;
    wire N__26405;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26393;
    wire N__26390;
    wire N__26387;
    wire N__26384;
    wire N__26381;
    wire N__26378;
    wire N__26375;
    wire N__26372;
    wire N__26369;
    wire N__26366;
    wire N__26363;
    wire N__26360;
    wire N__26357;
    wire N__26354;
    wire N__26351;
    wire N__26348;
    wire N__26345;
    wire N__26342;
    wire N__26339;
    wire N__26336;
    wire N__26333;
    wire N__26330;
    wire N__26327;
    wire N__26324;
    wire N__26321;
    wire N__26318;
    wire N__26315;
    wire N__26312;
    wire N__26309;
    wire N__26306;
    wire N__26303;
    wire N__26300;
    wire N__26297;
    wire N__26294;
    wire N__26291;
    wire N__26288;
    wire N__26285;
    wire N__26282;
    wire N__26279;
    wire N__26276;
    wire N__26273;
    wire N__26270;
    wire N__26267;
    wire N__26264;
    wire N__26261;
    wire N__26258;
    wire N__26255;
    wire N__26252;
    wire N__26249;
    wire N__26246;
    wire N__26243;
    wire N__26240;
    wire N__26237;
    wire N__26236;
    wire N__26233;
    wire N__26232;
    wire N__26229;
    wire N__26222;
    wire N__26221;
    wire N__26218;
    wire N__26215;
    wire N__26212;
    wire N__26207;
    wire N__26204;
    wire N__26203;
    wire N__26202;
    wire N__26201;
    wire N__26200;
    wire N__26199;
    wire N__26198;
    wire N__26197;
    wire N__26196;
    wire N__26195;
    wire N__26194;
    wire N__26193;
    wire N__26192;
    wire N__26189;
    wire N__26186;
    wire N__26177;
    wire N__26170;
    wire N__26161;
    wire N__26160;
    wire N__26159;
    wire N__26158;
    wire N__26157;
    wire N__26156;
    wire N__26155;
    wire N__26154;
    wire N__26153;
    wire N__26152;
    wire N__26151;
    wire N__26150;
    wire N__26149;
    wire N__26148;
    wire N__26147;
    wire N__26146;
    wire N__26145;
    wire N__26144;
    wire N__26143;
    wire N__26142;
    wire N__26139;
    wire N__26130;
    wire N__26121;
    wire N__26112;
    wire N__26103;
    wire N__26094;
    wire N__26087;
    wire N__26084;
    wire N__26081;
    wire N__26070;
    wire N__26067;
    wire N__26062;
    wire N__26059;
    wire N__26056;
    wire N__26053;
    wire N__26048;
    wire N__26045;
    wire N__26044;
    wire N__26041;
    wire N__26040;
    wire N__26033;
    wire N__26032;
    wire N__26029;
    wire N__26026;
    wire N__26023;
    wire N__26018;
    wire N__26015;
    wire N__26012;
    wire N__26009;
    wire N__26006;
    wire N__26003;
    wire N__26000;
    wire N__25997;
    wire N__25996;
    wire N__25993;
    wire N__25990;
    wire N__25987;
    wire N__25984;
    wire N__25983;
    wire N__25978;
    wire N__25975;
    wire N__25972;
    wire N__25967;
    wire N__25964;
    wire N__25963;
    wire N__25960;
    wire N__25957;
    wire N__25956;
    wire N__25951;
    wire N__25948;
    wire N__25945;
    wire N__25940;
    wire N__25937;
    wire N__25936;
    wire N__25931;
    wire N__25930;
    wire N__25927;
    wire N__25924;
    wire N__25921;
    wire N__25916;
    wire N__25913;
    wire N__25912;
    wire N__25909;
    wire N__25904;
    wire N__25903;
    wire N__25900;
    wire N__25897;
    wire N__25894;
    wire N__25889;
    wire N__25886;
    wire N__25885;
    wire N__25882;
    wire N__25877;
    wire N__25876;
    wire N__25873;
    wire N__25870;
    wire N__25867;
    wire N__25862;
    wire N__25859;
    wire N__25858;
    wire N__25853;
    wire N__25852;
    wire N__25849;
    wire N__25846;
    wire N__25843;
    wire N__25838;
    wire N__25835;
    wire N__25832;
    wire N__25829;
    wire N__25826;
    wire N__25825;
    wire N__25822;
    wire N__25819;
    wire N__25816;
    wire N__25811;
    wire N__25808;
    wire N__25807;
    wire N__25804;
    wire N__25801;
    wire N__25798;
    wire N__25793;
    wire N__25790;
    wire N__25789;
    wire N__25786;
    wire N__25783;
    wire N__25780;
    wire N__25775;
    wire N__25772;
    wire N__25771;
    wire N__25768;
    wire N__25765;
    wire N__25762;
    wire N__25757;
    wire N__25754;
    wire N__25753;
    wire N__25750;
    wire N__25747;
    wire N__25744;
    wire N__25739;
    wire N__25736;
    wire N__25735;
    wire N__25732;
    wire N__25729;
    wire N__25726;
    wire N__25721;
    wire N__25718;
    wire N__25717;
    wire N__25716;
    wire N__25713;
    wire N__25708;
    wire N__25703;
    wire N__25700;
    wire N__25699;
    wire N__25698;
    wire N__25695;
    wire N__25690;
    wire N__25685;
    wire N__25682;
    wire N__25681;
    wire N__25678;
    wire N__25675;
    wire N__25672;
    wire N__25667;
    wire N__25664;
    wire N__25661;
    wire N__25658;
    wire N__25655;
    wire N__25654;
    wire N__25651;
    wire N__25648;
    wire N__25645;
    wire N__25640;
    wire N__25637;
    wire N__25634;
    wire N__25633;
    wire N__25630;
    wire N__25627;
    wire N__25624;
    wire N__25619;
    wire N__25616;
    wire N__25615;
    wire N__25612;
    wire N__25609;
    wire N__25606;
    wire N__25601;
    wire N__25598;
    wire N__25597;
    wire N__25594;
    wire N__25591;
    wire N__25588;
    wire N__25583;
    wire N__25580;
    wire N__25577;
    wire N__25576;
    wire N__25573;
    wire N__25570;
    wire N__25567;
    wire N__25562;
    wire N__25559;
    wire N__25558;
    wire N__25555;
    wire N__25552;
    wire N__25549;
    wire N__25544;
    wire N__25541;
    wire N__25540;
    wire N__25537;
    wire N__25534;
    wire N__25531;
    wire N__25526;
    wire N__25523;
    wire N__25520;
    wire N__25517;
    wire N__25514;
    wire N__25511;
    wire N__25508;
    wire N__25505;
    wire N__25502;
    wire N__25499;
    wire N__25496;
    wire N__25493;
    wire N__25490;
    wire N__25487;
    wire N__25484;
    wire N__25481;
    wire N__25478;
    wire N__25475;
    wire N__25472;
    wire N__25469;
    wire N__25466;
    wire N__25463;
    wire N__25460;
    wire N__25459;
    wire N__25456;
    wire N__25453;
    wire N__25448;
    wire N__25445;
    wire N__25442;
    wire N__25439;
    wire N__25436;
    wire N__25433;
    wire N__25430;
    wire N__25427;
    wire N__25424;
    wire N__25421;
    wire N__25420;
    wire N__25417;
    wire N__25416;
    wire N__25413;
    wire N__25410;
    wire N__25407;
    wire N__25400;
    wire N__25397;
    wire N__25394;
    wire N__25391;
    wire N__25388;
    wire N__25385;
    wire N__25382;
    wire N__25379;
    wire N__25376;
    wire N__25373;
    wire N__25370;
    wire N__25367;
    wire N__25364;
    wire N__25361;
    wire N__25358;
    wire N__25355;
    wire N__25352;
    wire N__25349;
    wire N__25346;
    wire N__25343;
    wire N__25340;
    wire N__25337;
    wire N__25334;
    wire N__25331;
    wire N__25328;
    wire N__25325;
    wire N__25322;
    wire N__25319;
    wire N__25316;
    wire N__25313;
    wire N__25310;
    wire N__25307;
    wire N__25304;
    wire N__25301;
    wire N__25298;
    wire N__25295;
    wire N__25292;
    wire N__25289;
    wire N__25286;
    wire N__25283;
    wire N__25280;
    wire N__25277;
    wire N__25274;
    wire N__25271;
    wire N__25268;
    wire N__25265;
    wire N__25262;
    wire N__25259;
    wire N__25256;
    wire N__25253;
    wire N__25250;
    wire N__25247;
    wire N__25244;
    wire N__25241;
    wire N__25238;
    wire N__25235;
    wire N__25232;
    wire N__25229;
    wire N__25226;
    wire N__25223;
    wire N__25220;
    wire N__25217;
    wire N__25214;
    wire N__25211;
    wire N__25208;
    wire N__25205;
    wire N__25202;
    wire N__25199;
    wire N__25196;
    wire N__25193;
    wire N__25190;
    wire N__25187;
    wire N__25184;
    wire N__25181;
    wire N__25178;
    wire N__25175;
    wire N__25172;
    wire N__25169;
    wire N__25166;
    wire N__25165;
    wire N__25164;
    wire N__25161;
    wire N__25158;
    wire N__25155;
    wire N__25154;
    wire N__25149;
    wire N__25146;
    wire N__25143;
    wire N__25140;
    wire N__25137;
    wire N__25134;
    wire N__25127;
    wire N__25124;
    wire N__25123;
    wire N__25122;
    wire N__25119;
    wire N__25116;
    wire N__25113;
    wire N__25108;
    wire N__25103;
    wire N__25102;
    wire N__25101;
    wire N__25098;
    wire N__25095;
    wire N__25092;
    wire N__25089;
    wire N__25084;
    wire N__25081;
    wire N__25080;
    wire N__25077;
    wire N__25074;
    wire N__25071;
    wire N__25068;
    wire N__25063;
    wire N__25058;
    wire N__25057;
    wire N__25054;
    wire N__25053;
    wire N__25050;
    wire N__25047;
    wire N__25044;
    wire N__25037;
    wire N__25036;
    wire N__25035;
    wire N__25028;
    wire N__25025;
    wire N__25022;
    wire N__25021;
    wire N__25020;
    wire N__25013;
    wire N__25010;
    wire N__25007;
    wire N__25004;
    wire N__25001;
    wire N__24998;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24986;
    wire N__24983;
    wire N__24980;
    wire N__24977;
    wire N__24974;
    wire N__24971;
    wire N__24968;
    wire N__24965;
    wire N__24962;
    wire N__24959;
    wire N__24956;
    wire N__24953;
    wire N__24952;
    wire N__24947;
    wire N__24944;
    wire N__24941;
    wire N__24938;
    wire N__24937;
    wire N__24934;
    wire N__24931;
    wire N__24926;
    wire N__24923;
    wire N__24922;
    wire N__24917;
    wire N__24916;
    wire N__24913;
    wire N__24910;
    wire N__24909;
    wire N__24906;
    wire N__24903;
    wire N__24900;
    wire N__24895;
    wire N__24890;
    wire N__24887;
    wire N__24884;
    wire N__24881;
    wire N__24878;
    wire N__24875;
    wire N__24872;
    wire N__24869;
    wire N__24866;
    wire N__24863;
    wire N__24860;
    wire N__24857;
    wire N__24854;
    wire N__24851;
    wire N__24848;
    wire N__24845;
    wire N__24842;
    wire N__24839;
    wire N__24836;
    wire N__24833;
    wire N__24830;
    wire N__24827;
    wire N__24824;
    wire N__24821;
    wire N__24818;
    wire N__24815;
    wire N__24812;
    wire N__24809;
    wire N__24806;
    wire N__24803;
    wire N__24800;
    wire N__24797;
    wire N__24794;
    wire N__24791;
    wire N__24788;
    wire N__24787;
    wire N__24786;
    wire N__24783;
    wire N__24780;
    wire N__24777;
    wire N__24774;
    wire N__24769;
    wire N__24766;
    wire N__24763;
    wire N__24758;
    wire N__24755;
    wire N__24752;
    wire N__24749;
    wire N__24746;
    wire N__24743;
    wire N__24740;
    wire N__24737;
    wire N__24734;
    wire N__24731;
    wire N__24728;
    wire N__24725;
    wire N__24722;
    wire N__24719;
    wire N__24716;
    wire N__24713;
    wire N__24710;
    wire N__24707;
    wire N__24704;
    wire N__24701;
    wire N__24698;
    wire N__24697;
    wire N__24696;
    wire N__24693;
    wire N__24690;
    wire N__24687;
    wire N__24684;
    wire N__24679;
    wire N__24674;
    wire N__24671;
    wire N__24668;
    wire N__24665;
    wire N__24662;
    wire N__24659;
    wire N__24656;
    wire N__24653;
    wire N__24650;
    wire N__24647;
    wire N__24644;
    wire N__24641;
    wire N__24638;
    wire N__24635;
    wire N__24632;
    wire N__24629;
    wire N__24626;
    wire N__24623;
    wire N__24620;
    wire N__24619;
    wire N__24618;
    wire N__24615;
    wire N__24610;
    wire N__24605;
    wire N__24602;
    wire N__24599;
    wire N__24596;
    wire N__24593;
    wire N__24590;
    wire N__24587;
    wire N__24584;
    wire N__24581;
    wire N__24578;
    wire N__24575;
    wire N__24572;
    wire N__24569;
    wire N__24568;
    wire N__24567;
    wire N__24560;
    wire N__24557;
    wire N__24554;
    wire N__24551;
    wire N__24548;
    wire N__24545;
    wire N__24542;
    wire N__24539;
    wire N__24536;
    wire N__24533;
    wire N__24530;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24518;
    wire N__24515;
    wire N__24512;
    wire N__24509;
    wire N__24506;
    wire N__24503;
    wire N__24500;
    wire N__24499;
    wire N__24496;
    wire N__24493;
    wire N__24490;
    wire N__24487;
    wire N__24484;
    wire N__24483;
    wire N__24478;
    wire N__24475;
    wire N__24470;
    wire N__24467;
    wire N__24464;
    wire N__24461;
    wire N__24458;
    wire N__24455;
    wire N__24452;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24440;
    wire N__24437;
    wire N__24436;
    wire N__24435;
    wire N__24432;
    wire N__24427;
    wire N__24422;
    wire N__24421;
    wire N__24418;
    wire N__24415;
    wire N__24412;
    wire N__24409;
    wire N__24404;
    wire N__24401;
    wire N__24398;
    wire N__24395;
    wire N__24394;
    wire N__24391;
    wire N__24388;
    wire N__24387;
    wire N__24382;
    wire N__24379;
    wire N__24378;
    wire N__24375;
    wire N__24372;
    wire N__24369;
    wire N__24366;
    wire N__24361;
    wire N__24356;
    wire N__24353;
    wire N__24350;
    wire N__24347;
    wire N__24344;
    wire N__24341;
    wire N__24338;
    wire N__24335;
    wire N__24332;
    wire N__24329;
    wire N__24326;
    wire N__24323;
    wire N__24320;
    wire N__24317;
    wire N__24314;
    wire N__24311;
    wire N__24308;
    wire N__24305;
    wire N__24302;
    wire N__24299;
    wire N__24296;
    wire N__24293;
    wire N__24290;
    wire N__24287;
    wire N__24284;
    wire N__24283;
    wire N__24282;
    wire N__24279;
    wire N__24276;
    wire N__24273;
    wire N__24270;
    wire N__24263;
    wire N__24262;
    wire N__24259;
    wire N__24256;
    wire N__24253;
    wire N__24250;
    wire N__24249;
    wire N__24246;
    wire N__24243;
    wire N__24240;
    wire N__24237;
    wire N__24232;
    wire N__24231;
    wire N__24228;
    wire N__24225;
    wire N__24222;
    wire N__24215;
    wire N__24212;
    wire N__24209;
    wire N__24206;
    wire N__24203;
    wire N__24200;
    wire N__24197;
    wire N__24194;
    wire N__24191;
    wire N__24188;
    wire N__24187;
    wire N__24186;
    wire N__24185;
    wire N__24178;
    wire N__24175;
    wire N__24170;
    wire N__24167;
    wire N__24164;
    wire N__24161;
    wire N__24158;
    wire N__24155;
    wire N__24152;
    wire N__24149;
    wire N__24148;
    wire N__24147;
    wire N__24144;
    wire N__24139;
    wire N__24136;
    wire N__24135;
    wire N__24132;
    wire N__24129;
    wire N__24126;
    wire N__24123;
    wire N__24118;
    wire N__24113;
    wire N__24110;
    wire N__24107;
    wire N__24104;
    wire N__24101;
    wire N__24098;
    wire N__24097;
    wire N__24092;
    wire N__24089;
    wire N__24086;
    wire N__24085;
    wire N__24082;
    wire N__24079;
    wire N__24074;
    wire N__24071;
    wire N__24068;
    wire N__24065;
    wire N__24062;
    wire N__24059;
    wire N__24058;
    wire N__24057;
    wire N__24054;
    wire N__24051;
    wire N__24048;
    wire N__24043;
    wire N__24042;
    wire N__24037;
    wire N__24034;
    wire N__24029;
    wire N__24026;
    wire N__24023;
    wire N__24022;
    wire N__24021;
    wire N__24018;
    wire N__24015;
    wire N__24012;
    wire N__24009;
    wire N__24006;
    wire N__24005;
    wire N__24000;
    wire N__23997;
    wire N__23994;
    wire N__23991;
    wire N__23986;
    wire N__23981;
    wire N__23978;
    wire N__23975;
    wire N__23972;
    wire N__23969;
    wire N__23966;
    wire N__23963;
    wire N__23960;
    wire N__23957;
    wire N__23956;
    wire N__23955;
    wire N__23952;
    wire N__23949;
    wire N__23946;
    wire N__23939;
    wire N__23938;
    wire N__23937;
    wire N__23934;
    wire N__23933;
    wire N__23930;
    wire N__23927;
    wire N__23924;
    wire N__23921;
    wire N__23918;
    wire N__23915;
    wire N__23912;
    wire N__23909;
    wire N__23904;
    wire N__23899;
    wire N__23896;
    wire N__23891;
    wire N__23888;
    wire N__23885;
    wire N__23884;
    wire N__23883;
    wire N__23880;
    wire N__23877;
    wire N__23874;
    wire N__23869;
    wire N__23864;
    wire N__23863;
    wire N__23860;
    wire N__23857;
    wire N__23856;
    wire N__23853;
    wire N__23852;
    wire N__23849;
    wire N__23846;
    wire N__23843;
    wire N__23840;
    wire N__23831;
    wire N__23828;
    wire N__23825;
    wire N__23822;
    wire N__23819;
    wire N__23816;
    wire N__23813;
    wire N__23810;
    wire N__23807;
    wire N__23804;
    wire N__23801;
    wire N__23800;
    wire N__23797;
    wire N__23794;
    wire N__23789;
    wire N__23788;
    wire N__23787;
    wire N__23780;
    wire N__23777;
    wire N__23776;
    wire N__23775;
    wire N__23768;
    wire N__23765;
    wire N__23762;
    wire N__23759;
    wire N__23756;
    wire N__23753;
    wire N__23752;
    wire N__23749;
    wire N__23746;
    wire N__23741;
    wire N__23738;
    wire N__23737;
    wire N__23736;
    wire N__23733;
    wire N__23730;
    wire N__23727;
    wire N__23724;
    wire N__23721;
    wire N__23714;
    wire N__23713;
    wire N__23710;
    wire N__23707;
    wire N__23704;
    wire N__23703;
    wire N__23700;
    wire N__23699;
    wire N__23696;
    wire N__23693;
    wire N__23690;
    wire N__23687;
    wire N__23678;
    wire N__23677;
    wire N__23674;
    wire N__23671;
    wire N__23670;
    wire N__23667;
    wire N__23664;
    wire N__23661;
    wire N__23656;
    wire N__23651;
    wire N__23650;
    wire N__23647;
    wire N__23644;
    wire N__23643;
    wire N__23640;
    wire N__23637;
    wire N__23636;
    wire N__23633;
    wire N__23628;
    wire N__23625;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23611;
    wire N__23610;
    wire N__23607;
    wire N__23604;
    wire N__23601;
    wire N__23598;
    wire N__23591;
    wire N__23590;
    wire N__23589;
    wire N__23586;
    wire N__23583;
    wire N__23580;
    wire N__23579;
    wire N__23576;
    wire N__23571;
    wire N__23568;
    wire N__23565;
    wire N__23562;
    wire N__23559;
    wire N__23556;
    wire N__23551;
    wire N__23546;
    wire N__23543;
    wire N__23542;
    wire N__23537;
    wire N__23534;
    wire N__23533;
    wire N__23532;
    wire N__23529;
    wire N__23526;
    wire N__23523;
    wire N__23520;
    wire N__23513;
    wire N__23512;
    wire N__23511;
    wire N__23510;
    wire N__23507;
    wire N__23504;
    wire N__23499;
    wire N__23496;
    wire N__23493;
    wire N__23490;
    wire N__23487;
    wire N__23484;
    wire N__23481;
    wire N__23474;
    wire N__23471;
    wire N__23468;
    wire N__23465;
    wire N__23464;
    wire N__23463;
    wire N__23460;
    wire N__23457;
    wire N__23454;
    wire N__23449;
    wire N__23446;
    wire N__23441;
    wire N__23440;
    wire N__23439;
    wire N__23436;
    wire N__23433;
    wire N__23432;
    wire N__23429;
    wire N__23426;
    wire N__23423;
    wire N__23420;
    wire N__23417;
    wire N__23412;
    wire N__23409;
    wire N__23406;
    wire N__23403;
    wire N__23400;
    wire N__23397;
    wire N__23392;
    wire N__23389;
    wire N__23384;
    wire N__23381;
    wire N__23380;
    wire N__23379;
    wire N__23376;
    wire N__23373;
    wire N__23370;
    wire N__23365;
    wire N__23360;
    wire N__23359;
    wire N__23354;
    wire N__23351;
    wire N__23350;
    wire N__23347;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23335;
    wire N__23332;
    wire N__23329;
    wire N__23324;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23309;
    wire N__23306;
    wire N__23303;
    wire N__23300;
    wire N__23297;
    wire N__23294;
    wire N__23293;
    wire N__23292;
    wire N__23289;
    wire N__23286;
    wire N__23283;
    wire N__23282;
    wire N__23277;
    wire N__23274;
    wire N__23271;
    wire N__23268;
    wire N__23265;
    wire N__23262;
    wire N__23259;
    wire N__23254;
    wire N__23249;
    wire N__23246;
    wire N__23243;
    wire N__23240;
    wire N__23239;
    wire N__23236;
    wire N__23235;
    wire N__23234;
    wire N__23231;
    wire N__23228;
    wire N__23223;
    wire N__23220;
    wire N__23213;
    wire N__23212;
    wire N__23209;
    wire N__23206;
    wire N__23201;
    wire N__23198;
    wire N__23197;
    wire N__23194;
    wire N__23191;
    wire N__23188;
    wire N__23185;
    wire N__23180;
    wire N__23179;
    wire N__23178;
    wire N__23175;
    wire N__23172;
    wire N__23169;
    wire N__23166;
    wire N__23163;
    wire N__23162;
    wire N__23159;
    wire N__23154;
    wire N__23151;
    wire N__23148;
    wire N__23145;
    wire N__23142;
    wire N__23135;
    wire N__23134;
    wire N__23133;
    wire N__23130;
    wire N__23127;
    wire N__23124;
    wire N__23117;
    wire N__23116;
    wire N__23115;
    wire N__23112;
    wire N__23109;
    wire N__23106;
    wire N__23099;
    wire N__23098;
    wire N__23097;
    wire N__23094;
    wire N__23093;
    wire N__23090;
    wire N__23087;
    wire N__23084;
    wire N__23081;
    wire N__23078;
    wire N__23069;
    wire N__23066;
    wire N__23065;
    wire N__23064;
    wire N__23061;
    wire N__23058;
    wire N__23055;
    wire N__23048;
    wire N__23045;
    wire N__23042;
    wire N__23041;
    wire N__23040;
    wire N__23039;
    wire N__23036;
    wire N__23033;
    wire N__23028;
    wire N__23021;
    wire N__23020;
    wire N__23019;
    wire N__23016;
    wire N__23013;
    wire N__23010;
    wire N__23003;
    wire N__23000;
    wire N__22999;
    wire N__22998;
    wire N__22997;
    wire N__22994;
    wire N__22991;
    wire N__22986;
    wire N__22979;
    wire N__22976;
    wire N__22973;
    wire N__22972;
    wire N__22971;
    wire N__22968;
    wire N__22965;
    wire N__22962;
    wire N__22957;
    wire N__22952;
    wire N__22949;
    wire N__22948;
    wire N__22945;
    wire N__22944;
    wire N__22941;
    wire N__22938;
    wire N__22935;
    wire N__22928;
    wire N__22925;
    wire N__22922;
    wire N__22921;
    wire N__22918;
    wire N__22915;
    wire N__22912;
    wire N__22909;
    wire N__22904;
    wire N__22901;
    wire N__22900;
    wire N__22897;
    wire N__22894;
    wire N__22891;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22876;
    wire N__22871;
    wire N__22868;
    wire N__22867;
    wire N__22864;
    wire N__22861;
    wire N__22858;
    wire N__22855;
    wire N__22850;
    wire N__22847;
    wire N__22846;
    wire N__22843;
    wire N__22840;
    wire N__22837;
    wire N__22834;
    wire N__22831;
    wire N__22828;
    wire N__22825;
    wire N__22822;
    wire N__22817;
    wire N__22814;
    wire N__22811;
    wire N__22808;
    wire N__22805;
    wire N__22804;
    wire N__22801;
    wire N__22798;
    wire N__22795;
    wire N__22792;
    wire N__22789;
    wire N__22786;
    wire N__22783;
    wire N__22780;
    wire N__22775;
    wire N__22772;
    wire N__22769;
    wire N__22766;
    wire N__22763;
    wire N__22760;
    wire N__22757;
    wire N__22754;
    wire N__22751;
    wire N__22748;
    wire N__22745;
    wire N__22742;
    wire N__22739;
    wire N__22736;
    wire N__22733;
    wire N__22730;
    wire N__22727;
    wire N__22724;
    wire N__22721;
    wire N__22718;
    wire N__22715;
    wire N__22712;
    wire N__22709;
    wire N__22706;
    wire N__22703;
    wire N__22700;
    wire N__22697;
    wire N__22694;
    wire N__22691;
    wire N__22688;
    wire N__22685;
    wire N__22682;
    wire N__22679;
    wire N__22676;
    wire N__22673;
    wire N__22670;
    wire N__22667;
    wire N__22664;
    wire N__22661;
    wire N__22658;
    wire N__22655;
    wire N__22652;
    wire N__22649;
    wire N__22646;
    wire N__22643;
    wire N__22640;
    wire N__22637;
    wire N__22636;
    wire N__22633;
    wire N__22630;
    wire N__22627;
    wire N__22622;
    wire N__22619;
    wire N__22616;
    wire N__22613;
    wire N__22610;
    wire N__22607;
    wire N__22604;
    wire N__22601;
    wire N__22598;
    wire N__22595;
    wire N__22592;
    wire N__22589;
    wire N__22586;
    wire N__22583;
    wire N__22580;
    wire N__22577;
    wire N__22574;
    wire N__22571;
    wire N__22568;
    wire N__22565;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22553;
    wire N__22550;
    wire N__22547;
    wire N__22544;
    wire N__22541;
    wire N__22538;
    wire N__22535;
    wire N__22532;
    wire N__22529;
    wire N__22526;
    wire N__22523;
    wire N__22520;
    wire N__22517;
    wire N__22514;
    wire N__22511;
    wire N__22510;
    wire N__22507;
    wire N__22504;
    wire N__22499;
    wire N__22496;
    wire N__22493;
    wire N__22490;
    wire N__22487;
    wire N__22484;
    wire N__22481;
    wire N__22478;
    wire N__22475;
    wire N__22472;
    wire N__22469;
    wire N__22466;
    wire N__22463;
    wire N__22460;
    wire N__22457;
    wire N__22454;
    wire N__22451;
    wire N__22448;
    wire N__22445;
    wire N__22442;
    wire N__22439;
    wire N__22436;
    wire N__22433;
    wire N__22430;
    wire N__22427;
    wire N__22424;
    wire N__22421;
    wire N__22418;
    wire N__22415;
    wire N__22412;
    wire N__22409;
    wire N__22406;
    wire N__22403;
    wire N__22400;
    wire N__22397;
    wire N__22394;
    wire N__22391;
    wire N__22388;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22376;
    wire N__22373;
    wire N__22370;
    wire N__22367;
    wire N__22364;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22346;
    wire N__22343;
    wire N__22340;
    wire N__22337;
    wire N__22334;
    wire N__22331;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22301;
    wire N__22298;
    wire N__22295;
    wire N__22292;
    wire N__22289;
    wire N__22286;
    wire N__22283;
    wire N__22280;
    wire N__22277;
    wire N__22274;
    wire N__22271;
    wire N__22268;
    wire N__22265;
    wire N__22262;
    wire N__22259;
    wire N__22256;
    wire N__22253;
    wire N__22250;
    wire N__22247;
    wire N__22244;
    wire N__22241;
    wire N__22238;
    wire N__22235;
    wire N__22232;
    wire N__22229;
    wire N__22226;
    wire N__22223;
    wire N__22220;
    wire N__22217;
    wire N__22214;
    wire N__22211;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22169;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22157;
    wire N__22154;
    wire N__22151;
    wire N__22148;
    wire N__22145;
    wire N__22142;
    wire N__22139;
    wire N__22136;
    wire N__22133;
    wire N__22130;
    wire N__22127;
    wire N__22124;
    wire N__22121;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22109;
    wire N__22106;
    wire N__22103;
    wire N__22100;
    wire N__22097;
    wire N__22094;
    wire N__22091;
    wire N__22088;
    wire N__22085;
    wire N__22082;
    wire N__22079;
    wire N__22076;
    wire N__22073;
    wire N__22070;
    wire N__22067;
    wire N__22064;
    wire N__22061;
    wire N__22058;
    wire N__22055;
    wire N__22052;
    wire N__22049;
    wire N__22046;
    wire N__22043;
    wire N__22040;
    wire N__22037;
    wire N__22034;
    wire N__22031;
    wire N__22028;
    wire N__22025;
    wire N__22022;
    wire N__22021;
    wire N__22018;
    wire N__22015;
    wire N__22012;
    wire N__22009;
    wire N__22004;
    wire N__22001;
    wire N__22000;
    wire N__21997;
    wire N__21994;
    wire N__21991;
    wire N__21988;
    wire N__21983;
    wire N__21982;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21965;
    wire N__21962;
    wire N__21959;
    wire N__21956;
    wire N__21955;
    wire N__21952;
    wire N__21951;
    wire N__21948;
    wire N__21945;
    wire N__21942;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21928;
    wire N__21927;
    wire N__21924;
    wire N__21921;
    wire N__21918;
    wire N__21915;
    wire N__21908;
    wire N__21905;
    wire N__21904;
    wire N__21901;
    wire N__21898;
    wire N__21893;
    wire N__21890;
    wire N__21887;
    wire N__21884;
    wire N__21881;
    wire N__21878;
    wire N__21875;
    wire N__21872;
    wire N__21869;
    wire N__21868;
    wire N__21867;
    wire N__21864;
    wire N__21861;
    wire N__21858;
    wire N__21851;
    wire N__21848;
    wire N__21847;
    wire N__21844;
    wire N__21843;
    wire N__21840;
    wire N__21837;
    wire N__21834;
    wire N__21827;
    wire N__21824;
    wire N__21823;
    wire N__21820;
    wire N__21819;
    wire N__21816;
    wire N__21813;
    wire N__21810;
    wire N__21803;
    wire N__21800;
    wire N__21799;
    wire N__21796;
    wire N__21795;
    wire N__21792;
    wire N__21789;
    wire N__21786;
    wire N__21779;
    wire N__21776;
    wire N__21775;
    wire N__21772;
    wire N__21771;
    wire N__21768;
    wire N__21765;
    wire N__21762;
    wire N__21755;
    wire N__21752;
    wire N__21751;
    wire N__21748;
    wire N__21747;
    wire N__21744;
    wire N__21741;
    wire N__21738;
    wire N__21731;
    wire N__21728;
    wire N__21727;
    wire N__21724;
    wire N__21723;
    wire N__21720;
    wire N__21717;
    wire N__21714;
    wire N__21707;
    wire N__21704;
    wire N__21703;
    wire N__21700;
    wire N__21699;
    wire N__21696;
    wire N__21693;
    wire N__21690;
    wire N__21683;
    wire N__21680;
    wire N__21679;
    wire N__21676;
    wire N__21673;
    wire N__21668;
    wire N__21665;
    wire N__21664;
    wire N__21661;
    wire N__21660;
    wire N__21657;
    wire N__21654;
    wire N__21651;
    wire N__21644;
    wire N__21641;
    wire N__21640;
    wire N__21637;
    wire N__21636;
    wire N__21633;
    wire N__21630;
    wire N__21627;
    wire N__21620;
    wire N__21617;
    wire N__21616;
    wire N__21613;
    wire N__21612;
    wire N__21609;
    wire N__21606;
    wire N__21603;
    wire N__21596;
    wire N__21593;
    wire N__21592;
    wire N__21589;
    wire N__21588;
    wire N__21585;
    wire N__21582;
    wire N__21579;
    wire N__21572;
    wire N__21569;
    wire N__21568;
    wire N__21565;
    wire N__21564;
    wire N__21561;
    wire N__21558;
    wire N__21555;
    wire N__21548;
    wire N__21545;
    wire N__21544;
    wire N__21541;
    wire N__21540;
    wire N__21537;
    wire N__21534;
    wire N__21531;
    wire N__21524;
    wire N__21521;
    wire N__21520;
    wire N__21517;
    wire N__21516;
    wire N__21513;
    wire N__21510;
    wire N__21507;
    wire N__21500;
    wire N__21497;
    wire N__21496;
    wire N__21493;
    wire N__21492;
    wire N__21489;
    wire N__21486;
    wire N__21483;
    wire N__21476;
    wire N__21473;
    wire N__21472;
    wire N__21469;
    wire N__21468;
    wire N__21465;
    wire N__21462;
    wire N__21459;
    wire N__21452;
    wire N__21451;
    wire N__21448;
    wire N__21447;
    wire N__21444;
    wire N__21441;
    wire N__21438;
    wire N__21431;
    wire N__21428;
    wire N__21427;
    wire N__21424;
    wire N__21423;
    wire N__21420;
    wire N__21417;
    wire N__21414;
    wire N__21407;
    wire N__21404;
    wire N__21403;
    wire N__21400;
    wire N__21399;
    wire N__21396;
    wire N__21393;
    wire N__21390;
    wire N__21383;
    wire N__21380;
    wire N__21379;
    wire N__21376;
    wire N__21375;
    wire N__21372;
    wire N__21369;
    wire N__21366;
    wire N__21359;
    wire N__21356;
    wire N__21355;
    wire N__21352;
    wire N__21351;
    wire N__21348;
    wire N__21345;
    wire N__21342;
    wire N__21335;
    wire N__21332;
    wire N__21331;
    wire N__21328;
    wire N__21327;
    wire N__21324;
    wire N__21321;
    wire N__21318;
    wire N__21311;
    wire N__21308;
    wire N__21307;
    wire N__21304;
    wire N__21303;
    wire N__21300;
    wire N__21297;
    wire N__21294;
    wire N__21287;
    wire N__21284;
    wire N__21283;
    wire N__21280;
    wire N__21279;
    wire N__21276;
    wire N__21273;
    wire N__21270;
    wire N__21263;
    wire N__21260;
    wire N__21257;
    wire N__21256;
    wire N__21255;
    wire N__21252;
    wire N__21249;
    wire N__21246;
    wire N__21239;
    wire N__21236;
    wire N__21233;
    wire N__21232;
    wire N__21231;
    wire N__21228;
    wire N__21225;
    wire N__21222;
    wire N__21217;
    wire N__21212;
    wire N__21209;
    wire N__21208;
    wire N__21207;
    wire N__21204;
    wire N__21201;
    wire N__21198;
    wire N__21193;
    wire N__21188;
    wire N__21185;
    wire N__21182;
    wire N__21179;
    wire N__21176;
    wire N__21173;
    wire N__21172;
    wire N__21169;
    wire N__21166;
    wire N__21165;
    wire N__21160;
    wire N__21157;
    wire N__21154;
    wire N__21149;
    wire N__21146;
    wire N__21145;
    wire N__21142;
    wire N__21139;
    wire N__21136;
    wire N__21131;
    wire N__21128;
    wire N__21127;
    wire N__21126;
    wire N__21123;
    wire N__21120;
    wire N__21117;
    wire N__21112;
    wire N__21107;
    wire N__21104;
    wire N__21103;
    wire N__21100;
    wire N__21097;
    wire N__21094;
    wire N__21089;
    wire N__21086;
    wire N__21085;
    wire N__21084;
    wire N__21081;
    wire N__21078;
    wire N__21075;
    wire N__21070;
    wire N__21065;
    wire N__21062;
    wire N__21059;
    wire N__21056;
    wire N__21053;
    wire N__21050;
    wire N__21049;
    wire N__21046;
    wire N__21043;
    wire N__21042;
    wire N__21037;
    wire N__21034;
    wire N__21031;
    wire N__21026;
    wire N__21023;
    wire N__21020;
    wire N__21019;
    wire N__21018;
    wire N__21015;
    wire N__21012;
    wire N__21009;
    wire N__21004;
    wire N__20999;
    wire N__20996;
    wire N__20995;
    wire N__20994;
    wire N__20989;
    wire N__20986;
    wire N__20983;
    wire N__20978;
    wire N__20975;
    wire N__20974;
    wire N__20973;
    wire N__20968;
    wire N__20965;
    wire N__20962;
    wire N__20957;
    wire N__20954;
    wire N__20953;
    wire N__20950;
    wire N__20949;
    wire N__20946;
    wire N__20943;
    wire N__20940;
    wire N__20935;
    wire N__20930;
    wire N__20927;
    wire N__20926;
    wire N__20923;
    wire N__20920;
    wire N__20915;
    wire N__20914;
    wire N__20911;
    wire N__20908;
    wire N__20905;
    wire N__20900;
    wire N__20897;
    wire N__20896;
    wire N__20893;
    wire N__20890;
    wire N__20889;
    wire N__20884;
    wire N__20881;
    wire N__20878;
    wire N__20873;
    wire N__20870;
    wire N__20867;
    wire N__20866;
    wire N__20863;
    wire N__20860;
    wire N__20859;
    wire N__20854;
    wire N__20851;
    wire N__20848;
    wire N__20843;
    wire N__20840;
    wire N__20837;
    wire N__20836;
    wire N__20833;
    wire N__20830;
    wire N__20829;
    wire N__20826;
    wire N__20823;
    wire N__20820;
    wire N__20815;
    wire N__20810;
    wire N__20807;
    wire N__20806;
    wire N__20801;
    wire N__20800;
    wire N__20797;
    wire N__20794;
    wire N__20791;
    wire N__20786;
    wire N__20783;
    wire N__20782;
    wire N__20781;
    wire N__20776;
    wire N__20773;
    wire N__20770;
    wire N__20765;
    wire N__20762;
    wire N__20761;
    wire N__20758;
    wire N__20755;
    wire N__20754;
    wire N__20749;
    wire N__20746;
    wire N__20743;
    wire N__20738;
    wire N__20735;
    wire N__20734;
    wire N__20731;
    wire N__20728;
    wire N__20727;
    wire N__20722;
    wire N__20719;
    wire N__20716;
    wire N__20711;
    wire N__20708;
    wire N__20705;
    wire N__20704;
    wire N__20701;
    wire N__20698;
    wire N__20697;
    wire N__20692;
    wire N__20689;
    wire N__20686;
    wire N__20681;
    wire N__20678;
    wire N__20675;
    wire N__20674;
    wire N__20671;
    wire N__20668;
    wire N__20667;
    wire N__20662;
    wire N__20659;
    wire N__20656;
    wire N__20651;
    wire N__20648;
    wire N__20645;
    wire N__20644;
    wire N__20643;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20629;
    wire N__20624;
    wire N__20621;
    wire N__20618;
    wire N__20617;
    wire N__20614;
    wire N__20611;
    wire N__20608;
    wire N__20607;
    wire N__20602;
    wire N__20599;
    wire N__20596;
    wire N__20591;
    wire N__20588;
    wire N__20587;
    wire N__20582;
    wire N__20581;
    wire N__20578;
    wire N__20575;
    wire N__20572;
    wire N__20567;
    wire N__20564;
    wire N__20563;
    wire N__20560;
    wire N__20557;
    wire N__20556;
    wire N__20551;
    wire N__20548;
    wire N__20545;
    wire N__20540;
    wire N__20537;
    wire N__20536;
    wire N__20533;
    wire N__20530;
    wire N__20529;
    wire N__20524;
    wire N__20521;
    wire N__20518;
    wire N__20513;
    wire N__20510;
    wire N__20509;
    wire N__20504;
    wire N__20503;
    wire N__20500;
    wire N__20497;
    wire N__20494;
    wire N__20489;
    wire N__20486;
    wire N__20485;
    wire N__20480;
    wire N__20479;
    wire N__20476;
    wire N__20473;
    wire N__20470;
    wire N__20465;
    wire N__20462;
    wire N__20461;
    wire N__20458;
    wire N__20455;
    wire N__20452;
    wire N__20449;
    wire N__20448;
    wire N__20443;
    wire N__20440;
    wire N__20437;
    wire N__20432;
    wire N__20431;
    wire N__20430;
    wire N__20427;
    wire N__20424;
    wire N__20421;
    wire N__20418;
    wire N__20415;
    wire N__20414;
    wire N__20411;
    wire N__20406;
    wire N__20403;
    wire N__20396;
    wire N__20393;
    wire N__20390;
    wire N__20387;
    wire N__20384;
    wire N__20381;
    wire N__20378;
    wire N__20375;
    wire N__20372;
    wire N__20369;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20330;
    wire N__20327;
    wire N__20324;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20312;
    wire N__20309;
    wire N__20308;
    wire N__20305;
    wire N__20302;
    wire N__20299;
    wire N__20296;
    wire N__20293;
    wire N__20290;
    wire N__20287;
    wire N__20282;
    wire N__20279;
    wire N__20276;
    wire N__20273;
    wire N__20270;
    wire N__20267;
    wire N__20264;
    wire N__20261;
    wire N__20258;
    wire N__20255;
    wire N__20252;
    wire N__20249;
    wire N__20246;
    wire N__20243;
    wire N__20240;
    wire N__20237;
    wire N__20234;
    wire N__20231;
    wire N__20228;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20213;
    wire N__20210;
    wire N__20207;
    wire N__20204;
    wire N__20201;
    wire N__20198;
    wire N__20195;
    wire N__20192;
    wire N__20189;
    wire N__20186;
    wire N__20183;
    wire N__20180;
    wire N__20177;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20165;
    wire N__20162;
    wire N__20159;
    wire N__20156;
    wire N__20153;
    wire N__20150;
    wire N__20147;
    wire N__20144;
    wire N__20141;
    wire N__20138;
    wire N__20135;
    wire N__20132;
    wire N__20129;
    wire N__20126;
    wire N__20123;
    wire N__20122;
    wire N__20119;
    wire N__20114;
    wire N__20111;
    wire N__20108;
    wire N__20107;
    wire N__20102;
    wire N__20099;
    wire N__20096;
    wire N__20093;
    wire N__20090;
    wire N__20087;
    wire N__20084;
    wire N__20081;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20066;
    wire N__20063;
    wire N__20060;
    wire N__20057;
    wire N__20056;
    wire N__20055;
    wire N__20052;
    wire N__20049;
    wire N__20046;
    wire N__20043;
    wire N__20040;
    wire N__20033;
    wire N__20030;
    wire N__20027;
    wire N__20024;
    wire N__20021;
    wire N__20018;
    wire N__20015;
    wire N__20012;
    wire N__20009;
    wire N__20008;
    wire N__20005;
    wire N__20002;
    wire N__20001;
    wire N__20000;
    wire N__19999;
    wire N__19998;
    wire N__19997;
    wire N__19992;
    wire N__19987;
    wire N__19984;
    wire N__19983;
    wire N__19982;
    wire N__19981;
    wire N__19980;
    wire N__19979;
    wire N__19978;
    wire N__19977;
    wire N__19976;
    wire N__19973;
    wire N__19970;
    wire N__19969;
    wire N__19968;
    wire N__19967;
    wire N__19966;
    wire N__19965;
    wire N__19964;
    wire N__19963;
    wire N__19962;
    wire N__19961;
    wire N__19960;
    wire N__19959;
    wire N__19958;
    wire N__19953;
    wire N__19950;
    wire N__19947;
    wire N__19940;
    wire N__19931;
    wire N__19928;
    wire N__19927;
    wire N__19926;
    wire N__19925;
    wire N__19922;
    wire N__19907;
    wire N__19896;
    wire N__19895;
    wire N__19892;
    wire N__19887;
    wire N__19882;
    wire N__19879;
    wire N__19872;
    wire N__19865;
    wire N__19862;
    wire N__19847;
    wire N__19844;
    wire N__19841;
    wire N__19838;
    wire N__19835;
    wire N__19832;
    wire N__19831;
    wire N__19830;
    wire N__19829;
    wire N__19828;
    wire N__19825;
    wire N__19824;
    wire N__19823;
    wire N__19822;
    wire N__19821;
    wire N__19820;
    wire N__19819;
    wire N__19818;
    wire N__19817;
    wire N__19816;
    wire N__19815;
    wire N__19814;
    wire N__19811;
    wire N__19808;
    wire N__19807;
    wire N__19806;
    wire N__19805;
    wire N__19804;
    wire N__19803;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19789;
    wire N__19788;
    wire N__19785;
    wire N__19782;
    wire N__19779;
    wire N__19778;
    wire N__19777;
    wire N__19776;
    wire N__19773;
    wire N__19770;
    wire N__19767;
    wire N__19764;
    wire N__19761;
    wire N__19758;
    wire N__19755;
    wire N__19752;
    wire N__19749;
    wire N__19748;
    wire N__19747;
    wire N__19744;
    wire N__19741;
    wire N__19740;
    wire N__19739;
    wire N__19738;
    wire N__19735;
    wire N__19732;
    wire N__19729;
    wire N__19726;
    wire N__19721;
    wire N__19712;
    wire N__19697;
    wire N__19694;
    wire N__19687;
    wire N__19684;
    wire N__19677;
    wire N__19674;
    wire N__19663;
    wire N__19658;
    wire N__19649;
    wire N__19646;
    wire N__19635;
    wire N__19632;
    wire N__19629;
    wire N__19626;
    wire N__19623;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19598;
    wire N__19595;
    wire N__19592;
    wire N__19589;
    wire N__19586;
    wire N__19583;
    wire N__19580;
    wire N__19577;
    wire N__19574;
    wire N__19571;
    wire N__19568;
    wire N__19565;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19553;
    wire N__19550;
    wire N__19547;
    wire N__19544;
    wire N__19541;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19520;
    wire N__19517;
    wire N__19514;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19502;
    wire N__19499;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19484;
    wire N__19481;
    wire N__19478;
    wire N__19475;
    wire N__19472;
    wire N__19469;
    wire N__19466;
    wire N__19463;
    wire N__19460;
    wire N__19457;
    wire N__19454;
    wire N__19451;
    wire N__19448;
    wire N__19445;
    wire N__19442;
    wire N__19439;
    wire N__19436;
    wire N__19433;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19412;
    wire N__19409;
    wire N__19406;
    wire N__19403;
    wire N__19400;
    wire N__19397;
    wire N__19394;
    wire N__19391;
    wire N__19388;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19349;
    wire N__19346;
    wire N__19343;
    wire N__19340;
    wire N__19337;
    wire N__19334;
    wire N__19331;
    wire N__19328;
    wire N__19325;
    wire N__19322;
    wire N__19319;
    wire N__19316;
    wire N__19313;
    wire N__19310;
    wire N__19307;
    wire N__19304;
    wire N__19301;
    wire N__19298;
    wire N__19295;
    wire N__19292;
    wire N__19289;
    wire N__19286;
    wire N__19283;
    wire N__19280;
    wire N__19277;
    wire N__19274;
    wire N__19271;
    wire N__19268;
    wire N__19265;
    wire N__19262;
    wire N__19259;
    wire N__19256;
    wire N__19253;
    wire N__19250;
    wire N__19247;
    wire N__19244;
    wire N__19241;
    wire N__19238;
    wire N__19235;
    wire N__19232;
    wire N__19229;
    wire N__19226;
    wire N__19223;
    wire N__19220;
    wire N__19217;
    wire N__19214;
    wire N__19211;
    wire N__19208;
    wire N__19205;
    wire N__19202;
    wire N__19199;
    wire N__19196;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire N__19178;
    wire N__19175;
    wire N__19172;
    wire N__19169;
    wire N__19166;
    wire N__19163;
    wire N__19160;
    wire N__19157;
    wire N__19154;
    wire N__19151;
    wire N__19148;
    wire N__19145;
    wire N__19142;
    wire N__19139;
    wire N__19136;
    wire N__19133;
    wire N__19130;
    wire N__19127;
    wire N__19124;
    wire N__19121;
    wire N__19118;
    wire N__19115;
    wire N__19112;
    wire N__19109;
    wire N__19106;
    wire N__19103;
    wire N__19100;
    wire N__19097;
    wire N__19094;
    wire N__19091;
    wire N__19088;
    wire N__19085;
    wire N__19082;
    wire N__19079;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19058;
    wire N__19055;
    wire N__19052;
    wire N__19049;
    wire N__19046;
    wire N__19043;
    wire N__19040;
    wire N__19037;
    wire N__19034;
    wire N__19031;
    wire N__19028;
    wire N__19025;
    wire N__19022;
    wire N__19019;
    wire N__19016;
    wire N__19013;
    wire N__19010;
    wire N__19007;
    wire N__19004;
    wire N__19001;
    wire N__18998;
    wire N__18995;
    wire N__18992;
    wire N__18989;
    wire N__18986;
    wire N__18983;
    wire N__18980;
    wire N__18977;
    wire N__18974;
    wire N__18971;
    wire N__18968;
    wire N__18965;
    wire N__18962;
    wire N__18959;
    wire N__18956;
    wire N__18953;
    wire N__18950;
    wire N__18947;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18935;
    wire N__18932;
    wire N__18929;
    wire N__18926;
    wire N__18923;
    wire N__18920;
    wire N__18917;
    wire N__18914;
    wire N__18911;
    wire N__18908;
    wire N__18905;
    wire N__18902;
    wire N__18899;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18866;
    wire N__18863;
    wire N__18860;
    wire N__18857;
    wire N__18854;
    wire N__18851;
    wire N__18848;
    wire N__18845;
    wire N__18842;
    wire N__18839;
    wire N__18836;
    wire N__18835;
    wire N__18830;
    wire N__18827;
    wire N__18824;
    wire N__18821;
    wire N__18820;
    wire N__18817;
    wire N__18814;
    wire N__18809;
    wire N__18806;
    wire N__18803;
    wire N__18800;
    wire N__18797;
    wire N__18794;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18779;
    wire N__18776;
    wire N__18773;
    wire N__18770;
    wire N__18767;
    wire N__18764;
    wire N__18761;
    wire N__18758;
    wire N__18755;
    wire N__18752;
    wire N__18749;
    wire N__18746;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18734;
    wire N__18731;
    wire N__18728;
    wire N__18725;
    wire N__18722;
    wire N__18719;
    wire N__18716;
    wire N__18713;
    wire N__18710;
    wire N__18707;
    wire N__18704;
    wire N__18701;
    wire N__18698;
    wire N__18695;
    wire N__18692;
    wire N__18689;
    wire N__18686;
    wire N__18683;
    wire N__18680;
    wire N__18677;
    wire N__18674;
    wire N__18671;
    wire N__18668;
    wire N__18665;
    wire N__18664;
    wire N__18663;
    wire N__18662;
    wire N__18661;
    wire N__18660;
    wire N__18659;
    wire N__18658;
    wire N__18657;
    wire N__18656;
    wire N__18655;
    wire N__18654;
    wire N__18651;
    wire N__18648;
    wire N__18645;
    wire N__18642;
    wire N__18639;
    wire N__18636;
    wire N__18633;
    wire N__18630;
    wire N__18627;
    wire N__18624;
    wire N__18621;
    wire N__18618;
    wire N__18615;
    wire N__18608;
    wire N__18599;
    wire N__18594;
    wire N__18589;
    wire N__18578;
    wire N__18575;
    wire N__18572;
    wire N__18569;
    wire N__18566;
    wire N__18563;
    wire N__18560;
    wire N__18557;
    wire N__18554;
    wire N__18551;
    wire N__18548;
    wire N__18545;
    wire N__18542;
    wire N__18539;
    wire N__18536;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18482;
    wire N__18479;
    wire N__18476;
    wire N__18473;
    wire N__18470;
    wire N__18467;
    wire N__18464;
    wire N__18461;
    wire N__18458;
    wire N__18455;
    wire N__18452;
    wire N__18449;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18431;
    wire N__18428;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18395;
    wire N__18392;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18380;
    wire N__18377;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18365;
    wire N__18362;
    wire N__18359;
    wire N__18356;
    wire N__18353;
    wire N__18350;
    wire N__18347;
    wire N__18344;
    wire N__18341;
    wire N__18338;
    wire N__18335;
    wire N__18332;
    wire N__18329;
    wire N__18326;
    wire N__18323;
    wire delay_tr_input_ibuf_gb_io_gb_input;
    wire delay_hc_input_ibuf_gb_io_gb_input;
    wire GNDG0;
    wire VCCG0;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_0 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_15 ;
    wire bfn_1_11_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_8 ;
    wire bfn_1_12_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ;
    wire rgb_drv_RNOZ0;
    wire delay_hc_input_c_g;
    wire \current_shift_inst.PI_CTRL.un1_integrator ;
    wire bfn_3_13_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_2 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_3 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_5 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_6 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_8 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire bfn_3_14_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_10 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_11 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_12 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_13 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_14 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_16 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_17 ;
    wire bfn_3_15_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_18 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_19 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_21 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_22 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_24 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_25 ;
    wire bfn_3_16_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_26 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_28 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_29 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_30 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire N_38_i_i;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_44_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_2 ;
    wire \current_shift_inst.PI_CTRL.N_77_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_43 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.N_46 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.N_47 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire elapsed_time_ns_1_RNIUVBN9_0_11;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axb_0 ;
    wire bfn_7_13_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_7 ;
    wire bfn_7_14_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_13 ;
    wire bfn_7_20_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire bfn_7_21_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire bfn_7_22_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire bfn_7_23_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_12 ;
    wire il_max_comp1_c;
    wire bfn_8_7_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire bfn_8_8_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire bfn_8_9_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire bfn_8_10_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire bfn_8_11_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ;
    wire bfn_8_12_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_8_13_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire bfn_8_14_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ;
    wire \current_shift_inst.elapsed_time_ns_s1_fast_31 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire bfn_8_19_0_;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire bfn_8_20_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire bfn_8_21_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire bfn_8_22_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire s4_phy_c;
    wire GB_BUFFER_clock_output_0_THRU_CO;
    wire il_min_comp1_c;
    wire elapsed_time_ns_1_RNI24CN9_0_15;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ;
    wire elapsed_time_ns_1_RNIK63T9_0_8_cascade_;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_1 ;
    wire bfn_9_11_0_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_9 ;
    wire bfn_9_12_0_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt18 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ;
    wire bfn_9_13_0_;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_30 ;
    wire \current_shift_inst.control_input_18 ;
    wire bfn_9_14_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ;
    wire \current_shift_inst.control_input_cry_0 ;
    wire \current_shift_inst.control_input_axb_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ;
    wire \current_shift_inst.control_input_cry_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ;
    wire \current_shift_inst.control_input_cry_2 ;
    wire \current_shift_inst.control_input_axb_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ;
    wire \current_shift_inst.control_input_cry_3 ;
    wire \current_shift_inst.control_input_axb_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ;
    wire \current_shift_inst.control_input_cry_4 ;
    wire \current_shift_inst.control_input_axb_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ;
    wire \current_shift_inst.control_input_cry_5 ;
    wire \current_shift_inst.control_input_axb_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ;
    wire \current_shift_inst.control_input_cry_6 ;
    wire \current_shift_inst.control_input_cry_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ;
    wire bfn_9_15_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ;
    wire \current_shift_inst.control_input_cry_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ;
    wire \current_shift_inst.control_input_cry_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ;
    wire \current_shift_inst.control_input_cry_10 ;
    wire \current_shift_inst.control_input_axb_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ;
    wire \current_shift_inst.control_input_cry_11 ;
    wire \current_shift_inst.control_input_cry_12 ;
    wire \current_shift_inst.control_input_31 ;
    wire \current_shift_inst.control_input_axb_1 ;
    wire \current_shift_inst.control_input_axb_3 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ;
    wire bfn_9_16_0_;
    wire \current_shift_inst.un10_control_input_cry_0 ;
    wire \current_shift_inst.un10_control_input_cry_1 ;
    wire \current_shift_inst.un10_control_input_cry_2 ;
    wire \current_shift_inst.un10_control_input_cry_3 ;
    wire \current_shift_inst.un10_control_input_cry_4 ;
    wire \current_shift_inst.un10_control_input_cry_5 ;
    wire \current_shift_inst.un10_control_input_cry_6 ;
    wire \current_shift_inst.un10_control_input_cry_7 ;
    wire \current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ;
    wire bfn_9_17_0_;
    wire \current_shift_inst.un10_control_input_cry_8 ;
    wire \current_shift_inst.un10_control_input_cry_9 ;
    wire \current_shift_inst.un10_control_input_cry_10 ;
    wire \current_shift_inst.un10_control_input_cry_11 ;
    wire \current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_12 ;
    wire \current_shift_inst.un10_control_input_cry_13 ;
    wire \current_shift_inst.un10_control_input_cry_14 ;
    wire \current_shift_inst.un10_control_input_cry_15 ;
    wire bfn_9_18_0_;
    wire \current_shift_inst.un10_control_input_cry_16 ;
    wire \current_shift_inst.un10_control_input_cry_17 ;
    wire \current_shift_inst.un10_control_input_cry_18 ;
    wire \current_shift_inst.un10_control_input_cry_19 ;
    wire \current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_20 ;
    wire \current_shift_inst.un10_control_input_cry_21 ;
    wire \current_shift_inst.un10_control_input_cry_22 ;
    wire \current_shift_inst.un10_control_input_cry_23 ;
    wire bfn_9_19_0_;
    wire \current_shift_inst.un10_control_input_cry_24 ;
    wire \current_shift_inst.un10_control_input_cry_25 ;
    wire \current_shift_inst.un10_control_input_cry_26 ;
    wire \current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_27 ;
    wire \current_shift_inst.un10_control_input_cry_28 ;
    wire \current_shift_inst.un10_control_input_cry_29 ;
    wire \current_shift_inst.un10_control_input_cry_30 ;
    wire \current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_2 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_11 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_1 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_10 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_13 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ;
    wire elapsed_time_ns_1_RNIH33T9_0_5;
    wire elapsed_time_ns_1_RNIG23T9_0_4;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ;
    wire elapsed_time_ns_1_RNIE03T9_0_2;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ;
    wire elapsed_time_ns_1_RNIF13T9_0_3;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ;
    wire elapsed_time_ns_1_RNI68CN9_0_19;
    wire elapsed_time_ns_1_RNI57CN9_0_18;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ;
    wire elapsed_time_ns_1_RNIK63T9_0_8;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ;
    wire elapsed_time_ns_1_RNITUBN9_0_10;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ;
    wire elapsed_time_ns_1_RNIL73T9_0_9;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ;
    wire elapsed_time_ns_1_RNI7ADN9_0_29;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ;
    wire elapsed_time_ns_1_RNI02CN9_0_13;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ;
    wire elapsed_time_ns_1_RNIV2EN9_0_30;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ;
    wire elapsed_time_ns_1_RNI04EN9_0_31;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ;
    wire elapsed_time_ns_1_RNIDV2T9_0_1;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_df30_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt30 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ;
    wire \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt16 ;
    wire \current_shift_inst.elapsed_time_ns_s1_22 ;
    wire il_min_comp1_D1;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire \current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt26 ;
    wire \current_shift_inst.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ;
    wire \current_shift_inst.control_input_axb_0 ;
    wire \current_shift_inst.control_input_axb_0_cascade_ ;
    wire \current_shift_inst.N_1288_i ;
    wire \current_shift_inst.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_1 ;
    wire \current_shift_inst.un4_control_input1_2 ;
    wire bfn_10_18_0_;
    wire \current_shift_inst.un4_control_input_1_axb_2 ;
    wire \current_shift_inst.un4_control_input_1_cry_1 ;
    wire \current_shift_inst.un4_control_input_1_axb_3 ;
    wire \current_shift_inst.un4_control_input_1_cry_2 ;
    wire \current_shift_inst.un4_control_input_1_axb_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_3 ;
    wire \current_shift_inst.un4_control_input_1_axb_5 ;
    wire \current_shift_inst.un4_control_input1_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_4 ;
    wire \current_shift_inst.un4_control_input_1_axb_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_5 ;
    wire \current_shift_inst.un4_control_input_1_axb_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_6 ;
    wire \current_shift_inst.un4_control_input_1_axb_8 ;
    wire \current_shift_inst.un4_control_input_1_cry_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_8 ;
    wire \current_shift_inst.un4_control_input_1_axb_9 ;
    wire \current_shift_inst.un4_control_input1_10 ;
    wire bfn_10_19_0_;
    wire \current_shift_inst.un4_control_input_1_axb_10 ;
    wire \current_shift_inst.un4_control_input_1_cry_9 ;
    wire \current_shift_inst.un4_control_input_1_cry_10 ;
    wire \current_shift_inst.un4_control_input_1_axb_12 ;
    wire \current_shift_inst.un4_control_input_1_cry_11 ;
    wire \current_shift_inst.un4_control_input_1_axb_13 ;
    wire \current_shift_inst.un4_control_input_1_cry_12 ;
    wire \current_shift_inst.un4_control_input_1_cry_13 ;
    wire \current_shift_inst.un4_control_input_1_axb_15 ;
    wire \current_shift_inst.un4_control_input1_16 ;
    wire \current_shift_inst.un4_control_input_1_cry_14 ;
    wire \current_shift_inst.un4_control_input_1_axb_16 ;
    wire \current_shift_inst.un4_control_input_1_cry_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_16 ;
    wire \current_shift_inst.un4_control_input_1_axb_17 ;
    wire bfn_10_20_0_;
    wire \current_shift_inst.un4_control_input_1_cry_17 ;
    wire \current_shift_inst.un4_control_input_1_axb_19 ;
    wire \current_shift_inst.un4_control_input_1_cry_18 ;
    wire \current_shift_inst.un4_control_input_1_axb_20 ;
    wire \current_shift_inst.un4_control_input_1_cry_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_21 ;
    wire \current_shift_inst.un4_control_input1_22 ;
    wire \current_shift_inst.un4_control_input_1_cry_20 ;
    wire \current_shift_inst.un4_control_input_1_axb_22 ;
    wire \current_shift_inst.un4_control_input_1_cry_21 ;
    wire \current_shift_inst.un4_control_input_1_axb_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_22 ;
    wire \current_shift_inst.un4_control_input_1_axb_24 ;
    wire \current_shift_inst.un4_control_input_1_cry_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_24 ;
    wire \current_shift_inst.un4_control_input_1_axb_25 ;
    wire bfn_10_21_0_;
    wire \current_shift_inst.un4_control_input_1_cry_25 ;
    wire \current_shift_inst.un4_control_input_1_cry_26 ;
    wire \current_shift_inst.un4_control_input_1_axb_28 ;
    wire \current_shift_inst.un4_control_input_1_cry_27 ;
    wire \current_shift_inst.un4_control_input_1_axb_29 ;
    wire \current_shift_inst.un4_control_input_1_cry_28 ;
    wire \current_shift_inst.un4_control_input1_31 ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_ ;
    wire \current_shift_inst.un4_control_input_1_axb_18 ;
    wire \current_shift_inst.un4_control_input_1_axb_27 ;
    wire \current_shift_inst.un4_control_input_1_axb_26 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ;
    wire elapsed_time_ns_1_RNII43T9_0_6;
    wire elapsed_time_ns_1_RNII43T9_0_6_cascade_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ;
    wire elapsed_time_ns_1_RNI46CN9_0_17;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ;
    wire elapsed_time_ns_1_RNIJ53T9_0_7;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_df30_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire bfn_11_7_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire bfn_11_8_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt18 ;
    wire bfn_11_9_0_;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt26 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt28 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ;
    wire bfn_11_11_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ;
    wire bfn_11_12_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ;
    wire bfn_11_13_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ;
    wire bfn_11_14_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ;
    wire bfn_11_15_0_;
    wire \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_0_s1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1 ;
    wire \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ;
    wire bfn_11_16_0_;
    wire \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_8_s1 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1 ;
    wire bfn_11_17_0_;
    wire \current_shift_inst.un38_control_input_cry_16_s1 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ;
    wire \current_shift_inst.un38_control_input_0_s1_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s1 ;
    wire \current_shift_inst.un38_control_input_cry_23_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_24 ;
    wire bfn_11_18_0_;
    wire \current_shift_inst.un38_control_input_0_s1_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_26 ;
    wire \current_shift_inst.un38_control_input_cry_25_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s1 ;
    wire \current_shift_inst.un38_control_input_cry_27_s1 ;
    wire \current_shift_inst.un38_control_input_cry_28_s1 ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ;
    wire \current_shift_inst.un38_control_input_cry_29_s1 ;
    wire \current_shift_inst.un38_control_input_cry_30_s1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.un4_control_input1_9 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ;
    wire \current_shift_inst.un4_control_input_1_axb_11 ;
    wire \current_shift_inst.un4_control_input_1_axb_14 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ;
    wire \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ;
    wire \current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ;
    wire \current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_27 ;
    wire \current_shift_inst.un4_control_input1_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ;
    wire \current_shift_inst.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.un4_control_input1_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_26 ;
    wire \current_shift_inst.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.un4_control_input1_29 ;
    wire \current_shift_inst.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.un4_control_input1_25 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31_rep1 ;
    wire \current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_14 ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_11_23_0_;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_11_24_0_;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire s3_phy_c;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ;
    wire elapsed_time_ns_1_RNI35CN9_0_16;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ;
    wire bfn_12_6_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire bfn_12_7_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire bfn_12_8_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ;
    wire bfn_12_9_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst2.state_RNIG7JFZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.runningZ0 ;
    wire \phase_controller_inst2.start_timer_hcZ0 ;
    wire \phase_controller_inst2.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst2.stoper_hc.un2_start_0_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.start_latchedZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire elapsed_time_ns_1_RNI58DN9_0_27;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt24 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ;
    wire elapsed_time_ns_1_RNIV0CN9_0_12;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ;
    wire elapsed_time_ns_1_RNI36DN9_0_25;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire elapsed_time_ns_1_RNI47DN9_0_26;
    wire \phase_controller_inst2.stoper_hc.un1_start_g ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ;
    wire \current_shift_inst.un38_control_input_5_0 ;
    wire bfn_12_13_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2 ;
    wire \current_shift_inst.un38_control_input_5_1 ;
    wire \current_shift_inst.un38_control_input_cry_0_s0 ;
    wire \current_shift_inst.un38_control_input_cry_1_s0 ;
    wire \current_shift_inst.un38_control_input_cry_2_s0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0 ;
    wire \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ;
    wire bfn_12_14_0_;
    wire \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_8_s0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0 ;
    wire bfn_12_15_0_;
    wire \current_shift_inst.un38_control_input_cry_16_s0 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ;
    wire \current_shift_inst.un38_control_input_0_s0_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s0 ;
    wire \current_shift_inst.un38_control_input_cry_23_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ;
    wire \current_shift_inst.un38_control_input_0_s0_24 ;
    wire bfn_12_16_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ;
    wire \current_shift_inst.un38_control_input_0_s0_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ;
    wire \current_shift_inst.un38_control_input_0_s0_26 ;
    wire \current_shift_inst.un38_control_input_cry_25_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ;
    wire \current_shift_inst.un38_control_input_0_s0_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ;
    wire \current_shift_inst.un38_control_input_cry_27_s0 ;
    wire \current_shift_inst.un38_control_input_cry_28_s0 ;
    wire \current_shift_inst.un38_control_input_cry_29_s0 ;
    wire \current_shift_inst.un38_control_input_axb_31_s0 ;
    wire \current_shift_inst.un38_control_input_0_s1_31 ;
    wire \current_shift_inst.un38_control_input_cry_30_s0 ;
    wire \current_shift_inst.control_input_axb_11 ;
    wire \current_shift_inst.un38_control_input_0_s1_28 ;
    wire \current_shift_inst.un38_control_input_0_s0_28 ;
    wire \current_shift_inst.control_input_axb_8 ;
    wire \current_shift_inst.un38_control_input_0_s1_29 ;
    wire \current_shift_inst.un38_control_input_0_s0_29 ;
    wire \current_shift_inst.control_input_axb_9 ;
    wire \current_shift_inst.un38_control_input_0_s1_30 ;
    wire \current_shift_inst.un38_control_input_0_s0_30 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ;
    wire \current_shift_inst.control_input_axb_10 ;
    wire \delay_measurement_inst.delay_hc_timer.N_199_i ;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.N_198_i ;
    wire \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.un4_control_input1_4 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ;
    wire \current_shift_inst.un4_control_input1_8 ;
    wire \current_shift_inst.elapsed_time_ns_s1_8 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.un4_control_input1_7 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.un4_control_input1_17 ;
    wire \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.un4_control_input1_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ;
    wire \current_shift_inst.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.un4_control_input1_12 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_11 ;
    wire \current_shift_inst.un4_control_input1_11 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_23 ;
    wire \current_shift_inst.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ;
    wire \current_shift_inst.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.un4_control_input1_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.un4_control_input1_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ;
    wire \current_shift_inst.un4_control_input1_24 ;
    wire \current_shift_inst.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ;
    wire \current_shift_inst.elapsed_time_ns_s1_19 ;
    wire \current_shift_inst.un4_control_input1_19 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ;
    wire bfn_12_21_0_;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire bfn_12_22_0_;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_2_1_16 ;
    wire \pwm_generator_inst.un2_threshold_2_1_15 ;
    wire \pwm_generator_inst.threshold_3 ;
    wire \pwm_generator_inst.threshold_4 ;
    wire \pwm_generator_inst.threshold_5 ;
    wire \pwm_generator_inst.un14_counter_6 ;
    wire \pwm_generator_inst.un14_counter_7 ;
    wire \pwm_generator_inst.un14_counter_1 ;
    wire \pwm_generator_inst.threshold_0 ;
    wire \pwm_generator_inst.threshold_2 ;
    wire \pwm_generator_inst.un14_counter_8 ;
    wire N_19_1;
    wire \pwm_generator_inst.threshold_9 ;
    wire \pll_inst.red_c_i ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ;
    wire elapsed_time_ns_1_RNI13CN9_0_14;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt16 ;
    wire \phase_controller_inst2.tr_time_passed ;
    wire \phase_controller_inst2.stateZ0Z_0 ;
    wire \phase_controller_inst2.state_RNI9M3OZ0Z_0_cascade_ ;
    wire \phase_controller_inst2.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_inst2.stateZ0Z_3 ;
    wire il_max_comp2_c;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt22 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ;
    wire elapsed_time_ns_1_RNI14DN9_0_23;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ;
    wire elapsed_time_ns_1_RNI03DN9_0_22;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt20 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ;
    wire elapsed_time_ns_1_RNIU0DN9_0_20;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ;
    wire elapsed_time_ns_1_RNI69DN9_0_28;
    wire elapsed_time_ns_1_RNI69DN9_0_28_cascade_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ;
    wire il_min_comp2_c;
    wire \phase_controller_inst2.hc_time_passed ;
    wire \phase_controller_inst2.stateZ0Z_2 ;
    wire \phase_controller_inst2.stateZ0Z_1 ;
    wire \phase_controller_inst2.state_RNI9M3OZ0Z_0 ;
    wire \phase_controller_inst2.start_timer_tr_RNO_0_0_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.runningZ0 ;
    wire \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_df30 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ;
    wire elapsed_time_ns_1_RNI0AOBB_0_13_cascade_;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31 ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_18 ;
    wire \current_shift_inst.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.un4_control_input1_5 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.un4_control_input1_13 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.un4_control_input1_15 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.un4_control_input1_14 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ;
    wire il_max_comp1_D1;
    wire \current_shift_inst.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.un4_control_input1_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire \current_shift_inst.timer_s1.N_162_i_g ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1 ;
    wire \current_shift_inst.un4_control_input1_1 ;
    wire \current_shift_inst.un4_control_input1_1_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_s1_1 ;
    wire \current_shift_inst.un38_control_input_cry_0_s0_sf ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.un38_control_input_5_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_3 ;
    wire \current_shift_inst.un4_control_input1_3 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ;
    wire \current_shift_inst.timer_s1.N_162_i ;
    wire \current_shift_inst.timer_s1.N_163_i ;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.un1_counterlto2_0_cascade_ ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \current_shift_inst.timer_s1.running_i ;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.un1_counterlto9_2_cascade_ ;
    wire \pwm_generator_inst.un1_counterlt9 ;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_6 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_8 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ;
    wire bfn_13_24_0_;
    wire \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_0 ;
    wire \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_1 ;
    wire \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_2 ;
    wire \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_3 ;
    wire \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_4 ;
    wire \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ;
    wire \pwm_generator_inst.un19_threshold_cry_5 ;
    wire \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ;
    wire \pwm_generator_inst.un19_threshold_cry_6 ;
    wire \pwm_generator_inst.un19_threshold_cry_7 ;
    wire \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ;
    wire bfn_13_25_0_;
    wire \pwm_generator_inst.un19_threshold_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433 ;
    wire \pwm_generator_inst.un19_threshold_axb_5 ;
    wire \pwm_generator_inst.un19_threshold_axb_3 ;
    wire \pwm_generator_inst.un19_threshold_axb_6 ;
    wire \pwm_generator_inst.un19_threshold_axb_4 ;
    wire \pwm_generator_inst.un19_threshold_axb_0 ;
    wire \pwm_generator_inst.un19_threshold_axb_8 ;
    wire \pwm_generator_inst.un19_threshold_axb_2 ;
    wire \pwm_generator_inst.un19_threshold_axb_7 ;
    wire \pwm_generator_inst.un2_threshold_2_0 ;
    wire \pwm_generator_inst.un2_threshold_1_15 ;
    wire bfn_13_28_0_;
    wire \pwm_generator_inst.un2_threshold_2_1 ;
    wire \pwm_generator_inst.un2_threshold_1_16 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_2_2 ;
    wire \pwm_generator_inst.un2_threshold_1_17 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_2_3 ;
    wire \pwm_generator_inst.un2_threshold_1_18 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_2_4 ;
    wire \pwm_generator_inst.un2_threshold_1_19 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_2_5 ;
    wire \pwm_generator_inst.un2_threshold_1_20 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_2_6 ;
    wire \pwm_generator_inst.un2_threshold_1_21 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_2_7 ;
    wire \pwm_generator_inst.un2_threshold_1_22 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_2_8 ;
    wire \pwm_generator_inst.un2_threshold_1_23 ;
    wire bfn_13_29_0_;
    wire \pwm_generator_inst.un2_threshold_2_9 ;
    wire \pwm_generator_inst.un2_threshold_1_24 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_2_10 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_2_11 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_2_12 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_2_13 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_2_14 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_1_25 ;
    wire \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_14 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15 ;
    wire \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ;
    wire bfn_13_30_0_;
    wire \phase_controller_inst2.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst2.start_timer_trZ0 ;
    wire \phase_controller_inst2.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst1.stoper_hc.runningZ0 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_1 ;
    wire bfn_14_7_0_;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_9 ;
    wire bfn_14_8_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt16 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_16 ;
    wire bfn_14_9_0_;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ;
    wire bfn_14_10_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ;
    wire bfn_14_11_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ;
    wire bfn_14_12_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ;
    wire bfn_14_13_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ;
    wire bfn_14_14_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire bfn_14_15_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire bfn_14_16_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire bfn_14_17_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_3 ;
    wire state_ns_i_a3_1;
    wire il_max_comp1_D2;
    wire \current_shift_inst.PI_CTRL.prop_term_1_5 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_4 ;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_9 ;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_0 ;
    wire bfn_14_25_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_2 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_7 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_8 ;
    wire bfn_14_26_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_9 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ;
    wire \pwm_generator_inst.un19_threshold_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_10 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_11 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_12 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_13 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_14 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_15 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_16 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ;
    wire bfn_14_27_0_;
    wire \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_16 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_17 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_axb_18 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_17 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_15 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_12 ;
    wire \pwm_generator_inst.un3_threshold ;
    wire bfn_14_28_0_;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_0 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_1 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_2 ;
    wire \pwm_generator_inst.un3_threshold_axbZ0Z_4 ;
    wire \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ;
    wire \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ;
    wire \pwm_generator_inst.un3_threshold_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ;
    wire \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ;
    wire \pwm_generator_inst.un3_threshold_cry_5 ;
    wire CONSTANT_ONE_NET;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ;
    wire \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ;
    wire \pwm_generator_inst.un3_threshold_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ;
    wire \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ;
    wire bfn_14_29_0_;
    wire \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_8 ;
    wire \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_9 ;
    wire \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_10 ;
    wire \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_11 ;
    wire \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_15 ;
    wire \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ;
    wire bfn_14_30_0_;
    wire \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_16 ;
    wire \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_17 ;
    wire \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_cry_19 ;
    wire \pwm_generator_inst.un3_threshold_cry_19_THRU_CO ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire elapsed_time_ns_1_RNI25DN9_0_24;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt18 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt24 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt20 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt22 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ;
    wire elapsed_time_ns_1_RNIV8OBB_0_12_cascade_;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ;
    wire elapsed_time_ns_1_RNI0AOBB_0_13;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire bfn_15_14_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire bfn_15_15_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire bfn_15_16_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire bfn_15_17_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire \phase_controller_inst1.start_timer_hc_0_sqmuxa ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_7 ;
    wire s1_phy_c;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire state_3;
    wire T01_c;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire bfn_15_23_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire bfn_15_24_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire bfn_15_25_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire bfn_15_26_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_14 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt26 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3 ;
    wire elapsed_time_ns_1_RNIV1DN9_0_21;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ;
    wire elapsed_time_ns_1_RNIT6OBB_0_10;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ;
    wire elapsed_time_ns_1_RNIT6OBB_0_10_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ;
    wire elapsed_time_ns_1_RNIV8OBB_0_12;
    wire \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ;
    wire elapsed_time_ns_1_RNI3DOBB_0_16;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ;
    wire elapsed_time_ns_1_RNI4EOBB_0_17;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ;
    wire elapsed_time_ns_1_RNIV9PBB_0_21;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ;
    wire elapsed_time_ns_1_RNI7IPBB_0_29;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire \phase_controller_inst1.stoper_hc.start_latchedZ0 ;
    wire delay_tr_input_c_g;
    wire \phase_controller_inst1.hc_time_passed ;
    wire \phase_controller_inst1.start_timer_tr_RNOZ0Z_0 ;
    wire \phase_controller_inst1.state_RNIE87FZ0Z_2 ;
    wire T45_c;
    wire il_min_comp1_D2;
    wire T23_c;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire s2_phy_c;
    wire start_stop_c;
    wire phase_controller_inst1_state_4;
    wire \phase_controller_inst1.stoper_tr.runningZ0 ;
    wire elapsed_time_ns_1_RNI2COBB_0_15;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ;
    wire elapsed_time_ns_1_RNI5FOBB_0_18;
    wire elapsed_time_ns_1_RNI5FOBB_0_18_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ;
    wire elapsed_time_ns_1_RNIU8PBB_0_20;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ;
    wire elapsed_time_ns_1_RNIDC91B_0_1;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ;
    wire elapsed_time_ns_1_RNIED91B_0_2;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ;
    wire elapsed_time_ns_1_RNIFE91B_0_3;
    wire elapsed_time_ns_1_RNIGF91B_0_4;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ;
    wire bfn_17_11_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire bfn_17_12_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire bfn_17_13_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ;
    wire bfn_17_14_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire elapsed_time_ns_1_RNI5GPBB_0_27;
    wire elapsed_time_ns_1_RNI6HPBB_0_28;
    wire elapsed_time_ns_1_RNI6HPBB_0_28_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ;
    wire \delay_measurement_inst.delay_tr_timer.N_200_i ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.N_201_i ;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire T12_c;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire \phase_controller_inst1.state_RNI7NN7Z0Z_0 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_10 ;
    wire elapsed_time_ns_1_RNILK91B_0_9;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ;
    wire elapsed_time_ns_1_RNIIH91B_0_6;
    wire elapsed_time_ns_1_RNI3EPBB_0_25;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ;
    wire elapsed_time_ns_1_RNIHG91B_0_5;
    wire elapsed_time_ns_1_RNIKJ91B_0_8;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ;
    wire elapsed_time_ns_1_RNIJI91B_0_7;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ;
    wire elapsed_time_ns_1_RNI6GOBB_0_19;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_18_10_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_18_11_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt16 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt18 ;
    wire bfn_18_12_0_;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_30 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt24 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ;
    wire elapsed_time_ns_1_RNI2DPBB_0_24;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt30 ;
    wire elapsed_time_ns_1_RNIVAQBB_0_30;
    wire elapsed_time_ns_1_RNIVAQBB_0_30_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_df30 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ;
    wire elapsed_time_ns_1_RNI0CQBB_0_31;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ;
    wire elapsed_time_ns_1_RNI1BOBB_0_14;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst1.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst1.tr_time_passed ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.un1_start_g ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire elapsed_time_ns_1_RNI4FPBB_0_26;
    wire elapsed_time_ns_1_RNIU7OBB_0_11;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt22 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ;
    wire elapsed_time_ns_1_RNI1CPBB_0_23;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_0 ;
    wire elapsed_time_ns_1_RNI0BPBB_0_22;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ;
    wire \pwm_generator_inst.N_16 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4 ;
    wire \current_shift_inst.PI_CTRL.N_27_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0 ;
    wire \current_shift_inst.PI_CTRL.N_98 ;
    wire \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ;
    wire \pwm_generator_inst.N_17 ;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ;
    wire \pwm_generator_inst.un1_duty_inputlt3 ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire pwm_duty_input_7;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire pwm_duty_input_8;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire pwm_duty_input_0;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire pwm_duty_input_3;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire pwm_duty_input_1;
    wire \current_shift_inst.PI_CTRL.N_97 ;
    wire \current_shift_inst.PI_CTRL.N_96 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_3 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire pwm_duty_input_2;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire pwm_duty_input_6;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire pwm_duty_input_5;
    wire \current_shift_inst.PI_CTRL.N_91 ;
    wire \current_shift_inst.PI_CTRL.N_27 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire pwm_duty_input_4;
    wire \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.N_159 ;
    wire pwm_duty_input_9;
    wire _gnd_net_;
    wire clock_output_0;
    wire red_c_g;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__20075),
            .RESETB(N__30797),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clock_output_0));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .A_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .D_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .C_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .B_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__37884),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__37881),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({N__26826,N__26834,N__26825,N__26832,N__26824,N__26831,N__26823,N__26833,N__26820,N__26827,N__26819,N__26828,N__26822,N__26829,N__26821,N__26830}),
            .C({dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31}),
            .B({dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,N__37883,dangling_wire_45,N__37882}),
            .OHOLDTOP(),
            .O({dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,\current_shift_inst.PI_CTRL.integrator_1_0_2_15 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_14 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_13 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_12 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_11 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_10 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_9 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_8 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_7 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_6 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_5 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_4 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_3 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_2 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_1 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__37791),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__37784),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77}),
            .ADDSUBBOT(),
            .A({dangling_wire_78,N__30965,N__30958,N__30963,N__30957,N__30964,N__30956,N__30966,N__30953,N__30959,N__30952,N__30960,N__30954,N__30961,N__30955,N__30962}),
            .C({dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94}),
            .B({dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,N__37790,N__37787,dangling_wire_102,dangling_wire_103,dangling_wire_104,N__37785,N__37789,N__37786,N__37788}),
            .OHOLDTOP(),
            .O({dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,\pwm_generator_inst.un2_threshold_2_1_16 ,\pwm_generator_inst.un2_threshold_2_1_15 ,\pwm_generator_inst.un2_threshold_2_14 ,\pwm_generator_inst.un2_threshold_2_13 ,\pwm_generator_inst.un2_threshold_2_12 ,\pwm_generator_inst.un2_threshold_2_11 ,\pwm_generator_inst.un2_threshold_2_10 ,\pwm_generator_inst.un2_threshold_2_9 ,\pwm_generator_inst.un2_threshold_2_8 ,\pwm_generator_inst.un2_threshold_2_7 ,\pwm_generator_inst.un2_threshold_2_6 ,\pwm_generator_inst.un2_threshold_2_5 ,\pwm_generator_inst.un2_threshold_2_4 ,\pwm_generator_inst.un2_threshold_2_3 ,\pwm_generator_inst.un2_threshold_2_2 ,\pwm_generator_inst.un2_threshold_2_1 ,\pwm_generator_inst.un2_threshold_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__37909),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__37885),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135}),
            .ADDSUBBOT(),
            .A({dangling_wire_136,N__30967,N__30970,N__30968,N__30971,N__30969,N__48825,N__47666,N__47726,N__49207,N__49158,N__49083,N__47571,N__49256,N__49346,N__47636}),
            .C({dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152}),
            .B({dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,N__37891,N__37888,dangling_wire_160,dangling_wire_161,dangling_wire_162,N__37886,N__37890,N__37887,N__37889}),
            .OHOLDTOP(),
            .O({dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167,dangling_wire_168,\pwm_generator_inst.un2_threshold_1_25 ,\pwm_generator_inst.un2_threshold_1_24 ,\pwm_generator_inst.un2_threshold_1_23 ,\pwm_generator_inst.un2_threshold_1_22 ,\pwm_generator_inst.un2_threshold_1_21 ,\pwm_generator_inst.un2_threshold_1_20 ,\pwm_generator_inst.un2_threshold_1_19 ,\pwm_generator_inst.un2_threshold_1_18 ,\pwm_generator_inst.un2_threshold_1_17 ,\pwm_generator_inst.un2_threshold_1_16 ,\pwm_generator_inst.un2_threshold_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.un3_threshold ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .A_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .D_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .C_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .B_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__37798),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__37795),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184}),
            .ADDSUBBOT(),
            .A({dangling_wire_185,N__26780,N__22846,N__20309,N__22921,N__22867,N__36830,N__33898,N__39389,N__33931,N__36931,N__36901,N__36316,N__22804,N__22900,N__47269}),
            .C({dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201}),
            .B({dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,N__37797,dangling_wire_215,N__37796}),
            .OHOLDTOP(),
            .O({dangling_wire_216,dangling_wire_217,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_18 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_17 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_16 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_15 ,\current_shift_inst.PI_CTRL.integrator_1_15 ,\current_shift_inst.PI_CTRL.integrator_1_14 ,\current_shift_inst.PI_CTRL.integrator_1_13 ,\current_shift_inst.PI_CTRL.integrator_1_12 ,\current_shift_inst.PI_CTRL.integrator_1_11 ,\current_shift_inst.PI_CTRL.integrator_1_10 ,\current_shift_inst.PI_CTRL.integrator_1_9 ,\current_shift_inst.PI_CTRL.integrator_1_8 ,\current_shift_inst.PI_CTRL.integrator_1_7 ,\current_shift_inst.PI_CTRL.integrator_1_6 ,\current_shift_inst.PI_CTRL.integrator_1_5 ,\current_shift_inst.PI_CTRL.integrator_1_4 ,\current_shift_inst.PI_CTRL.integrator_1_3 ,\current_shift_inst.PI_CTRL.integrator_1_2 ,\current_shift_inst.PI_CTRL.un1_integrator }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__49533),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__49535),
            .DIN(N__49534),
            .DOUT(N__49533),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__49535),
            .PADOUT(N__49534),
            .PADIN(N__49533),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clock_output_obuf_iopad (
            .OE(N__49524),
            .DIN(N__49523),
            .DOUT(N__49522),
            .PACKAGEPIN(clock_output));
    defparam clock_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam clock_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO clock_output_obuf_preio (
            .PADOEN(N__49524),
            .PADOUT(N__49523),
            .PADIN(N__49522),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21884),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T01_obuf_iopad (
            .OE(N__49515),
            .DIN(N__49514),
            .DOUT(N__49513),
            .PACKAGEPIN(T01));
    defparam T01_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T01_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T01_obuf_preio (
            .PADOEN(N__49515),
            .PADOUT(N__49514),
            .PADIN(N__49513),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__39272),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__49506),
            .DIN(N__49505),
            .DOUT(N__49504),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__49506),
            .PADOUT(N__49505),
            .PADIN(N__49504),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__49497),
            .DIN(N__49496),
            .DOUT(N__49495),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__49497),
            .PADOUT(N__49496),
            .PADIN(N__49495),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T23_obuf_iopad (
            .OE(N__49488),
            .DIN(N__49487),
            .DOUT(N__49486),
            .PACKAGEPIN(T23));
    defparam T23_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T23_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T23_obuf_preio (
            .PADOEN(N__49488),
            .PADOUT(N__49487),
            .PADIN(N__49486),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__42593),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__49479),
            .DIN(N__49478),
            .DOUT(N__49477),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__49479),
            .PADOUT(N__49478),
            .PADIN(N__49477),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__27389),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__49470),
            .DIN(N__49469),
            .DOUT(N__49468),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__49470),
            .PADOUT(N__49469),
            .PADIN(N__49468),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__49461),
            .DIN(N__49460),
            .DOUT(N__49459),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__49461),
            .PADOUT(N__49460),
            .PADIN(N__49459),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__43037),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T12_obuf_iopad (
            .OE(N__49452),
            .DIN(N__49451),
            .DOUT(N__49450),
            .PACKAGEPIN(T12));
    defparam T12_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T12_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T12_obuf_preio (
            .PADOEN(N__49452),
            .PADOUT(N__49451),
            .PADIN(N__49450),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__44603),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__49443),
            .DIN(N__49442),
            .DOUT(N__49441),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__49443),
            .PADOUT(N__49442),
            .PADIN(N__49441),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__49434),
            .DIN(N__49433),
            .DOUT(N__49432),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__49434),
            .PADOUT(N__49433),
            .PADIN(N__49432),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__39362),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__49425),
            .DIN(N__49424),
            .DOUT(N__49423),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__49425),
            .PADOUT(N__49424),
            .PADIN(N__49423),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21893),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__49416),
            .DIN(N__49415),
            .DOUT(N__49414),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__49416),
            .PADOUT(N__49415),
            .PADIN(N__49414),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__49407),
            .DIN(N__49406),
            .DOUT(N__49405),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__49407),
            .PADOUT(N__49406),
            .PADIN(N__49405),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__27365),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T45_obuf_iopad (
            .OE(N__49398),
            .DIN(N__49397),
            .DOUT(N__49396),
            .PACKAGEPIN(T45));
    defparam T45_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T45_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T45_obuf_preio (
            .PADOEN(N__49398),
            .PADOUT(N__49397),
            .PADIN(N__49396),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__42656),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_gb_io_iopad (
            .OE(N__49389),
            .DIN(N__49388),
            .DOUT(N__49387),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_gb_io_preio (
            .PADOEN(N__49389),
            .PADOUT(N__49388),
            .PADIN(N__49387),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_gb_io_iopad (
            .OE(N__49380),
            .DIN(N__49379),
            .DOUT(N__49378),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_gb_io_preio (
            .PADOEN(N__49380),
            .PADOUT(N__49379),
            .PADIN(N__49378),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__11861 (
            .O(N__49361),
            .I(N__49358));
    LocalMux I__11860 (
            .O(N__49358),
            .I(N__49355));
    Span4Mux_h I__11859 (
            .O(N__49355),
            .I(N__49352));
    Span4Mux_h I__11858 (
            .O(N__49352),
            .I(N__49349));
    Odrv4 I__11857 (
            .O(N__49349),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    InMux I__11856 (
            .O(N__49346),
            .I(N__49342));
    InMux I__11855 (
            .O(N__49345),
            .I(N__49339));
    LocalMux I__11854 (
            .O(N__49342),
            .I(N__49336));
    LocalMux I__11853 (
            .O(N__49339),
            .I(pwm_duty_input_1));
    Odrv4 I__11852 (
            .O(N__49336),
            .I(pwm_duty_input_1));
    InMux I__11851 (
            .O(N__49331),
            .I(N__49322));
    InMux I__11850 (
            .O(N__49330),
            .I(N__49322));
    InMux I__11849 (
            .O(N__49329),
            .I(N__49322));
    LocalMux I__11848 (
            .O(N__49322),
            .I(\current_shift_inst.PI_CTRL.N_97 ));
    CascadeMux I__11847 (
            .O(N__49319),
            .I(N__49313));
    InMux I__11846 (
            .O(N__49318),
            .I(N__49304));
    InMux I__11845 (
            .O(N__49317),
            .I(N__49304));
    InMux I__11844 (
            .O(N__49316),
            .I(N__49304));
    InMux I__11843 (
            .O(N__49313),
            .I(N__49304));
    LocalMux I__11842 (
            .O(N__49304),
            .I(N__49301));
    Span4Mux_s3_h I__11841 (
            .O(N__49301),
            .I(N__49297));
    InMux I__11840 (
            .O(N__49300),
            .I(N__49294));
    Odrv4 I__11839 (
            .O(N__49297),
            .I(\current_shift_inst.PI_CTRL.N_96 ));
    LocalMux I__11838 (
            .O(N__49294),
            .I(\current_shift_inst.PI_CTRL.N_96 ));
    CascadeMux I__11837 (
            .O(N__49289),
            .I(N__49285));
    CascadeMux I__11836 (
            .O(N__49288),
            .I(N__49282));
    InMux I__11835 (
            .O(N__49285),
            .I(N__49276));
    InMux I__11834 (
            .O(N__49282),
            .I(N__49276));
    InMux I__11833 (
            .O(N__49281),
            .I(N__49273));
    LocalMux I__11832 (
            .O(N__49276),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_3 ));
    LocalMux I__11831 (
            .O(N__49273),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_3 ));
    InMux I__11830 (
            .O(N__49268),
            .I(N__49265));
    LocalMux I__11829 (
            .O(N__49265),
            .I(N__49262));
    Span12Mux_s3_h I__11828 (
            .O(N__49262),
            .I(N__49259));
    Odrv12 I__11827 (
            .O(N__49259),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__11826 (
            .O(N__49256),
            .I(N__49253));
    LocalMux I__11825 (
            .O(N__49253),
            .I(N__49249));
    InMux I__11824 (
            .O(N__49252),
            .I(N__49246));
    Span4Mux_s1_h I__11823 (
            .O(N__49249),
            .I(N__49243));
    LocalMux I__11822 (
            .O(N__49246),
            .I(pwm_duty_input_2));
    Odrv4 I__11821 (
            .O(N__49243),
            .I(pwm_duty_input_2));
    CascadeMux I__11820 (
            .O(N__49238),
            .I(N__49235));
    InMux I__11819 (
            .O(N__49235),
            .I(N__49230));
    InMux I__11818 (
            .O(N__49234),
            .I(N__49225));
    InMux I__11817 (
            .O(N__49233),
            .I(N__49225));
    LocalMux I__11816 (
            .O(N__49230),
            .I(N__49222));
    LocalMux I__11815 (
            .O(N__49225),
            .I(N__49219));
    Span4Mux_s2_h I__11814 (
            .O(N__49222),
            .I(N__49214));
    Span4Mux_v I__11813 (
            .O(N__49219),
            .I(N__49214));
    Span4Mux_h I__11812 (
            .O(N__49214),
            .I(N__49211));
    Odrv4 I__11811 (
            .O(N__49211),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    CascadeMux I__11810 (
            .O(N__49208),
            .I(N__49204));
    InMux I__11809 (
            .O(N__49207),
            .I(N__49200));
    InMux I__11808 (
            .O(N__49204),
            .I(N__49195));
    InMux I__11807 (
            .O(N__49203),
            .I(N__49195));
    LocalMux I__11806 (
            .O(N__49200),
            .I(N__49192));
    LocalMux I__11805 (
            .O(N__49195),
            .I(pwm_duty_input_6));
    Odrv4 I__11804 (
            .O(N__49192),
            .I(pwm_duty_input_6));
    CascadeMux I__11803 (
            .O(N__49187),
            .I(N__49184));
    InMux I__11802 (
            .O(N__49184),
            .I(N__49181));
    LocalMux I__11801 (
            .O(N__49181),
            .I(N__49178));
    Span4Mux_v I__11800 (
            .O(N__49178),
            .I(N__49173));
    InMux I__11799 (
            .O(N__49177),
            .I(N__49168));
    InMux I__11798 (
            .O(N__49176),
            .I(N__49168));
    Sp12to4 I__11797 (
            .O(N__49173),
            .I(N__49163));
    LocalMux I__11796 (
            .O(N__49168),
            .I(N__49163));
    Odrv12 I__11795 (
            .O(N__49163),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    InMux I__11794 (
            .O(N__49160),
            .I(N__49153));
    InMux I__11793 (
            .O(N__49159),
            .I(N__49153));
    InMux I__11792 (
            .O(N__49158),
            .I(N__49150));
    LocalMux I__11791 (
            .O(N__49153),
            .I(pwm_duty_input_5));
    LocalMux I__11790 (
            .O(N__49150),
            .I(pwm_duty_input_5));
    InMux I__11789 (
            .O(N__49145),
            .I(N__49142));
    LocalMux I__11788 (
            .O(N__49142),
            .I(\current_shift_inst.PI_CTRL.N_91 ));
    InMux I__11787 (
            .O(N__49139),
            .I(N__49136));
    LocalMux I__11786 (
            .O(N__49136),
            .I(N__49133));
    Odrv12 I__11785 (
            .O(N__49133),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    CascadeMux I__11784 (
            .O(N__49130),
            .I(N__49127));
    InMux I__11783 (
            .O(N__49127),
            .I(N__49122));
    InMux I__11782 (
            .O(N__49126),
            .I(N__49117));
    InMux I__11781 (
            .O(N__49125),
            .I(N__49117));
    LocalMux I__11780 (
            .O(N__49122),
            .I(N__49111));
    LocalMux I__11779 (
            .O(N__49117),
            .I(N__49111));
    InMux I__11778 (
            .O(N__49116),
            .I(N__49108));
    Span4Mux_s2_h I__11777 (
            .O(N__49111),
            .I(N__49103));
    LocalMux I__11776 (
            .O(N__49108),
            .I(N__49103));
    Span4Mux_h I__11775 (
            .O(N__49103),
            .I(N__49100));
    Span4Mux_h I__11774 (
            .O(N__49100),
            .I(N__49097));
    Odrv4 I__11773 (
            .O(N__49097),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    CascadeMux I__11772 (
            .O(N__49094),
            .I(N__49091));
    InMux I__11771 (
            .O(N__49091),
            .I(N__49088));
    LocalMux I__11770 (
            .O(N__49088),
            .I(N__49084));
    InMux I__11769 (
            .O(N__49087),
            .I(N__49080));
    Span4Mux_h I__11768 (
            .O(N__49084),
            .I(N__49077));
    InMux I__11767 (
            .O(N__49083),
            .I(N__49074));
    LocalMux I__11766 (
            .O(N__49080),
            .I(pwm_duty_input_4));
    Odrv4 I__11765 (
            .O(N__49077),
            .I(pwm_duty_input_4));
    LocalMux I__11764 (
            .O(N__49074),
            .I(pwm_duty_input_4));
    CascadeMux I__11763 (
            .O(N__49067),
            .I(N__49059));
    CascadeMux I__11762 (
            .O(N__49066),
            .I(N__49056));
    CascadeMux I__11761 (
            .O(N__49065),
            .I(N__49051));
    InMux I__11760 (
            .O(N__49064),
            .I(N__49045));
    InMux I__11759 (
            .O(N__49063),
            .I(N__49045));
    InMux I__11758 (
            .O(N__49062),
            .I(N__49042));
    InMux I__11757 (
            .O(N__49059),
            .I(N__49039));
    InMux I__11756 (
            .O(N__49056),
            .I(N__49036));
    InMux I__11755 (
            .O(N__49055),
            .I(N__49031));
    InMux I__11754 (
            .O(N__49054),
            .I(N__49031));
    InMux I__11753 (
            .O(N__49051),
            .I(N__49026));
    InMux I__11752 (
            .O(N__49050),
            .I(N__49026));
    LocalMux I__11751 (
            .O(N__49045),
            .I(N__49021));
    LocalMux I__11750 (
            .O(N__49042),
            .I(N__49021));
    LocalMux I__11749 (
            .O(N__49039),
            .I(N__49018));
    LocalMux I__11748 (
            .O(N__49036),
            .I(N__49015));
    LocalMux I__11747 (
            .O(N__49031),
            .I(N__49010));
    LocalMux I__11746 (
            .O(N__49026),
            .I(N__49010));
    Span4Mux_v I__11745 (
            .O(N__49021),
            .I(N__49007));
    Span4Mux_s3_h I__11744 (
            .O(N__49018),
            .I(N__49004));
    Span4Mux_s3_h I__11743 (
            .O(N__49015),
            .I(N__49001));
    Span4Mux_s3_h I__11742 (
            .O(N__49010),
            .I(N__48998));
    Span4Mux_h I__11741 (
            .O(N__49007),
            .I(N__48995));
    Span4Mux_h I__11740 (
            .O(N__49004),
            .I(N__48990));
    Span4Mux_h I__11739 (
            .O(N__49001),
            .I(N__48990));
    Span4Mux_h I__11738 (
            .O(N__48998),
            .I(N__48987));
    Odrv4 I__11737 (
            .O(N__48995),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ));
    Odrv4 I__11736 (
            .O(N__48990),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ));
    Odrv4 I__11735 (
            .O(N__48987),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ));
    InMux I__11734 (
            .O(N__48980),
            .I(N__48973));
    InMux I__11733 (
            .O(N__48979),
            .I(N__48968));
    InMux I__11732 (
            .O(N__48978),
            .I(N__48968));
    InMux I__11731 (
            .O(N__48977),
            .I(N__48963));
    InMux I__11730 (
            .O(N__48976),
            .I(N__48963));
    LocalMux I__11729 (
            .O(N__48973),
            .I(N__48953));
    LocalMux I__11728 (
            .O(N__48968),
            .I(N__48953));
    LocalMux I__11727 (
            .O(N__48963),
            .I(N__48950));
    InMux I__11726 (
            .O(N__48962),
            .I(N__48947));
    InMux I__11725 (
            .O(N__48961),
            .I(N__48940));
    InMux I__11724 (
            .O(N__48960),
            .I(N__48940));
    InMux I__11723 (
            .O(N__48959),
            .I(N__48940));
    InMux I__11722 (
            .O(N__48958),
            .I(N__48937));
    Span4Mux_v I__11721 (
            .O(N__48953),
            .I(N__48930));
    Span4Mux_s1_h I__11720 (
            .O(N__48950),
            .I(N__48930));
    LocalMux I__11719 (
            .O(N__48947),
            .I(N__48930));
    LocalMux I__11718 (
            .O(N__48940),
            .I(N__48927));
    LocalMux I__11717 (
            .O(N__48937),
            .I(N__48924));
    Span4Mux_h I__11716 (
            .O(N__48930),
            .I(N__48919));
    Span4Mux_h I__11715 (
            .O(N__48927),
            .I(N__48919));
    Span4Mux_h I__11714 (
            .O(N__48924),
            .I(N__48916));
    Span4Mux_h I__11713 (
            .O(N__48919),
            .I(N__48913));
    Odrv4 I__11712 (
            .O(N__48916),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__11711 (
            .O(N__48913),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    CascadeMux I__11710 (
            .O(N__48908),
            .I(N__48904));
    CascadeMux I__11709 (
            .O(N__48907),
            .I(N__48901));
    InMux I__11708 (
            .O(N__48904),
            .I(N__48897));
    InMux I__11707 (
            .O(N__48901),
            .I(N__48894));
    InMux I__11706 (
            .O(N__48900),
            .I(N__48891));
    LocalMux I__11705 (
            .O(N__48897),
            .I(N__48888));
    LocalMux I__11704 (
            .O(N__48894),
            .I(N__48883));
    LocalMux I__11703 (
            .O(N__48891),
            .I(N__48883));
    Span4Mux_s3_h I__11702 (
            .O(N__48888),
            .I(N__48878));
    Span4Mux_v I__11701 (
            .O(N__48883),
            .I(N__48878));
    Span4Mux_h I__11700 (
            .O(N__48878),
            .I(N__48875));
    Odrv4 I__11699 (
            .O(N__48875),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    InMux I__11698 (
            .O(N__48872),
            .I(N__48864));
    InMux I__11697 (
            .O(N__48871),
            .I(N__48859));
    InMux I__11696 (
            .O(N__48870),
            .I(N__48859));
    InMux I__11695 (
            .O(N__48869),
            .I(N__48852));
    InMux I__11694 (
            .O(N__48868),
            .I(N__48852));
    InMux I__11693 (
            .O(N__48867),
            .I(N__48852));
    LocalMux I__11692 (
            .O(N__48864),
            .I(N__48846));
    LocalMux I__11691 (
            .O(N__48859),
            .I(N__48846));
    LocalMux I__11690 (
            .O(N__48852),
            .I(N__48843));
    InMux I__11689 (
            .O(N__48851),
            .I(N__48840));
    Span4Mux_v I__11688 (
            .O(N__48846),
            .I(N__48833));
    Span4Mux_s1_h I__11687 (
            .O(N__48843),
            .I(N__48833));
    LocalMux I__11686 (
            .O(N__48840),
            .I(N__48833));
    Span4Mux_h I__11685 (
            .O(N__48833),
            .I(N__48830));
    Odrv4 I__11684 (
            .O(N__48830),
            .I(\current_shift_inst.PI_CTRL.N_159 ));
    InMux I__11683 (
            .O(N__48827),
            .I(N__48820));
    InMux I__11682 (
            .O(N__48826),
            .I(N__48820));
    InMux I__11681 (
            .O(N__48825),
            .I(N__48817));
    LocalMux I__11680 (
            .O(N__48820),
            .I(pwm_duty_input_9));
    LocalMux I__11679 (
            .O(N__48817),
            .I(pwm_duty_input_9));
    InMux I__11678 (
            .O(N__48812),
            .I(N__48809));
    LocalMux I__11677 (
            .O(N__48809),
            .I(N__48643));
    ClkMux I__11676 (
            .O(N__48808),
            .I(N__48314));
    ClkMux I__11675 (
            .O(N__48807),
            .I(N__48314));
    ClkMux I__11674 (
            .O(N__48806),
            .I(N__48314));
    ClkMux I__11673 (
            .O(N__48805),
            .I(N__48314));
    ClkMux I__11672 (
            .O(N__48804),
            .I(N__48314));
    ClkMux I__11671 (
            .O(N__48803),
            .I(N__48314));
    ClkMux I__11670 (
            .O(N__48802),
            .I(N__48314));
    ClkMux I__11669 (
            .O(N__48801),
            .I(N__48314));
    ClkMux I__11668 (
            .O(N__48800),
            .I(N__48314));
    ClkMux I__11667 (
            .O(N__48799),
            .I(N__48314));
    ClkMux I__11666 (
            .O(N__48798),
            .I(N__48314));
    ClkMux I__11665 (
            .O(N__48797),
            .I(N__48314));
    ClkMux I__11664 (
            .O(N__48796),
            .I(N__48314));
    ClkMux I__11663 (
            .O(N__48795),
            .I(N__48314));
    ClkMux I__11662 (
            .O(N__48794),
            .I(N__48314));
    ClkMux I__11661 (
            .O(N__48793),
            .I(N__48314));
    ClkMux I__11660 (
            .O(N__48792),
            .I(N__48314));
    ClkMux I__11659 (
            .O(N__48791),
            .I(N__48314));
    ClkMux I__11658 (
            .O(N__48790),
            .I(N__48314));
    ClkMux I__11657 (
            .O(N__48789),
            .I(N__48314));
    ClkMux I__11656 (
            .O(N__48788),
            .I(N__48314));
    ClkMux I__11655 (
            .O(N__48787),
            .I(N__48314));
    ClkMux I__11654 (
            .O(N__48786),
            .I(N__48314));
    ClkMux I__11653 (
            .O(N__48785),
            .I(N__48314));
    ClkMux I__11652 (
            .O(N__48784),
            .I(N__48314));
    ClkMux I__11651 (
            .O(N__48783),
            .I(N__48314));
    ClkMux I__11650 (
            .O(N__48782),
            .I(N__48314));
    ClkMux I__11649 (
            .O(N__48781),
            .I(N__48314));
    ClkMux I__11648 (
            .O(N__48780),
            .I(N__48314));
    ClkMux I__11647 (
            .O(N__48779),
            .I(N__48314));
    ClkMux I__11646 (
            .O(N__48778),
            .I(N__48314));
    ClkMux I__11645 (
            .O(N__48777),
            .I(N__48314));
    ClkMux I__11644 (
            .O(N__48776),
            .I(N__48314));
    ClkMux I__11643 (
            .O(N__48775),
            .I(N__48314));
    ClkMux I__11642 (
            .O(N__48774),
            .I(N__48314));
    ClkMux I__11641 (
            .O(N__48773),
            .I(N__48314));
    ClkMux I__11640 (
            .O(N__48772),
            .I(N__48314));
    ClkMux I__11639 (
            .O(N__48771),
            .I(N__48314));
    ClkMux I__11638 (
            .O(N__48770),
            .I(N__48314));
    ClkMux I__11637 (
            .O(N__48769),
            .I(N__48314));
    ClkMux I__11636 (
            .O(N__48768),
            .I(N__48314));
    ClkMux I__11635 (
            .O(N__48767),
            .I(N__48314));
    ClkMux I__11634 (
            .O(N__48766),
            .I(N__48314));
    ClkMux I__11633 (
            .O(N__48765),
            .I(N__48314));
    ClkMux I__11632 (
            .O(N__48764),
            .I(N__48314));
    ClkMux I__11631 (
            .O(N__48763),
            .I(N__48314));
    ClkMux I__11630 (
            .O(N__48762),
            .I(N__48314));
    ClkMux I__11629 (
            .O(N__48761),
            .I(N__48314));
    ClkMux I__11628 (
            .O(N__48760),
            .I(N__48314));
    ClkMux I__11627 (
            .O(N__48759),
            .I(N__48314));
    ClkMux I__11626 (
            .O(N__48758),
            .I(N__48314));
    ClkMux I__11625 (
            .O(N__48757),
            .I(N__48314));
    ClkMux I__11624 (
            .O(N__48756),
            .I(N__48314));
    ClkMux I__11623 (
            .O(N__48755),
            .I(N__48314));
    ClkMux I__11622 (
            .O(N__48754),
            .I(N__48314));
    ClkMux I__11621 (
            .O(N__48753),
            .I(N__48314));
    ClkMux I__11620 (
            .O(N__48752),
            .I(N__48314));
    ClkMux I__11619 (
            .O(N__48751),
            .I(N__48314));
    ClkMux I__11618 (
            .O(N__48750),
            .I(N__48314));
    ClkMux I__11617 (
            .O(N__48749),
            .I(N__48314));
    ClkMux I__11616 (
            .O(N__48748),
            .I(N__48314));
    ClkMux I__11615 (
            .O(N__48747),
            .I(N__48314));
    ClkMux I__11614 (
            .O(N__48746),
            .I(N__48314));
    ClkMux I__11613 (
            .O(N__48745),
            .I(N__48314));
    ClkMux I__11612 (
            .O(N__48744),
            .I(N__48314));
    ClkMux I__11611 (
            .O(N__48743),
            .I(N__48314));
    ClkMux I__11610 (
            .O(N__48742),
            .I(N__48314));
    ClkMux I__11609 (
            .O(N__48741),
            .I(N__48314));
    ClkMux I__11608 (
            .O(N__48740),
            .I(N__48314));
    ClkMux I__11607 (
            .O(N__48739),
            .I(N__48314));
    ClkMux I__11606 (
            .O(N__48738),
            .I(N__48314));
    ClkMux I__11605 (
            .O(N__48737),
            .I(N__48314));
    ClkMux I__11604 (
            .O(N__48736),
            .I(N__48314));
    ClkMux I__11603 (
            .O(N__48735),
            .I(N__48314));
    ClkMux I__11602 (
            .O(N__48734),
            .I(N__48314));
    ClkMux I__11601 (
            .O(N__48733),
            .I(N__48314));
    ClkMux I__11600 (
            .O(N__48732),
            .I(N__48314));
    ClkMux I__11599 (
            .O(N__48731),
            .I(N__48314));
    ClkMux I__11598 (
            .O(N__48730),
            .I(N__48314));
    ClkMux I__11597 (
            .O(N__48729),
            .I(N__48314));
    ClkMux I__11596 (
            .O(N__48728),
            .I(N__48314));
    ClkMux I__11595 (
            .O(N__48727),
            .I(N__48314));
    ClkMux I__11594 (
            .O(N__48726),
            .I(N__48314));
    ClkMux I__11593 (
            .O(N__48725),
            .I(N__48314));
    ClkMux I__11592 (
            .O(N__48724),
            .I(N__48314));
    ClkMux I__11591 (
            .O(N__48723),
            .I(N__48314));
    ClkMux I__11590 (
            .O(N__48722),
            .I(N__48314));
    ClkMux I__11589 (
            .O(N__48721),
            .I(N__48314));
    ClkMux I__11588 (
            .O(N__48720),
            .I(N__48314));
    ClkMux I__11587 (
            .O(N__48719),
            .I(N__48314));
    ClkMux I__11586 (
            .O(N__48718),
            .I(N__48314));
    ClkMux I__11585 (
            .O(N__48717),
            .I(N__48314));
    ClkMux I__11584 (
            .O(N__48716),
            .I(N__48314));
    ClkMux I__11583 (
            .O(N__48715),
            .I(N__48314));
    ClkMux I__11582 (
            .O(N__48714),
            .I(N__48314));
    ClkMux I__11581 (
            .O(N__48713),
            .I(N__48314));
    ClkMux I__11580 (
            .O(N__48712),
            .I(N__48314));
    ClkMux I__11579 (
            .O(N__48711),
            .I(N__48314));
    ClkMux I__11578 (
            .O(N__48710),
            .I(N__48314));
    ClkMux I__11577 (
            .O(N__48709),
            .I(N__48314));
    ClkMux I__11576 (
            .O(N__48708),
            .I(N__48314));
    ClkMux I__11575 (
            .O(N__48707),
            .I(N__48314));
    ClkMux I__11574 (
            .O(N__48706),
            .I(N__48314));
    ClkMux I__11573 (
            .O(N__48705),
            .I(N__48314));
    ClkMux I__11572 (
            .O(N__48704),
            .I(N__48314));
    ClkMux I__11571 (
            .O(N__48703),
            .I(N__48314));
    ClkMux I__11570 (
            .O(N__48702),
            .I(N__48314));
    ClkMux I__11569 (
            .O(N__48701),
            .I(N__48314));
    ClkMux I__11568 (
            .O(N__48700),
            .I(N__48314));
    ClkMux I__11567 (
            .O(N__48699),
            .I(N__48314));
    ClkMux I__11566 (
            .O(N__48698),
            .I(N__48314));
    ClkMux I__11565 (
            .O(N__48697),
            .I(N__48314));
    ClkMux I__11564 (
            .O(N__48696),
            .I(N__48314));
    ClkMux I__11563 (
            .O(N__48695),
            .I(N__48314));
    ClkMux I__11562 (
            .O(N__48694),
            .I(N__48314));
    ClkMux I__11561 (
            .O(N__48693),
            .I(N__48314));
    ClkMux I__11560 (
            .O(N__48692),
            .I(N__48314));
    ClkMux I__11559 (
            .O(N__48691),
            .I(N__48314));
    ClkMux I__11558 (
            .O(N__48690),
            .I(N__48314));
    ClkMux I__11557 (
            .O(N__48689),
            .I(N__48314));
    ClkMux I__11556 (
            .O(N__48688),
            .I(N__48314));
    ClkMux I__11555 (
            .O(N__48687),
            .I(N__48314));
    ClkMux I__11554 (
            .O(N__48686),
            .I(N__48314));
    ClkMux I__11553 (
            .O(N__48685),
            .I(N__48314));
    ClkMux I__11552 (
            .O(N__48684),
            .I(N__48314));
    ClkMux I__11551 (
            .O(N__48683),
            .I(N__48314));
    ClkMux I__11550 (
            .O(N__48682),
            .I(N__48314));
    ClkMux I__11549 (
            .O(N__48681),
            .I(N__48314));
    ClkMux I__11548 (
            .O(N__48680),
            .I(N__48314));
    ClkMux I__11547 (
            .O(N__48679),
            .I(N__48314));
    ClkMux I__11546 (
            .O(N__48678),
            .I(N__48314));
    ClkMux I__11545 (
            .O(N__48677),
            .I(N__48314));
    ClkMux I__11544 (
            .O(N__48676),
            .I(N__48314));
    ClkMux I__11543 (
            .O(N__48675),
            .I(N__48314));
    ClkMux I__11542 (
            .O(N__48674),
            .I(N__48314));
    ClkMux I__11541 (
            .O(N__48673),
            .I(N__48314));
    ClkMux I__11540 (
            .O(N__48672),
            .I(N__48314));
    ClkMux I__11539 (
            .O(N__48671),
            .I(N__48314));
    ClkMux I__11538 (
            .O(N__48670),
            .I(N__48314));
    ClkMux I__11537 (
            .O(N__48669),
            .I(N__48314));
    ClkMux I__11536 (
            .O(N__48668),
            .I(N__48314));
    ClkMux I__11535 (
            .O(N__48667),
            .I(N__48314));
    ClkMux I__11534 (
            .O(N__48666),
            .I(N__48314));
    ClkMux I__11533 (
            .O(N__48665),
            .I(N__48314));
    ClkMux I__11532 (
            .O(N__48664),
            .I(N__48314));
    ClkMux I__11531 (
            .O(N__48663),
            .I(N__48314));
    ClkMux I__11530 (
            .O(N__48662),
            .I(N__48314));
    ClkMux I__11529 (
            .O(N__48661),
            .I(N__48314));
    ClkMux I__11528 (
            .O(N__48660),
            .I(N__48314));
    ClkMux I__11527 (
            .O(N__48659),
            .I(N__48314));
    ClkMux I__11526 (
            .O(N__48658),
            .I(N__48314));
    ClkMux I__11525 (
            .O(N__48657),
            .I(N__48314));
    ClkMux I__11524 (
            .O(N__48656),
            .I(N__48314));
    ClkMux I__11523 (
            .O(N__48655),
            .I(N__48314));
    ClkMux I__11522 (
            .O(N__48654),
            .I(N__48314));
    ClkMux I__11521 (
            .O(N__48653),
            .I(N__48314));
    ClkMux I__11520 (
            .O(N__48652),
            .I(N__48314));
    ClkMux I__11519 (
            .O(N__48651),
            .I(N__48314));
    ClkMux I__11518 (
            .O(N__48650),
            .I(N__48314));
    ClkMux I__11517 (
            .O(N__48649),
            .I(N__48314));
    ClkMux I__11516 (
            .O(N__48648),
            .I(N__48314));
    ClkMux I__11515 (
            .O(N__48647),
            .I(N__48314));
    ClkMux I__11514 (
            .O(N__48646),
            .I(N__48314));
    Glb2LocalMux I__11513 (
            .O(N__48643),
            .I(N__48314));
    GlobalMux I__11512 (
            .O(N__48314),
            .I(clock_output_0));
    InMux I__11511 (
            .O(N__48311),
            .I(N__48305));
    InMux I__11510 (
            .O(N__48310),
            .I(N__48302));
    InMux I__11509 (
            .O(N__48309),
            .I(N__48299));
    InMux I__11508 (
            .O(N__48308),
            .I(N__48296));
    LocalMux I__11507 (
            .O(N__48305),
            .I(N__48293));
    LocalMux I__11506 (
            .O(N__48302),
            .I(N__48290));
    LocalMux I__11505 (
            .O(N__48299),
            .I(N__48287));
    LocalMux I__11504 (
            .O(N__48296),
            .I(N__48283));
    Glb2LocalMux I__11503 (
            .O(N__48293),
            .I(N__47786));
    Glb2LocalMux I__11502 (
            .O(N__48290),
            .I(N__47786));
    Glb2LocalMux I__11501 (
            .O(N__48287),
            .I(N__47786));
    SRMux I__11500 (
            .O(N__48286),
            .I(N__47786));
    Glb2LocalMux I__11499 (
            .O(N__48283),
            .I(N__47786));
    SRMux I__11498 (
            .O(N__48282),
            .I(N__47786));
    SRMux I__11497 (
            .O(N__48281),
            .I(N__47786));
    SRMux I__11496 (
            .O(N__48280),
            .I(N__47786));
    SRMux I__11495 (
            .O(N__48279),
            .I(N__47786));
    SRMux I__11494 (
            .O(N__48278),
            .I(N__47786));
    SRMux I__11493 (
            .O(N__48277),
            .I(N__47786));
    SRMux I__11492 (
            .O(N__48276),
            .I(N__47786));
    SRMux I__11491 (
            .O(N__48275),
            .I(N__47786));
    SRMux I__11490 (
            .O(N__48274),
            .I(N__47786));
    SRMux I__11489 (
            .O(N__48273),
            .I(N__47786));
    SRMux I__11488 (
            .O(N__48272),
            .I(N__47786));
    SRMux I__11487 (
            .O(N__48271),
            .I(N__47786));
    SRMux I__11486 (
            .O(N__48270),
            .I(N__47786));
    SRMux I__11485 (
            .O(N__48269),
            .I(N__47786));
    SRMux I__11484 (
            .O(N__48268),
            .I(N__47786));
    SRMux I__11483 (
            .O(N__48267),
            .I(N__47786));
    SRMux I__11482 (
            .O(N__48266),
            .I(N__47786));
    SRMux I__11481 (
            .O(N__48265),
            .I(N__47786));
    SRMux I__11480 (
            .O(N__48264),
            .I(N__47786));
    SRMux I__11479 (
            .O(N__48263),
            .I(N__47786));
    SRMux I__11478 (
            .O(N__48262),
            .I(N__47786));
    SRMux I__11477 (
            .O(N__48261),
            .I(N__47786));
    SRMux I__11476 (
            .O(N__48260),
            .I(N__47786));
    SRMux I__11475 (
            .O(N__48259),
            .I(N__47786));
    SRMux I__11474 (
            .O(N__48258),
            .I(N__47786));
    SRMux I__11473 (
            .O(N__48257),
            .I(N__47786));
    SRMux I__11472 (
            .O(N__48256),
            .I(N__47786));
    SRMux I__11471 (
            .O(N__48255),
            .I(N__47786));
    SRMux I__11470 (
            .O(N__48254),
            .I(N__47786));
    SRMux I__11469 (
            .O(N__48253),
            .I(N__47786));
    SRMux I__11468 (
            .O(N__48252),
            .I(N__47786));
    SRMux I__11467 (
            .O(N__48251),
            .I(N__47786));
    SRMux I__11466 (
            .O(N__48250),
            .I(N__47786));
    SRMux I__11465 (
            .O(N__48249),
            .I(N__47786));
    SRMux I__11464 (
            .O(N__48248),
            .I(N__47786));
    SRMux I__11463 (
            .O(N__48247),
            .I(N__47786));
    SRMux I__11462 (
            .O(N__48246),
            .I(N__47786));
    SRMux I__11461 (
            .O(N__48245),
            .I(N__47786));
    SRMux I__11460 (
            .O(N__48244),
            .I(N__47786));
    SRMux I__11459 (
            .O(N__48243),
            .I(N__47786));
    SRMux I__11458 (
            .O(N__48242),
            .I(N__47786));
    SRMux I__11457 (
            .O(N__48241),
            .I(N__47786));
    SRMux I__11456 (
            .O(N__48240),
            .I(N__47786));
    SRMux I__11455 (
            .O(N__48239),
            .I(N__47786));
    SRMux I__11454 (
            .O(N__48238),
            .I(N__47786));
    SRMux I__11453 (
            .O(N__48237),
            .I(N__47786));
    SRMux I__11452 (
            .O(N__48236),
            .I(N__47786));
    SRMux I__11451 (
            .O(N__48235),
            .I(N__47786));
    SRMux I__11450 (
            .O(N__48234),
            .I(N__47786));
    SRMux I__11449 (
            .O(N__48233),
            .I(N__47786));
    SRMux I__11448 (
            .O(N__48232),
            .I(N__47786));
    SRMux I__11447 (
            .O(N__48231),
            .I(N__47786));
    SRMux I__11446 (
            .O(N__48230),
            .I(N__47786));
    SRMux I__11445 (
            .O(N__48229),
            .I(N__47786));
    SRMux I__11444 (
            .O(N__48228),
            .I(N__47786));
    SRMux I__11443 (
            .O(N__48227),
            .I(N__47786));
    SRMux I__11442 (
            .O(N__48226),
            .I(N__47786));
    SRMux I__11441 (
            .O(N__48225),
            .I(N__47786));
    SRMux I__11440 (
            .O(N__48224),
            .I(N__47786));
    SRMux I__11439 (
            .O(N__48223),
            .I(N__47786));
    SRMux I__11438 (
            .O(N__48222),
            .I(N__47786));
    SRMux I__11437 (
            .O(N__48221),
            .I(N__47786));
    SRMux I__11436 (
            .O(N__48220),
            .I(N__47786));
    SRMux I__11435 (
            .O(N__48219),
            .I(N__47786));
    SRMux I__11434 (
            .O(N__48218),
            .I(N__47786));
    SRMux I__11433 (
            .O(N__48217),
            .I(N__47786));
    SRMux I__11432 (
            .O(N__48216),
            .I(N__47786));
    SRMux I__11431 (
            .O(N__48215),
            .I(N__47786));
    SRMux I__11430 (
            .O(N__48214),
            .I(N__47786));
    SRMux I__11429 (
            .O(N__48213),
            .I(N__47786));
    SRMux I__11428 (
            .O(N__48212),
            .I(N__47786));
    SRMux I__11427 (
            .O(N__48211),
            .I(N__47786));
    SRMux I__11426 (
            .O(N__48210),
            .I(N__47786));
    SRMux I__11425 (
            .O(N__48209),
            .I(N__47786));
    SRMux I__11424 (
            .O(N__48208),
            .I(N__47786));
    SRMux I__11423 (
            .O(N__48207),
            .I(N__47786));
    SRMux I__11422 (
            .O(N__48206),
            .I(N__47786));
    SRMux I__11421 (
            .O(N__48205),
            .I(N__47786));
    SRMux I__11420 (
            .O(N__48204),
            .I(N__47786));
    SRMux I__11419 (
            .O(N__48203),
            .I(N__47786));
    SRMux I__11418 (
            .O(N__48202),
            .I(N__47786));
    SRMux I__11417 (
            .O(N__48201),
            .I(N__47786));
    SRMux I__11416 (
            .O(N__48200),
            .I(N__47786));
    SRMux I__11415 (
            .O(N__48199),
            .I(N__47786));
    SRMux I__11414 (
            .O(N__48198),
            .I(N__47786));
    SRMux I__11413 (
            .O(N__48197),
            .I(N__47786));
    SRMux I__11412 (
            .O(N__48196),
            .I(N__47786));
    SRMux I__11411 (
            .O(N__48195),
            .I(N__47786));
    SRMux I__11410 (
            .O(N__48194),
            .I(N__47786));
    SRMux I__11409 (
            .O(N__48193),
            .I(N__47786));
    SRMux I__11408 (
            .O(N__48192),
            .I(N__47786));
    SRMux I__11407 (
            .O(N__48191),
            .I(N__47786));
    SRMux I__11406 (
            .O(N__48190),
            .I(N__47786));
    SRMux I__11405 (
            .O(N__48189),
            .I(N__47786));
    SRMux I__11404 (
            .O(N__48188),
            .I(N__47786));
    SRMux I__11403 (
            .O(N__48187),
            .I(N__47786));
    SRMux I__11402 (
            .O(N__48186),
            .I(N__47786));
    SRMux I__11401 (
            .O(N__48185),
            .I(N__47786));
    SRMux I__11400 (
            .O(N__48184),
            .I(N__47786));
    SRMux I__11399 (
            .O(N__48183),
            .I(N__47786));
    SRMux I__11398 (
            .O(N__48182),
            .I(N__47786));
    SRMux I__11397 (
            .O(N__48181),
            .I(N__47786));
    SRMux I__11396 (
            .O(N__48180),
            .I(N__47786));
    SRMux I__11395 (
            .O(N__48179),
            .I(N__47786));
    SRMux I__11394 (
            .O(N__48178),
            .I(N__47786));
    SRMux I__11393 (
            .O(N__48177),
            .I(N__47786));
    SRMux I__11392 (
            .O(N__48176),
            .I(N__47786));
    SRMux I__11391 (
            .O(N__48175),
            .I(N__47786));
    SRMux I__11390 (
            .O(N__48174),
            .I(N__47786));
    SRMux I__11389 (
            .O(N__48173),
            .I(N__47786));
    SRMux I__11388 (
            .O(N__48172),
            .I(N__47786));
    SRMux I__11387 (
            .O(N__48171),
            .I(N__47786));
    SRMux I__11386 (
            .O(N__48170),
            .I(N__47786));
    SRMux I__11385 (
            .O(N__48169),
            .I(N__47786));
    SRMux I__11384 (
            .O(N__48168),
            .I(N__47786));
    SRMux I__11383 (
            .O(N__48167),
            .I(N__47786));
    SRMux I__11382 (
            .O(N__48166),
            .I(N__47786));
    SRMux I__11381 (
            .O(N__48165),
            .I(N__47786));
    SRMux I__11380 (
            .O(N__48164),
            .I(N__47786));
    SRMux I__11379 (
            .O(N__48163),
            .I(N__47786));
    SRMux I__11378 (
            .O(N__48162),
            .I(N__47786));
    SRMux I__11377 (
            .O(N__48161),
            .I(N__47786));
    SRMux I__11376 (
            .O(N__48160),
            .I(N__47786));
    SRMux I__11375 (
            .O(N__48159),
            .I(N__47786));
    SRMux I__11374 (
            .O(N__48158),
            .I(N__47786));
    SRMux I__11373 (
            .O(N__48157),
            .I(N__47786));
    SRMux I__11372 (
            .O(N__48156),
            .I(N__47786));
    SRMux I__11371 (
            .O(N__48155),
            .I(N__47786));
    SRMux I__11370 (
            .O(N__48154),
            .I(N__47786));
    SRMux I__11369 (
            .O(N__48153),
            .I(N__47786));
    SRMux I__11368 (
            .O(N__48152),
            .I(N__47786));
    SRMux I__11367 (
            .O(N__48151),
            .I(N__47786));
    SRMux I__11366 (
            .O(N__48150),
            .I(N__47786));
    SRMux I__11365 (
            .O(N__48149),
            .I(N__47786));
    SRMux I__11364 (
            .O(N__48148),
            .I(N__47786));
    SRMux I__11363 (
            .O(N__48147),
            .I(N__47786));
    SRMux I__11362 (
            .O(N__48146),
            .I(N__47786));
    SRMux I__11361 (
            .O(N__48145),
            .I(N__47786));
    SRMux I__11360 (
            .O(N__48144),
            .I(N__47786));
    SRMux I__11359 (
            .O(N__48143),
            .I(N__47786));
    SRMux I__11358 (
            .O(N__48142),
            .I(N__47786));
    SRMux I__11357 (
            .O(N__48141),
            .I(N__47786));
    SRMux I__11356 (
            .O(N__48140),
            .I(N__47786));
    SRMux I__11355 (
            .O(N__48139),
            .I(N__47786));
    SRMux I__11354 (
            .O(N__48138),
            .I(N__47786));
    SRMux I__11353 (
            .O(N__48137),
            .I(N__47786));
    SRMux I__11352 (
            .O(N__48136),
            .I(N__47786));
    SRMux I__11351 (
            .O(N__48135),
            .I(N__47786));
    SRMux I__11350 (
            .O(N__48134),
            .I(N__47786));
    SRMux I__11349 (
            .O(N__48133),
            .I(N__47786));
    SRMux I__11348 (
            .O(N__48132),
            .I(N__47786));
    SRMux I__11347 (
            .O(N__48131),
            .I(N__47786));
    SRMux I__11346 (
            .O(N__48130),
            .I(N__47786));
    SRMux I__11345 (
            .O(N__48129),
            .I(N__47786));
    SRMux I__11344 (
            .O(N__48128),
            .I(N__47786));
    SRMux I__11343 (
            .O(N__48127),
            .I(N__47786));
    SRMux I__11342 (
            .O(N__48126),
            .I(N__47786));
    SRMux I__11341 (
            .O(N__48125),
            .I(N__47786));
    SRMux I__11340 (
            .O(N__48124),
            .I(N__47786));
    SRMux I__11339 (
            .O(N__48123),
            .I(N__47786));
    SRMux I__11338 (
            .O(N__48122),
            .I(N__47786));
    SRMux I__11337 (
            .O(N__48121),
            .I(N__47786));
    GlobalMux I__11336 (
            .O(N__47786),
            .I(N__47783));
    gio2CtrlBuf I__11335 (
            .O(N__47783),
            .I(red_c_g));
    InMux I__11334 (
            .O(N__47780),
            .I(N__47777));
    LocalMux I__11333 (
            .O(N__47777),
            .I(\pwm_generator_inst.un1_duty_inputlt3 ));
    InMux I__11332 (
            .O(N__47774),
            .I(N__47765));
    InMux I__11331 (
            .O(N__47773),
            .I(N__47765));
    InMux I__11330 (
            .O(N__47772),
            .I(N__47765));
    LocalMux I__11329 (
            .O(N__47765),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    CascadeMux I__11328 (
            .O(N__47762),
            .I(N__47759));
    InMux I__11327 (
            .O(N__47759),
            .I(N__47754));
    InMux I__11326 (
            .O(N__47758),
            .I(N__47749));
    InMux I__11325 (
            .O(N__47757),
            .I(N__47749));
    LocalMux I__11324 (
            .O(N__47754),
            .I(N__47746));
    LocalMux I__11323 (
            .O(N__47749),
            .I(N__47743));
    Span4Mux_v I__11322 (
            .O(N__47746),
            .I(N__47740));
    Span4Mux_h I__11321 (
            .O(N__47743),
            .I(N__47737));
    Sp12to4 I__11320 (
            .O(N__47740),
            .I(N__47734));
    Span4Mux_h I__11319 (
            .O(N__47737),
            .I(N__47731));
    Odrv12 I__11318 (
            .O(N__47734),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    Odrv4 I__11317 (
            .O(N__47731),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    InMux I__11316 (
            .O(N__47726),
            .I(N__47723));
    LocalMux I__11315 (
            .O(N__47723),
            .I(N__47718));
    InMux I__11314 (
            .O(N__47722),
            .I(N__47713));
    InMux I__11313 (
            .O(N__47721),
            .I(N__47713));
    Span4Mux_s0_h I__11312 (
            .O(N__47718),
            .I(N__47710));
    LocalMux I__11311 (
            .O(N__47713),
            .I(pwm_duty_input_7));
    Odrv4 I__11310 (
            .O(N__47710),
            .I(pwm_duty_input_7));
    CascadeMux I__11309 (
            .O(N__47705),
            .I(N__47701));
    CascadeMux I__11308 (
            .O(N__47704),
            .I(N__47698));
    InMux I__11307 (
            .O(N__47701),
            .I(N__47695));
    InMux I__11306 (
            .O(N__47698),
            .I(N__47692));
    LocalMux I__11305 (
            .O(N__47695),
            .I(N__47688));
    LocalMux I__11304 (
            .O(N__47692),
            .I(N__47685));
    InMux I__11303 (
            .O(N__47691),
            .I(N__47682));
    Span4Mux_h I__11302 (
            .O(N__47688),
            .I(N__47679));
    Span12Mux_s1_h I__11301 (
            .O(N__47685),
            .I(N__47674));
    LocalMux I__11300 (
            .O(N__47682),
            .I(N__47674));
    Span4Mux_h I__11299 (
            .O(N__47679),
            .I(N__47671));
    Odrv12 I__11298 (
            .O(N__47674),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    Odrv4 I__11297 (
            .O(N__47671),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    InMux I__11296 (
            .O(N__47666),
            .I(N__47661));
    InMux I__11295 (
            .O(N__47665),
            .I(N__47656));
    InMux I__11294 (
            .O(N__47664),
            .I(N__47656));
    LocalMux I__11293 (
            .O(N__47661),
            .I(N__47653));
    LocalMux I__11292 (
            .O(N__47656),
            .I(pwm_duty_input_8));
    Odrv4 I__11291 (
            .O(N__47653),
            .I(pwm_duty_input_8));
    InMux I__11290 (
            .O(N__47648),
            .I(N__47645));
    LocalMux I__11289 (
            .O(N__47645),
            .I(N__47642));
    Span4Mux_h I__11288 (
            .O(N__47642),
            .I(N__47639));
    Odrv4 I__11287 (
            .O(N__47639),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    InMux I__11286 (
            .O(N__47636),
            .I(N__47632));
    InMux I__11285 (
            .O(N__47635),
            .I(N__47629));
    LocalMux I__11284 (
            .O(N__47632),
            .I(N__47626));
    LocalMux I__11283 (
            .O(N__47629),
            .I(pwm_duty_input_0));
    Odrv4 I__11282 (
            .O(N__47626),
            .I(pwm_duty_input_0));
    InMux I__11281 (
            .O(N__47621),
            .I(N__47617));
    InMux I__11280 (
            .O(N__47620),
            .I(N__47614));
    LocalMux I__11279 (
            .O(N__47617),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ));
    LocalMux I__11278 (
            .O(N__47614),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ));
    InMux I__11277 (
            .O(N__47609),
            .I(N__47606));
    LocalMux I__11276 (
            .O(N__47606),
            .I(N__47601));
    InMux I__11275 (
            .O(N__47605),
            .I(N__47598));
    InMux I__11274 (
            .O(N__47604),
            .I(N__47595));
    Span4Mux_v I__11273 (
            .O(N__47601),
            .I(N__47590));
    LocalMux I__11272 (
            .O(N__47598),
            .I(N__47590));
    LocalMux I__11271 (
            .O(N__47595),
            .I(N__47587));
    Span4Mux_h I__11270 (
            .O(N__47590),
            .I(N__47584));
    Span12Mux_s4_h I__11269 (
            .O(N__47587),
            .I(N__47581));
    Span4Mux_h I__11268 (
            .O(N__47584),
            .I(N__47578));
    Odrv12 I__11267 (
            .O(N__47581),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    Odrv4 I__11266 (
            .O(N__47578),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__11265 (
            .O(N__47573),
            .I(N__47568));
    InMux I__11264 (
            .O(N__47572),
            .I(N__47565));
    InMux I__11263 (
            .O(N__47571),
            .I(N__47562));
    LocalMux I__11262 (
            .O(N__47568),
            .I(N__47559));
    LocalMux I__11261 (
            .O(N__47565),
            .I(N__47556));
    LocalMux I__11260 (
            .O(N__47562),
            .I(N__47553));
    Odrv4 I__11259 (
            .O(N__47559),
            .I(pwm_duty_input_3));
    Odrv4 I__11258 (
            .O(N__47556),
            .I(pwm_duty_input_3));
    Odrv4 I__11257 (
            .O(N__47553),
            .I(pwm_duty_input_3));
    InMux I__11256 (
            .O(N__47546),
            .I(N__47532));
    InMux I__11255 (
            .O(N__47545),
            .I(N__47532));
    InMux I__11254 (
            .O(N__47544),
            .I(N__47517));
    InMux I__11253 (
            .O(N__47543),
            .I(N__47517));
    InMux I__11252 (
            .O(N__47542),
            .I(N__47517));
    InMux I__11251 (
            .O(N__47541),
            .I(N__47517));
    InMux I__11250 (
            .O(N__47540),
            .I(N__47517));
    InMux I__11249 (
            .O(N__47539),
            .I(N__47517));
    InMux I__11248 (
            .O(N__47538),
            .I(N__47517));
    InMux I__11247 (
            .O(N__47537),
            .I(N__47514));
    LocalMux I__11246 (
            .O(N__47532),
            .I(N__47509));
    LocalMux I__11245 (
            .O(N__47517),
            .I(N__47509));
    LocalMux I__11244 (
            .O(N__47514),
            .I(N__47504));
    Span12Mux_s7_v I__11243 (
            .O(N__47509),
            .I(N__47504));
    Odrv12 I__11242 (
            .O(N__47504),
            .I(\pwm_generator_inst.N_16 ));
    InMux I__11241 (
            .O(N__47501),
            .I(N__47498));
    LocalMux I__11240 (
            .O(N__47498),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4 ));
    CascadeMux I__11239 (
            .O(N__47495),
            .I(\current_shift_inst.PI_CTRL.N_27_cascade_ ));
    InMux I__11238 (
            .O(N__47492),
            .I(N__47489));
    LocalMux I__11237 (
            .O(N__47489),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0 ));
    InMux I__11236 (
            .O(N__47486),
            .I(N__47483));
    LocalMux I__11235 (
            .O(N__47483),
            .I(\current_shift_inst.PI_CTRL.N_98 ));
    CascadeMux I__11234 (
            .O(N__47480),
            .I(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ));
    InMux I__11233 (
            .O(N__47477),
            .I(N__47464));
    InMux I__11232 (
            .O(N__47476),
            .I(N__47464));
    InMux I__11231 (
            .O(N__47475),
            .I(N__47448));
    InMux I__11230 (
            .O(N__47474),
            .I(N__47448));
    InMux I__11229 (
            .O(N__47473),
            .I(N__47448));
    InMux I__11228 (
            .O(N__47472),
            .I(N__47448));
    InMux I__11227 (
            .O(N__47471),
            .I(N__47448));
    InMux I__11226 (
            .O(N__47470),
            .I(N__47448));
    InMux I__11225 (
            .O(N__47469),
            .I(N__47448));
    LocalMux I__11224 (
            .O(N__47464),
            .I(N__47445));
    InMux I__11223 (
            .O(N__47463),
            .I(N__47442));
    LocalMux I__11222 (
            .O(N__47448),
            .I(N__47439));
    Span4Mux_v I__11221 (
            .O(N__47445),
            .I(N__47434));
    LocalMux I__11220 (
            .O(N__47442),
            .I(N__47434));
    Span4Mux_h I__11219 (
            .O(N__47439),
            .I(N__47431));
    Span4Mux_h I__11218 (
            .O(N__47434),
            .I(N__47428));
    Span4Mux_h I__11217 (
            .O(N__47431),
            .I(N__47425));
    Sp12to4 I__11216 (
            .O(N__47428),
            .I(N__47422));
    Span4Mux_h I__11215 (
            .O(N__47425),
            .I(N__47419));
    Odrv12 I__11214 (
            .O(N__47422),
            .I(\pwm_generator_inst.N_17 ));
    Odrv4 I__11213 (
            .O(N__47419),
            .I(\pwm_generator_inst.N_17 ));
    CascadeMux I__11212 (
            .O(N__47414),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ));
    InMux I__11211 (
            .O(N__47411),
            .I(N__47408));
    LocalMux I__11210 (
            .O(N__47408),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ));
    CascadeMux I__11209 (
            .O(N__47405),
            .I(N__47401));
    InMux I__11208 (
            .O(N__47404),
            .I(N__47396));
    InMux I__11207 (
            .O(N__47401),
            .I(N__47396));
    LocalMux I__11206 (
            .O(N__47396),
            .I(N__47392));
    InMux I__11205 (
            .O(N__47395),
            .I(N__47389));
    Span4Mux_h I__11204 (
            .O(N__47392),
            .I(N__47386));
    LocalMux I__11203 (
            .O(N__47389),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ));
    Odrv4 I__11202 (
            .O(N__47386),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ));
    CascadeMux I__11201 (
            .O(N__47381),
            .I(N__47377));
    InMux I__11200 (
            .O(N__47380),
            .I(N__47372));
    InMux I__11199 (
            .O(N__47377),
            .I(N__47372));
    LocalMux I__11198 (
            .O(N__47372),
            .I(N__47368));
    InMux I__11197 (
            .O(N__47371),
            .I(N__47365));
    Span4Mux_h I__11196 (
            .O(N__47368),
            .I(N__47362));
    LocalMux I__11195 (
            .O(N__47365),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ));
    Odrv4 I__11194 (
            .O(N__47362),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ));
    InMux I__11193 (
            .O(N__47357),
            .I(N__47354));
    LocalMux I__11192 (
            .O(N__47354),
            .I(N__47351));
    Odrv4 I__11191 (
            .O(N__47351),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ));
    InMux I__11190 (
            .O(N__47348),
            .I(N__47343));
    InMux I__11189 (
            .O(N__47347),
            .I(N__47340));
    InMux I__11188 (
            .O(N__47346),
            .I(N__47337));
    LocalMux I__11187 (
            .O(N__47343),
            .I(N__47334));
    LocalMux I__11186 (
            .O(N__47340),
            .I(N__47331));
    LocalMux I__11185 (
            .O(N__47337),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    Odrv12 I__11184 (
            .O(N__47334),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    Odrv4 I__11183 (
            .O(N__47331),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    InMux I__11182 (
            .O(N__47324),
            .I(N__47320));
    InMux I__11181 (
            .O(N__47323),
            .I(N__47316));
    LocalMux I__11180 (
            .O(N__47320),
            .I(N__47313));
    InMux I__11179 (
            .O(N__47319),
            .I(N__47310));
    LocalMux I__11178 (
            .O(N__47316),
            .I(N__47307));
    Span4Mux_h I__11177 (
            .O(N__47313),
            .I(N__47304));
    LocalMux I__11176 (
            .O(N__47310),
            .I(N__47299));
    Span4Mux_h I__11175 (
            .O(N__47307),
            .I(N__47299));
    Span4Mux_h I__11174 (
            .O(N__47304),
            .I(N__47295));
    Span4Mux_h I__11173 (
            .O(N__47299),
            .I(N__47292));
    InMux I__11172 (
            .O(N__47298),
            .I(N__47289));
    Odrv4 I__11171 (
            .O(N__47295),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    Odrv4 I__11170 (
            .O(N__47292),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    LocalMux I__11169 (
            .O(N__47289),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    InMux I__11168 (
            .O(N__47282),
            .I(N__47276));
    InMux I__11167 (
            .O(N__47281),
            .I(N__47276));
    LocalMux I__11166 (
            .O(N__47276),
            .I(N__47273));
    Odrv12 I__11165 (
            .O(N__47273),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ));
    InMux I__11164 (
            .O(N__47270),
            .I(N__47266));
    InMux I__11163 (
            .O(N__47269),
            .I(N__47263));
    LocalMux I__11162 (
            .O(N__47266),
            .I(N__47260));
    LocalMux I__11161 (
            .O(N__47263),
            .I(N__47257));
    Sp12to4 I__11160 (
            .O(N__47260),
            .I(N__47254));
    Span4Mux_v I__11159 (
            .O(N__47257),
            .I(N__47251));
    Span12Mux_v I__11158 (
            .O(N__47254),
            .I(N__47248));
    Sp12to4 I__11157 (
            .O(N__47251),
            .I(N__47245));
    Odrv12 I__11156 (
            .O(N__47248),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    Odrv12 I__11155 (
            .O(N__47245),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    InMux I__11154 (
            .O(N__47240),
            .I(N__47237));
    LocalMux I__11153 (
            .O(N__47237),
            .I(N__47234));
    Odrv4 I__11152 (
            .O(N__47234),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ));
    InMux I__11151 (
            .O(N__47231),
            .I(N__47227));
    InMux I__11150 (
            .O(N__47230),
            .I(N__47223));
    LocalMux I__11149 (
            .O(N__47227),
            .I(N__47220));
    InMux I__11148 (
            .O(N__47226),
            .I(N__47217));
    LocalMux I__11147 (
            .O(N__47223),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    Odrv12 I__11146 (
            .O(N__47220),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    LocalMux I__11145 (
            .O(N__47217),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    InMux I__11144 (
            .O(N__47210),
            .I(N__47206));
    InMux I__11143 (
            .O(N__47209),
            .I(N__47202));
    LocalMux I__11142 (
            .O(N__47206),
            .I(N__47199));
    InMux I__11141 (
            .O(N__47205),
            .I(N__47196));
    LocalMux I__11140 (
            .O(N__47202),
            .I(N__47192));
    Span4Mux_h I__11139 (
            .O(N__47199),
            .I(N__47189));
    LocalMux I__11138 (
            .O(N__47196),
            .I(N__47186));
    CascadeMux I__11137 (
            .O(N__47195),
            .I(N__47183));
    Span4Mux_v I__11136 (
            .O(N__47192),
            .I(N__47178));
    Span4Mux_h I__11135 (
            .O(N__47189),
            .I(N__47178));
    Span12Mux_v I__11134 (
            .O(N__47186),
            .I(N__47175));
    InMux I__11133 (
            .O(N__47183),
            .I(N__47172));
    Odrv4 I__11132 (
            .O(N__47178),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    Odrv12 I__11131 (
            .O(N__47175),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    LocalMux I__11130 (
            .O(N__47172),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__11129 (
            .O(N__47165),
            .I(N__47157));
    InMux I__11128 (
            .O(N__47164),
            .I(N__47154));
    InMux I__11127 (
            .O(N__47163),
            .I(N__47151));
    InMux I__11126 (
            .O(N__47162),
            .I(N__47148));
    InMux I__11125 (
            .O(N__47161),
            .I(N__47125));
    InMux I__11124 (
            .O(N__47160),
            .I(N__47125));
    LocalMux I__11123 (
            .O(N__47157),
            .I(N__47103));
    LocalMux I__11122 (
            .O(N__47154),
            .I(N__47096));
    LocalMux I__11121 (
            .O(N__47151),
            .I(N__47096));
    LocalMux I__11120 (
            .O(N__47148),
            .I(N__47096));
    InMux I__11119 (
            .O(N__47147),
            .I(N__47091));
    InMux I__11118 (
            .O(N__47146),
            .I(N__47091));
    CascadeMux I__11117 (
            .O(N__47145),
            .I(N__47085));
    InMux I__11116 (
            .O(N__47144),
            .I(N__47072));
    InMux I__11115 (
            .O(N__47143),
            .I(N__47072));
    InMux I__11114 (
            .O(N__47142),
            .I(N__47072));
    InMux I__11113 (
            .O(N__47141),
            .I(N__47072));
    InMux I__11112 (
            .O(N__47140),
            .I(N__47067));
    InMux I__11111 (
            .O(N__47139),
            .I(N__47067));
    InMux I__11110 (
            .O(N__47138),
            .I(N__47048));
    InMux I__11109 (
            .O(N__47137),
            .I(N__47045));
    InMux I__11108 (
            .O(N__47136),
            .I(N__47034));
    InMux I__11107 (
            .O(N__47135),
            .I(N__47034));
    InMux I__11106 (
            .O(N__47134),
            .I(N__47034));
    InMux I__11105 (
            .O(N__47133),
            .I(N__47034));
    InMux I__11104 (
            .O(N__47132),
            .I(N__47034));
    InMux I__11103 (
            .O(N__47131),
            .I(N__47029));
    InMux I__11102 (
            .O(N__47130),
            .I(N__47029));
    LocalMux I__11101 (
            .O(N__47125),
            .I(N__47026));
    InMux I__11100 (
            .O(N__47124),
            .I(N__47021));
    InMux I__11099 (
            .O(N__47123),
            .I(N__47021));
    InMux I__11098 (
            .O(N__47122),
            .I(N__47018));
    InMux I__11097 (
            .O(N__47121),
            .I(N__47013));
    InMux I__11096 (
            .O(N__47120),
            .I(N__47013));
    InMux I__11095 (
            .O(N__47119),
            .I(N__47004));
    InMux I__11094 (
            .O(N__47118),
            .I(N__47004));
    InMux I__11093 (
            .O(N__47117),
            .I(N__47004));
    InMux I__11092 (
            .O(N__47116),
            .I(N__47004));
    InMux I__11091 (
            .O(N__47115),
            .I(N__46995));
    InMux I__11090 (
            .O(N__47114),
            .I(N__46995));
    InMux I__11089 (
            .O(N__47113),
            .I(N__46995));
    InMux I__11088 (
            .O(N__47112),
            .I(N__46995));
    InMux I__11087 (
            .O(N__47111),
            .I(N__46985));
    InMux I__11086 (
            .O(N__47110),
            .I(N__46985));
    InMux I__11085 (
            .O(N__47109),
            .I(N__46978));
    InMux I__11084 (
            .O(N__47108),
            .I(N__46978));
    InMux I__11083 (
            .O(N__47107),
            .I(N__46978));
    InMux I__11082 (
            .O(N__47106),
            .I(N__46971));
    Span4Mux_v I__11081 (
            .O(N__47103),
            .I(N__46964));
    Span4Mux_v I__11080 (
            .O(N__47096),
            .I(N__46964));
    LocalMux I__11079 (
            .O(N__47091),
            .I(N__46964));
    InMux I__11078 (
            .O(N__47090),
            .I(N__46957));
    InMux I__11077 (
            .O(N__47089),
            .I(N__46957));
    InMux I__11076 (
            .O(N__47088),
            .I(N__46957));
    InMux I__11075 (
            .O(N__47085),
            .I(N__46954));
    InMux I__11074 (
            .O(N__47084),
            .I(N__46949));
    InMux I__11073 (
            .O(N__47083),
            .I(N__46949));
    InMux I__11072 (
            .O(N__47082),
            .I(N__46946));
    InMux I__11071 (
            .O(N__47081),
            .I(N__46943));
    LocalMux I__11070 (
            .O(N__47072),
            .I(N__46940));
    LocalMux I__11069 (
            .O(N__47067),
            .I(N__46937));
    InMux I__11068 (
            .O(N__47066),
            .I(N__46916));
    InMux I__11067 (
            .O(N__47065),
            .I(N__46916));
    InMux I__11066 (
            .O(N__47064),
            .I(N__46907));
    InMux I__11065 (
            .O(N__47063),
            .I(N__46907));
    InMux I__11064 (
            .O(N__47062),
            .I(N__46907));
    InMux I__11063 (
            .O(N__47061),
            .I(N__46907));
    InMux I__11062 (
            .O(N__47060),
            .I(N__46900));
    InMux I__11061 (
            .O(N__47059),
            .I(N__46900));
    InMux I__11060 (
            .O(N__47058),
            .I(N__46900));
    InMux I__11059 (
            .O(N__47057),
            .I(N__46893));
    InMux I__11058 (
            .O(N__47056),
            .I(N__46893));
    InMux I__11057 (
            .O(N__47055),
            .I(N__46893));
    InMux I__11056 (
            .O(N__47054),
            .I(N__46884));
    InMux I__11055 (
            .O(N__47053),
            .I(N__46884));
    InMux I__11054 (
            .O(N__47052),
            .I(N__46884));
    InMux I__11053 (
            .O(N__47051),
            .I(N__46884));
    LocalMux I__11052 (
            .O(N__47048),
            .I(N__46877));
    LocalMux I__11051 (
            .O(N__47045),
            .I(N__46877));
    LocalMux I__11050 (
            .O(N__47034),
            .I(N__46877));
    LocalMux I__11049 (
            .O(N__47029),
            .I(N__46870));
    Span4Mux_v I__11048 (
            .O(N__47026),
            .I(N__46870));
    LocalMux I__11047 (
            .O(N__47021),
            .I(N__46870));
    LocalMux I__11046 (
            .O(N__47018),
            .I(N__46861));
    LocalMux I__11045 (
            .O(N__47013),
            .I(N__46861));
    LocalMux I__11044 (
            .O(N__47004),
            .I(N__46861));
    LocalMux I__11043 (
            .O(N__46995),
            .I(N__46861));
    InMux I__11042 (
            .O(N__46994),
            .I(N__46850));
    InMux I__11041 (
            .O(N__46993),
            .I(N__46850));
    InMux I__11040 (
            .O(N__46992),
            .I(N__46850));
    InMux I__11039 (
            .O(N__46991),
            .I(N__46850));
    InMux I__11038 (
            .O(N__46990),
            .I(N__46850));
    LocalMux I__11037 (
            .O(N__46985),
            .I(N__46845));
    LocalMux I__11036 (
            .O(N__46978),
            .I(N__46845));
    InMux I__11035 (
            .O(N__46977),
            .I(N__46842));
    InMux I__11034 (
            .O(N__46976),
            .I(N__46834));
    InMux I__11033 (
            .O(N__46975),
            .I(N__46834));
    InMux I__11032 (
            .O(N__46974),
            .I(N__46834));
    LocalMux I__11031 (
            .O(N__46971),
            .I(N__46823));
    Span4Mux_h I__11030 (
            .O(N__46964),
            .I(N__46823));
    LocalMux I__11029 (
            .O(N__46957),
            .I(N__46823));
    LocalMux I__11028 (
            .O(N__46954),
            .I(N__46823));
    LocalMux I__11027 (
            .O(N__46949),
            .I(N__46823));
    LocalMux I__11026 (
            .O(N__46946),
            .I(N__46814));
    LocalMux I__11025 (
            .O(N__46943),
            .I(N__46814));
    Span4Mux_h I__11024 (
            .O(N__46940),
            .I(N__46814));
    Span4Mux_h I__11023 (
            .O(N__46937),
            .I(N__46814));
    InMux I__11022 (
            .O(N__46936),
            .I(N__46811));
    InMux I__11021 (
            .O(N__46935),
            .I(N__46808));
    InMux I__11020 (
            .O(N__46934),
            .I(N__46801));
    InMux I__11019 (
            .O(N__46933),
            .I(N__46801));
    InMux I__11018 (
            .O(N__46932),
            .I(N__46801));
    InMux I__11017 (
            .O(N__46931),
            .I(N__46796));
    InMux I__11016 (
            .O(N__46930),
            .I(N__46796));
    InMux I__11015 (
            .O(N__46929),
            .I(N__46785));
    InMux I__11014 (
            .O(N__46928),
            .I(N__46785));
    InMux I__11013 (
            .O(N__46927),
            .I(N__46785));
    InMux I__11012 (
            .O(N__46926),
            .I(N__46785));
    InMux I__11011 (
            .O(N__46925),
            .I(N__46785));
    InMux I__11010 (
            .O(N__46924),
            .I(N__46776));
    InMux I__11009 (
            .O(N__46923),
            .I(N__46776));
    InMux I__11008 (
            .O(N__46922),
            .I(N__46776));
    InMux I__11007 (
            .O(N__46921),
            .I(N__46776));
    LocalMux I__11006 (
            .O(N__46916),
            .I(N__46773));
    LocalMux I__11005 (
            .O(N__46907),
            .I(N__46764));
    LocalMux I__11004 (
            .O(N__46900),
            .I(N__46764));
    LocalMux I__11003 (
            .O(N__46893),
            .I(N__46764));
    LocalMux I__11002 (
            .O(N__46884),
            .I(N__46764));
    Span4Mux_v I__11001 (
            .O(N__46877),
            .I(N__46757));
    Span4Mux_v I__11000 (
            .O(N__46870),
            .I(N__46757));
    Span4Mux_v I__10999 (
            .O(N__46861),
            .I(N__46757));
    LocalMux I__10998 (
            .O(N__46850),
            .I(N__46750));
    Span12Mux_v I__10997 (
            .O(N__46845),
            .I(N__46750));
    LocalMux I__10996 (
            .O(N__46842),
            .I(N__46750));
    InMux I__10995 (
            .O(N__46841),
            .I(N__46747));
    LocalMux I__10994 (
            .O(N__46834),
            .I(N__46740));
    Span4Mux_v I__10993 (
            .O(N__46823),
            .I(N__46740));
    Span4Mux_v I__10992 (
            .O(N__46814),
            .I(N__46740));
    LocalMux I__10991 (
            .O(N__46811),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__10990 (
            .O(N__46808),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__10989 (
            .O(N__46801),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__10988 (
            .O(N__46796),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__10987 (
            .O(N__46785),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__10986 (
            .O(N__46776),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__10985 (
            .O(N__46773),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__10984 (
            .O(N__46764),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__10983 (
            .O(N__46757),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv12 I__10982 (
            .O(N__46750),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__10981 (
            .O(N__46747),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__10980 (
            .O(N__46740),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    InMux I__10979 (
            .O(N__46715),
            .I(N__46709));
    InMux I__10978 (
            .O(N__46714),
            .I(N__46709));
    LocalMux I__10977 (
            .O(N__46709),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ));
    CEMux I__10976 (
            .O(N__46706),
            .I(N__46703));
    LocalMux I__10975 (
            .O(N__46703),
            .I(N__46691));
    CEMux I__10974 (
            .O(N__46702),
            .I(N__46688));
    InMux I__10973 (
            .O(N__46701),
            .I(N__46672));
    CEMux I__10972 (
            .O(N__46700),
            .I(N__46669));
    CEMux I__10971 (
            .O(N__46699),
            .I(N__46666));
    CEMux I__10970 (
            .O(N__46698),
            .I(N__46658));
    InMux I__10969 (
            .O(N__46697),
            .I(N__46648));
    InMux I__10968 (
            .O(N__46696),
            .I(N__46648));
    InMux I__10967 (
            .O(N__46695),
            .I(N__46648));
    InMux I__10966 (
            .O(N__46694),
            .I(N__46648));
    Span4Mux_v I__10965 (
            .O(N__46691),
            .I(N__46643));
    LocalMux I__10964 (
            .O(N__46688),
            .I(N__46643));
    CEMux I__10963 (
            .O(N__46687),
            .I(N__46640));
    CEMux I__10962 (
            .O(N__46686),
            .I(N__46637));
    InMux I__10961 (
            .O(N__46685),
            .I(N__46628));
    InMux I__10960 (
            .O(N__46684),
            .I(N__46628));
    InMux I__10959 (
            .O(N__46683),
            .I(N__46628));
    InMux I__10958 (
            .O(N__46682),
            .I(N__46628));
    InMux I__10957 (
            .O(N__46681),
            .I(N__46619));
    InMux I__10956 (
            .O(N__46680),
            .I(N__46619));
    InMux I__10955 (
            .O(N__46679),
            .I(N__46619));
    InMux I__10954 (
            .O(N__46678),
            .I(N__46619));
    CEMux I__10953 (
            .O(N__46677),
            .I(N__46616));
    CEMux I__10952 (
            .O(N__46676),
            .I(N__46611));
    CEMux I__10951 (
            .O(N__46675),
            .I(N__46598));
    LocalMux I__10950 (
            .O(N__46672),
            .I(N__46595));
    LocalMux I__10949 (
            .O(N__46669),
            .I(N__46586));
    LocalMux I__10948 (
            .O(N__46666),
            .I(N__46583));
    CEMux I__10947 (
            .O(N__46665),
            .I(N__46580));
    InMux I__10946 (
            .O(N__46664),
            .I(N__46571));
    InMux I__10945 (
            .O(N__46663),
            .I(N__46571));
    InMux I__10944 (
            .O(N__46662),
            .I(N__46571));
    InMux I__10943 (
            .O(N__46661),
            .I(N__46571));
    LocalMux I__10942 (
            .O(N__46658),
            .I(N__46568));
    CEMux I__10941 (
            .O(N__46657),
            .I(N__46565));
    LocalMux I__10940 (
            .O(N__46648),
            .I(N__46562));
    Span4Mux_h I__10939 (
            .O(N__46643),
            .I(N__46557));
    LocalMux I__10938 (
            .O(N__46640),
            .I(N__46557));
    LocalMux I__10937 (
            .O(N__46637),
            .I(N__46554));
    LocalMux I__10936 (
            .O(N__46628),
            .I(N__46547));
    LocalMux I__10935 (
            .O(N__46619),
            .I(N__46547));
    LocalMux I__10934 (
            .O(N__46616),
            .I(N__46547));
    CEMux I__10933 (
            .O(N__46615),
            .I(N__46544));
    CEMux I__10932 (
            .O(N__46614),
            .I(N__46541));
    LocalMux I__10931 (
            .O(N__46611),
            .I(N__46538));
    InMux I__10930 (
            .O(N__46610),
            .I(N__46531));
    InMux I__10929 (
            .O(N__46609),
            .I(N__46531));
    InMux I__10928 (
            .O(N__46608),
            .I(N__46531));
    InMux I__10927 (
            .O(N__46607),
            .I(N__46522));
    InMux I__10926 (
            .O(N__46606),
            .I(N__46522));
    InMux I__10925 (
            .O(N__46605),
            .I(N__46522));
    InMux I__10924 (
            .O(N__46604),
            .I(N__46522));
    InMux I__10923 (
            .O(N__46603),
            .I(N__46515));
    InMux I__10922 (
            .O(N__46602),
            .I(N__46515));
    InMux I__10921 (
            .O(N__46601),
            .I(N__46515));
    LocalMux I__10920 (
            .O(N__46598),
            .I(N__46512));
    Span4Mux_h I__10919 (
            .O(N__46595),
            .I(N__46509));
    InMux I__10918 (
            .O(N__46594),
            .I(N__46500));
    InMux I__10917 (
            .O(N__46593),
            .I(N__46500));
    InMux I__10916 (
            .O(N__46592),
            .I(N__46500));
    InMux I__10915 (
            .O(N__46591),
            .I(N__46500));
    CEMux I__10914 (
            .O(N__46590),
            .I(N__46497));
    CEMux I__10913 (
            .O(N__46589),
            .I(N__46494));
    Span4Mux_h I__10912 (
            .O(N__46586),
            .I(N__46477));
    Span4Mux_h I__10911 (
            .O(N__46583),
            .I(N__46477));
    LocalMux I__10910 (
            .O(N__46580),
            .I(N__46477));
    LocalMux I__10909 (
            .O(N__46571),
            .I(N__46477));
    Span4Mux_v I__10908 (
            .O(N__46568),
            .I(N__46477));
    LocalMux I__10907 (
            .O(N__46565),
            .I(N__46477));
    Span4Mux_h I__10906 (
            .O(N__46562),
            .I(N__46477));
    Span4Mux_v I__10905 (
            .O(N__46557),
            .I(N__46477));
    Span4Mux_v I__10904 (
            .O(N__46554),
            .I(N__46474));
    Span4Mux_h I__10903 (
            .O(N__46547),
            .I(N__46471));
    LocalMux I__10902 (
            .O(N__46544),
            .I(N__46468));
    LocalMux I__10901 (
            .O(N__46541),
            .I(N__46465));
    Span4Mux_v I__10900 (
            .O(N__46538),
            .I(N__46454));
    LocalMux I__10899 (
            .O(N__46531),
            .I(N__46454));
    LocalMux I__10898 (
            .O(N__46522),
            .I(N__46454));
    LocalMux I__10897 (
            .O(N__46515),
            .I(N__46454));
    Span4Mux_h I__10896 (
            .O(N__46512),
            .I(N__46454));
    Span4Mux_v I__10895 (
            .O(N__46509),
            .I(N__46451));
    LocalMux I__10894 (
            .O(N__46500),
            .I(N__46448));
    LocalMux I__10893 (
            .O(N__46497),
            .I(N__46439));
    LocalMux I__10892 (
            .O(N__46494),
            .I(N__46439));
    Span4Mux_v I__10891 (
            .O(N__46477),
            .I(N__46439));
    Span4Mux_s3_h I__10890 (
            .O(N__46474),
            .I(N__46439));
    Span4Mux_v I__10889 (
            .O(N__46471),
            .I(N__46436));
    Span4Mux_h I__10888 (
            .O(N__46468),
            .I(N__46427));
    Span4Mux_h I__10887 (
            .O(N__46465),
            .I(N__46427));
    Span4Mux_v I__10886 (
            .O(N__46454),
            .I(N__46427));
    Span4Mux_h I__10885 (
            .O(N__46451),
            .I(N__46427));
    Span4Mux_v I__10884 (
            .O(N__46448),
            .I(N__46422));
    Span4Mux_h I__10883 (
            .O(N__46439),
            .I(N__46422));
    Odrv4 I__10882 (
            .O(N__46436),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__10881 (
            .O(N__46427),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__10880 (
            .O(N__46422),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    CascadeMux I__10879 (
            .O(N__46415),
            .I(N__46410));
    CascadeMux I__10878 (
            .O(N__46414),
            .I(N__46407));
    InMux I__10877 (
            .O(N__46413),
            .I(N__46400));
    InMux I__10876 (
            .O(N__46410),
            .I(N__46400));
    InMux I__10875 (
            .O(N__46407),
            .I(N__46400));
    LocalMux I__10874 (
            .O(N__46400),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ));
    InMux I__10873 (
            .O(N__46397),
            .I(N__46391));
    InMux I__10872 (
            .O(N__46396),
            .I(N__46388));
    InMux I__10871 (
            .O(N__46395),
            .I(N__46385));
    InMux I__10870 (
            .O(N__46394),
            .I(N__46382));
    LocalMux I__10869 (
            .O(N__46391),
            .I(N__46379));
    LocalMux I__10868 (
            .O(N__46388),
            .I(N__46374));
    LocalMux I__10867 (
            .O(N__46385),
            .I(N__46374));
    LocalMux I__10866 (
            .O(N__46382),
            .I(N__46371));
    Span4Mux_h I__10865 (
            .O(N__46379),
            .I(N__46368));
    Span4Mux_h I__10864 (
            .O(N__46374),
            .I(N__46365));
    Span4Mux_v I__10863 (
            .O(N__46371),
            .I(N__46362));
    Odrv4 I__10862 (
            .O(N__46368),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    Odrv4 I__10861 (
            .O(N__46365),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    Odrv4 I__10860 (
            .O(N__46362),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    InMux I__10859 (
            .O(N__46355),
            .I(N__46350));
    InMux I__10858 (
            .O(N__46354),
            .I(N__46347));
    InMux I__10857 (
            .O(N__46353),
            .I(N__46344));
    LocalMux I__10856 (
            .O(N__46350),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    LocalMux I__10855 (
            .O(N__46347),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    LocalMux I__10854 (
            .O(N__46344),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    InMux I__10853 (
            .O(N__46337),
            .I(N__46332));
    InMux I__10852 (
            .O(N__46336),
            .I(N__46329));
    InMux I__10851 (
            .O(N__46335),
            .I(N__46326));
    LocalMux I__10850 (
            .O(N__46332),
            .I(N__46323));
    LocalMux I__10849 (
            .O(N__46329),
            .I(N__46320));
    LocalMux I__10848 (
            .O(N__46326),
            .I(N__46316));
    Span4Mux_h I__10847 (
            .O(N__46323),
            .I(N__46313));
    Span4Mux_h I__10846 (
            .O(N__46320),
            .I(N__46310));
    InMux I__10845 (
            .O(N__46319),
            .I(N__46307));
    Odrv4 I__10844 (
            .O(N__46316),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    Odrv4 I__10843 (
            .O(N__46313),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    Odrv4 I__10842 (
            .O(N__46310),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    LocalMux I__10841 (
            .O(N__46307),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    InMux I__10840 (
            .O(N__46298),
            .I(N__46295));
    LocalMux I__10839 (
            .O(N__46295),
            .I(N__46292));
    Span4Mux_h I__10838 (
            .O(N__46292),
            .I(N__46288));
    InMux I__10837 (
            .O(N__46291),
            .I(N__46284));
    Span4Mux_h I__10836 (
            .O(N__46288),
            .I(N__46281));
    InMux I__10835 (
            .O(N__46287),
            .I(N__46278));
    LocalMux I__10834 (
            .O(N__46284),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    Odrv4 I__10833 (
            .O(N__46281),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    LocalMux I__10832 (
            .O(N__46278),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    InMux I__10831 (
            .O(N__46271),
            .I(N__46268));
    LocalMux I__10830 (
            .O(N__46268),
            .I(N__46264));
    InMux I__10829 (
            .O(N__46267),
            .I(N__46261));
    Sp12to4 I__10828 (
            .O(N__46264),
            .I(N__46256));
    LocalMux I__10827 (
            .O(N__46261),
            .I(N__46256));
    Odrv12 I__10826 (
            .O(N__46256),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ));
    CascadeMux I__10825 (
            .O(N__46253),
            .I(N__46250));
    InMux I__10824 (
            .O(N__46250),
            .I(N__46247));
    LocalMux I__10823 (
            .O(N__46247),
            .I(N__46243));
    InMux I__10822 (
            .O(N__46246),
            .I(N__46239));
    Span4Mux_v I__10821 (
            .O(N__46243),
            .I(N__46235));
    InMux I__10820 (
            .O(N__46242),
            .I(N__46232));
    LocalMux I__10819 (
            .O(N__46239),
            .I(N__46229));
    InMux I__10818 (
            .O(N__46238),
            .I(N__46225));
    Span4Mux_v I__10817 (
            .O(N__46235),
            .I(N__46222));
    LocalMux I__10816 (
            .O(N__46232),
            .I(N__46219));
    Span4Mux_v I__10815 (
            .O(N__46229),
            .I(N__46216));
    InMux I__10814 (
            .O(N__46228),
            .I(N__46213));
    LocalMux I__10813 (
            .O(N__46225),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    Odrv4 I__10812 (
            .O(N__46222),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    Odrv12 I__10811 (
            .O(N__46219),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    Odrv4 I__10810 (
            .O(N__46216),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    LocalMux I__10809 (
            .O(N__46213),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    InMux I__10808 (
            .O(N__46202),
            .I(N__46198));
    InMux I__10807 (
            .O(N__46201),
            .I(N__46195));
    LocalMux I__10806 (
            .O(N__46198),
            .I(N__46192));
    LocalMux I__10805 (
            .O(N__46195),
            .I(N__46186));
    Span4Mux_h I__10804 (
            .O(N__46192),
            .I(N__46183));
    InMux I__10803 (
            .O(N__46191),
            .I(N__46178));
    InMux I__10802 (
            .O(N__46190),
            .I(N__46178));
    InMux I__10801 (
            .O(N__46189),
            .I(N__46175));
    Span12Mux_s9_h I__10800 (
            .O(N__46186),
            .I(N__46168));
    Sp12to4 I__10799 (
            .O(N__46183),
            .I(N__46168));
    LocalMux I__10798 (
            .O(N__46178),
            .I(N__46168));
    LocalMux I__10797 (
            .O(N__46175),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    Odrv12 I__10796 (
            .O(N__46168),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    InMux I__10795 (
            .O(N__46163),
            .I(N__46160));
    LocalMux I__10794 (
            .O(N__46160),
            .I(N__46156));
    InMux I__10793 (
            .O(N__46159),
            .I(N__46153));
    Span4Mux_v I__10792 (
            .O(N__46156),
            .I(N__46150));
    LocalMux I__10791 (
            .O(N__46153),
            .I(N__46146));
    Span4Mux_v I__10790 (
            .O(N__46150),
            .I(N__46143));
    InMux I__10789 (
            .O(N__46149),
            .I(N__46140));
    Span4Mux_v I__10788 (
            .O(N__46146),
            .I(N__46137));
    Odrv4 I__10787 (
            .O(N__46143),
            .I(\phase_controller_inst1.tr_time_passed ));
    LocalMux I__10786 (
            .O(N__46140),
            .I(\phase_controller_inst1.tr_time_passed ));
    Odrv4 I__10785 (
            .O(N__46137),
            .I(\phase_controller_inst1.tr_time_passed ));
    InMux I__10784 (
            .O(N__46130),
            .I(N__46124));
    InMux I__10783 (
            .O(N__46129),
            .I(N__46124));
    LocalMux I__10782 (
            .O(N__46124),
            .I(N__46121));
    Odrv12 I__10781 (
            .O(N__46121),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ));
    CEMux I__10780 (
            .O(N__46118),
            .I(N__46082));
    CEMux I__10779 (
            .O(N__46117),
            .I(N__46082));
    CEMux I__10778 (
            .O(N__46116),
            .I(N__46082));
    CEMux I__10777 (
            .O(N__46115),
            .I(N__46082));
    CEMux I__10776 (
            .O(N__46114),
            .I(N__46082));
    CEMux I__10775 (
            .O(N__46113),
            .I(N__46082));
    CEMux I__10774 (
            .O(N__46112),
            .I(N__46082));
    CEMux I__10773 (
            .O(N__46111),
            .I(N__46082));
    CEMux I__10772 (
            .O(N__46110),
            .I(N__46082));
    CEMux I__10771 (
            .O(N__46109),
            .I(N__46082));
    CEMux I__10770 (
            .O(N__46108),
            .I(N__46082));
    CEMux I__10769 (
            .O(N__46107),
            .I(N__46082));
    GlobalMux I__10768 (
            .O(N__46082),
            .I(N__46079));
    gio2CtrlBuf I__10767 (
            .O(N__46079),
            .I(\phase_controller_inst2.stoper_tr.un1_start_g ));
    InMux I__10766 (
            .O(N__46076),
            .I(N__46072));
    InMux I__10765 (
            .O(N__46075),
            .I(N__46069));
    LocalMux I__10764 (
            .O(N__46072),
            .I(N__46065));
    LocalMux I__10763 (
            .O(N__46069),
            .I(N__46062));
    InMux I__10762 (
            .O(N__46068),
            .I(N__46059));
    Span4Mux_h I__10761 (
            .O(N__46065),
            .I(N__46056));
    Span4Mux_h I__10760 (
            .O(N__46062),
            .I(N__46053));
    LocalMux I__10759 (
            .O(N__46059),
            .I(N__46048));
    Span4Mux_v I__10758 (
            .O(N__46056),
            .I(N__46048));
    Span4Mux_v I__10757 (
            .O(N__46053),
            .I(N__46045));
    Span4Mux_h I__10756 (
            .O(N__46048),
            .I(N__46041));
    Span4Mux_h I__10755 (
            .O(N__46045),
            .I(N__46038));
    InMux I__10754 (
            .O(N__46044),
            .I(N__46035));
    Odrv4 I__10753 (
            .O(N__46041),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    Odrv4 I__10752 (
            .O(N__46038),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    LocalMux I__10751 (
            .O(N__46035),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__10750 (
            .O(N__46028),
            .I(N__46025));
    LocalMux I__10749 (
            .O(N__46025),
            .I(N__46021));
    InMux I__10748 (
            .O(N__46024),
            .I(N__46017));
    Span4Mux_h I__10747 (
            .O(N__46021),
            .I(N__46014));
    InMux I__10746 (
            .O(N__46020),
            .I(N__46011));
    LocalMux I__10745 (
            .O(N__46017),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    Odrv4 I__10744 (
            .O(N__46014),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    LocalMux I__10743 (
            .O(N__46011),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    InMux I__10742 (
            .O(N__46004),
            .I(N__46001));
    LocalMux I__10741 (
            .O(N__46001),
            .I(N__45997));
    InMux I__10740 (
            .O(N__46000),
            .I(N__45993));
    Span4Mux_h I__10739 (
            .O(N__45997),
            .I(N__45990));
    InMux I__10738 (
            .O(N__45996),
            .I(N__45987));
    LocalMux I__10737 (
            .O(N__45993),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    Odrv4 I__10736 (
            .O(N__45990),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    LocalMux I__10735 (
            .O(N__45987),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    InMux I__10734 (
            .O(N__45980),
            .I(N__45977));
    LocalMux I__10733 (
            .O(N__45977),
            .I(N__45971));
    InMux I__10732 (
            .O(N__45976),
            .I(N__45968));
    InMux I__10731 (
            .O(N__45975),
            .I(N__45965));
    InMux I__10730 (
            .O(N__45974),
            .I(N__45962));
    Span4Mux_h I__10729 (
            .O(N__45971),
            .I(N__45957));
    LocalMux I__10728 (
            .O(N__45968),
            .I(N__45957));
    LocalMux I__10727 (
            .O(N__45965),
            .I(N__45954));
    LocalMux I__10726 (
            .O(N__45962),
            .I(N__45949));
    Span4Mux_h I__10725 (
            .O(N__45957),
            .I(N__45949));
    Odrv4 I__10724 (
            .O(N__45954),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    Odrv4 I__10723 (
            .O(N__45949),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    CascadeMux I__10722 (
            .O(N__45944),
            .I(N__45941));
    InMux I__10721 (
            .O(N__45941),
            .I(N__45938));
    LocalMux I__10720 (
            .O(N__45938),
            .I(N__45935));
    Odrv4 I__10719 (
            .O(N__45935),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ));
    CascadeMux I__10718 (
            .O(N__45932),
            .I(N__45929));
    InMux I__10717 (
            .O(N__45929),
            .I(N__45926));
    LocalMux I__10716 (
            .O(N__45926),
            .I(N__45923));
    Odrv12 I__10715 (
            .O(N__45923),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt22 ));
    InMux I__10714 (
            .O(N__45920),
            .I(N__45914));
    InMux I__10713 (
            .O(N__45919),
            .I(N__45914));
    LocalMux I__10712 (
            .O(N__45914),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ));
    InMux I__10711 (
            .O(N__45911),
            .I(N__45908));
    LocalMux I__10710 (
            .O(N__45908),
            .I(N__45904));
    InMux I__10709 (
            .O(N__45907),
            .I(N__45901));
    Odrv4 I__10708 (
            .O(N__45904),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ));
    LocalMux I__10707 (
            .O(N__45901),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ));
    InMux I__10706 (
            .O(N__45896),
            .I(N__45892));
    InMux I__10705 (
            .O(N__45895),
            .I(N__45888));
    LocalMux I__10704 (
            .O(N__45892),
            .I(N__45885));
    InMux I__10703 (
            .O(N__45891),
            .I(N__45882));
    LocalMux I__10702 (
            .O(N__45888),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    Odrv4 I__10701 (
            .O(N__45885),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    LocalMux I__10700 (
            .O(N__45882),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    CascadeMux I__10699 (
            .O(N__45875),
            .I(N__45870));
    CascadeMux I__10698 (
            .O(N__45874),
            .I(N__45867));
    InMux I__10697 (
            .O(N__45873),
            .I(N__45864));
    InMux I__10696 (
            .O(N__45870),
            .I(N__45861));
    InMux I__10695 (
            .O(N__45867),
            .I(N__45858));
    LocalMux I__10694 (
            .O(N__45864),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    LocalMux I__10693 (
            .O(N__45861),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    LocalMux I__10692 (
            .O(N__45858),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    InMux I__10691 (
            .O(N__45851),
            .I(N__45847));
    InMux I__10690 (
            .O(N__45850),
            .I(N__45844));
    LocalMux I__10689 (
            .O(N__45847),
            .I(N__45841));
    LocalMux I__10688 (
            .O(N__45844),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ));
    Odrv4 I__10687 (
            .O(N__45841),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ));
    InMux I__10686 (
            .O(N__45836),
            .I(N__45833));
    LocalMux I__10685 (
            .O(N__45833),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ));
    CascadeMux I__10684 (
            .O(N__45830),
            .I(N__45826));
    InMux I__10683 (
            .O(N__45829),
            .I(N__45823));
    InMux I__10682 (
            .O(N__45826),
            .I(N__45820));
    LocalMux I__10681 (
            .O(N__45823),
            .I(N__45817));
    LocalMux I__10680 (
            .O(N__45820),
            .I(N__45814));
    Span4Mux_h I__10679 (
            .O(N__45817),
            .I(N__45811));
    Odrv4 I__10678 (
            .O(N__45814),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt30 ));
    Odrv4 I__10677 (
            .O(N__45811),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt30 ));
    InMux I__10676 (
            .O(N__45806),
            .I(N__45803));
    LocalMux I__10675 (
            .O(N__45803),
            .I(N__45799));
    InMux I__10674 (
            .O(N__45802),
            .I(N__45796));
    Odrv12 I__10673 (
            .O(N__45799),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    LocalMux I__10672 (
            .O(N__45796),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    CascadeMux I__10671 (
            .O(N__45791),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30_cascade_));
    InMux I__10670 (
            .O(N__45788),
            .I(N__45782));
    InMux I__10669 (
            .O(N__45787),
            .I(N__45777));
    InMux I__10668 (
            .O(N__45786),
            .I(N__45777));
    CascadeMux I__10667 (
            .O(N__45785),
            .I(N__45774));
    LocalMux I__10666 (
            .O(N__45782),
            .I(N__45771));
    LocalMux I__10665 (
            .O(N__45777),
            .I(N__45768));
    InMux I__10664 (
            .O(N__45774),
            .I(N__45765));
    Span4Mux_h I__10663 (
            .O(N__45771),
            .I(N__45758));
    Span4Mux_h I__10662 (
            .O(N__45768),
            .I(N__45758));
    LocalMux I__10661 (
            .O(N__45765),
            .I(N__45758));
    Odrv4 I__10660 (
            .O(N__45758),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    InMux I__10659 (
            .O(N__45755),
            .I(N__45752));
    LocalMux I__10658 (
            .O(N__45752),
            .I(N__45749));
    Odrv4 I__10657 (
            .O(N__45749),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30 ));
    InMux I__10656 (
            .O(N__45746),
            .I(N__45737));
    InMux I__10655 (
            .O(N__45745),
            .I(N__45737));
    InMux I__10654 (
            .O(N__45744),
            .I(N__45737));
    LocalMux I__10653 (
            .O(N__45737),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ));
    CascadeMux I__10652 (
            .O(N__45734),
            .I(N__45730));
    InMux I__10651 (
            .O(N__45733),
            .I(N__45725));
    InMux I__10650 (
            .O(N__45730),
            .I(N__45718));
    InMux I__10649 (
            .O(N__45729),
            .I(N__45718));
    InMux I__10648 (
            .O(N__45728),
            .I(N__45718));
    LocalMux I__10647 (
            .O(N__45725),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    LocalMux I__10646 (
            .O(N__45718),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    InMux I__10645 (
            .O(N__45713),
            .I(N__45707));
    InMux I__10644 (
            .O(N__45712),
            .I(N__45700));
    InMux I__10643 (
            .O(N__45711),
            .I(N__45700));
    InMux I__10642 (
            .O(N__45710),
            .I(N__45700));
    LocalMux I__10641 (
            .O(N__45707),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    LocalMux I__10640 (
            .O(N__45700),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    CascadeMux I__10639 (
            .O(N__45695),
            .I(N__45692));
    InMux I__10638 (
            .O(N__45692),
            .I(N__45689));
    LocalMux I__10637 (
            .O(N__45689),
            .I(N__45686));
    Span4Mux_h I__10636 (
            .O(N__45686),
            .I(N__45683));
    Odrv4 I__10635 (
            .O(N__45683),
            .I(\phase_controller_inst1.stoper_tr.un4_running_df30 ));
    InMux I__10634 (
            .O(N__45680),
            .I(N__45677));
    LocalMux I__10633 (
            .O(N__45677),
            .I(N__45674));
    Odrv12 I__10632 (
            .O(N__45674),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ));
    CascadeMux I__10631 (
            .O(N__45671),
            .I(N__45668));
    InMux I__10630 (
            .O(N__45668),
            .I(N__45665));
    LocalMux I__10629 (
            .O(N__45665),
            .I(N__45662));
    Span4Mux_h I__10628 (
            .O(N__45662),
            .I(N__45659));
    Odrv4 I__10627 (
            .O(N__45659),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt26 ));
    InMux I__10626 (
            .O(N__45656),
            .I(N__45653));
    LocalMux I__10625 (
            .O(N__45653),
            .I(N__45650));
    Odrv4 I__10624 (
            .O(N__45650),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ));
    CascadeMux I__10623 (
            .O(N__45647),
            .I(N__45644));
    InMux I__10622 (
            .O(N__45644),
            .I(N__45641));
    LocalMux I__10621 (
            .O(N__45641),
            .I(N__45638));
    Span4Mux_v I__10620 (
            .O(N__45638),
            .I(N__45635));
    Odrv4 I__10619 (
            .O(N__45635),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt28 ));
    InMux I__10618 (
            .O(N__45632),
            .I(N__45629));
    LocalMux I__10617 (
            .O(N__45629),
            .I(N__45626));
    Odrv4 I__10616 (
            .O(N__45626),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO ));
    InMux I__10615 (
            .O(N__45623),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ));
    InMux I__10614 (
            .O(N__45620),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30 ));
    InMux I__10613 (
            .O(N__45617),
            .I(N__45614));
    LocalMux I__10612 (
            .O(N__45614),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt24 ));
    CascadeMux I__10611 (
            .O(N__45611),
            .I(N__45607));
    InMux I__10610 (
            .O(N__45610),
            .I(N__45603));
    InMux I__10609 (
            .O(N__45607),
            .I(N__45598));
    InMux I__10608 (
            .O(N__45606),
            .I(N__45598));
    LocalMux I__10607 (
            .O(N__45603),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ));
    LocalMux I__10606 (
            .O(N__45598),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ));
    CascadeMux I__10605 (
            .O(N__45593),
            .I(N__45589));
    InMux I__10604 (
            .O(N__45592),
            .I(N__45584));
    InMux I__10603 (
            .O(N__45589),
            .I(N__45584));
    LocalMux I__10602 (
            .O(N__45584),
            .I(N__45581));
    Odrv12 I__10601 (
            .O(N__45581),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ));
    InMux I__10600 (
            .O(N__45578),
            .I(N__45573));
    InMux I__10599 (
            .O(N__45577),
            .I(N__45568));
    InMux I__10598 (
            .O(N__45576),
            .I(N__45568));
    LocalMux I__10597 (
            .O(N__45573),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ));
    LocalMux I__10596 (
            .O(N__45568),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ));
    CascadeMux I__10595 (
            .O(N__45563),
            .I(N__45560));
    InMux I__10594 (
            .O(N__45560),
            .I(N__45557));
    LocalMux I__10593 (
            .O(N__45557),
            .I(N__45554));
    Odrv4 I__10592 (
            .O(N__45554),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ));
    InMux I__10591 (
            .O(N__45551),
            .I(N__45547));
    InMux I__10590 (
            .O(N__45550),
            .I(N__45544));
    LocalMux I__10589 (
            .O(N__45547),
            .I(N__45541));
    LocalMux I__10588 (
            .O(N__45544),
            .I(N__45535));
    Span4Mux_v I__10587 (
            .O(N__45541),
            .I(N__45535));
    InMux I__10586 (
            .O(N__45540),
            .I(N__45532));
    Odrv4 I__10585 (
            .O(N__45535),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    LocalMux I__10584 (
            .O(N__45532),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    InMux I__10583 (
            .O(N__45527),
            .I(N__45524));
    LocalMux I__10582 (
            .O(N__45524),
            .I(N__45519));
    InMux I__10581 (
            .O(N__45523),
            .I(N__45516));
    InMux I__10580 (
            .O(N__45522),
            .I(N__45513));
    Span4Mux_v I__10579 (
            .O(N__45519),
            .I(N__45508));
    LocalMux I__10578 (
            .O(N__45516),
            .I(N__45508));
    LocalMux I__10577 (
            .O(N__45513),
            .I(N__45504));
    Span4Mux_h I__10576 (
            .O(N__45508),
            .I(N__45501));
    InMux I__10575 (
            .O(N__45507),
            .I(N__45498));
    Odrv12 I__10574 (
            .O(N__45504),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    Odrv4 I__10573 (
            .O(N__45501),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    LocalMux I__10572 (
            .O(N__45498),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__10571 (
            .O(N__45491),
            .I(N__45488));
    LocalMux I__10570 (
            .O(N__45488),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    InMux I__10569 (
            .O(N__45485),
            .I(N__45482));
    LocalMux I__10568 (
            .O(N__45482),
            .I(N__45479));
    Odrv12 I__10567 (
            .O(N__45479),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ));
    InMux I__10566 (
            .O(N__45476),
            .I(N__45472));
    InMux I__10565 (
            .O(N__45475),
            .I(N__45469));
    LocalMux I__10564 (
            .O(N__45472),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    LocalMux I__10563 (
            .O(N__45469),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    CascadeMux I__10562 (
            .O(N__45464),
            .I(N__45461));
    InMux I__10561 (
            .O(N__45461),
            .I(N__45458));
    LocalMux I__10560 (
            .O(N__45458),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    InMux I__10559 (
            .O(N__45455),
            .I(N__45451));
    InMux I__10558 (
            .O(N__45454),
            .I(N__45448));
    LocalMux I__10557 (
            .O(N__45451),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    LocalMux I__10556 (
            .O(N__45448),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__10555 (
            .O(N__45443),
            .I(N__45440));
    LocalMux I__10554 (
            .O(N__45440),
            .I(N__45437));
    Span4Mux_h I__10553 (
            .O(N__45437),
            .I(N__45434));
    Odrv4 I__10552 (
            .O(N__45434),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ));
    CascadeMux I__10551 (
            .O(N__45431),
            .I(N__45428));
    InMux I__10550 (
            .O(N__45428),
            .I(N__45425));
    LocalMux I__10549 (
            .O(N__45425),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    InMux I__10548 (
            .O(N__45422),
            .I(N__45418));
    InMux I__10547 (
            .O(N__45421),
            .I(N__45415));
    LocalMux I__10546 (
            .O(N__45418),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    LocalMux I__10545 (
            .O(N__45415),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    CascadeMux I__10544 (
            .O(N__45410),
            .I(N__45407));
    InMux I__10543 (
            .O(N__45407),
            .I(N__45404));
    LocalMux I__10542 (
            .O(N__45404),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    InMux I__10541 (
            .O(N__45401),
            .I(N__45398));
    LocalMux I__10540 (
            .O(N__45398),
            .I(N__45395));
    Odrv4 I__10539 (
            .O(N__45395),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ));
    InMux I__10538 (
            .O(N__45392),
            .I(N__45388));
    InMux I__10537 (
            .O(N__45391),
            .I(N__45385));
    LocalMux I__10536 (
            .O(N__45388),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    LocalMux I__10535 (
            .O(N__45385),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    CascadeMux I__10534 (
            .O(N__45380),
            .I(N__45377));
    InMux I__10533 (
            .O(N__45377),
            .I(N__45374));
    LocalMux I__10532 (
            .O(N__45374),
            .I(N__45371));
    Odrv4 I__10531 (
            .O(N__45371),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    InMux I__10530 (
            .O(N__45368),
            .I(N__45365));
    LocalMux I__10529 (
            .O(N__45365),
            .I(N__45362));
    Span4Mux_h I__10528 (
            .O(N__45362),
            .I(N__45359));
    Odrv4 I__10527 (
            .O(N__45359),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ));
    CascadeMux I__10526 (
            .O(N__45356),
            .I(N__45353));
    InMux I__10525 (
            .O(N__45353),
            .I(N__45350));
    LocalMux I__10524 (
            .O(N__45350),
            .I(N__45347));
    Span4Mux_h I__10523 (
            .O(N__45347),
            .I(N__45344));
    Odrv4 I__10522 (
            .O(N__45344),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt16 ));
    InMux I__10521 (
            .O(N__45341),
            .I(N__45338));
    LocalMux I__10520 (
            .O(N__45338),
            .I(N__45335));
    Span4Mux_v I__10519 (
            .O(N__45335),
            .I(N__45332));
    Odrv4 I__10518 (
            .O(N__45332),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ));
    CascadeMux I__10517 (
            .O(N__45329),
            .I(N__45326));
    InMux I__10516 (
            .O(N__45326),
            .I(N__45323));
    LocalMux I__10515 (
            .O(N__45323),
            .I(N__45320));
    Span4Mux_v I__10514 (
            .O(N__45320),
            .I(N__45317));
    Odrv4 I__10513 (
            .O(N__45317),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt18 ));
    InMux I__10512 (
            .O(N__45314),
            .I(N__45311));
    LocalMux I__10511 (
            .O(N__45311),
            .I(N__45308));
    Odrv4 I__10510 (
            .O(N__45308),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ));
    CascadeMux I__10509 (
            .O(N__45305),
            .I(N__45302));
    InMux I__10508 (
            .O(N__45302),
            .I(N__45299));
    LocalMux I__10507 (
            .O(N__45299),
            .I(N__45296));
    Odrv4 I__10506 (
            .O(N__45296),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt20 ));
    CascadeMux I__10505 (
            .O(N__45293),
            .I(N__45290));
    InMux I__10504 (
            .O(N__45290),
            .I(N__45287));
    LocalMux I__10503 (
            .O(N__45287),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ));
    InMux I__10502 (
            .O(N__45284),
            .I(N__45280));
    InMux I__10501 (
            .O(N__45283),
            .I(N__45277));
    LocalMux I__10500 (
            .O(N__45280),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__10499 (
            .O(N__45277),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__10498 (
            .O(N__45272),
            .I(N__45269));
    LocalMux I__10497 (
            .O(N__45269),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    InMux I__10496 (
            .O(N__45266),
            .I(N__45262));
    InMux I__10495 (
            .O(N__45265),
            .I(N__45259));
    LocalMux I__10494 (
            .O(N__45262),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__10493 (
            .O(N__45259),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    CascadeMux I__10492 (
            .O(N__45254),
            .I(N__45251));
    InMux I__10491 (
            .O(N__45251),
            .I(N__45248));
    LocalMux I__10490 (
            .O(N__45248),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ));
    InMux I__10489 (
            .O(N__45245),
            .I(N__45242));
    LocalMux I__10488 (
            .O(N__45242),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    InMux I__10487 (
            .O(N__45239),
            .I(N__45236));
    LocalMux I__10486 (
            .O(N__45236),
            .I(N__45233));
    Odrv12 I__10485 (
            .O(N__45233),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ));
    InMux I__10484 (
            .O(N__45230),
            .I(N__45226));
    InMux I__10483 (
            .O(N__45229),
            .I(N__45223));
    LocalMux I__10482 (
            .O(N__45226),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__10481 (
            .O(N__45223),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    CascadeMux I__10480 (
            .O(N__45218),
            .I(N__45215));
    InMux I__10479 (
            .O(N__45215),
            .I(N__45212));
    LocalMux I__10478 (
            .O(N__45212),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    InMux I__10477 (
            .O(N__45209),
            .I(N__45206));
    LocalMux I__10476 (
            .O(N__45206),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ));
    InMux I__10475 (
            .O(N__45203),
            .I(N__45199));
    InMux I__10474 (
            .O(N__45202),
            .I(N__45196));
    LocalMux I__10473 (
            .O(N__45199),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__10472 (
            .O(N__45196),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    CascadeMux I__10471 (
            .O(N__45191),
            .I(N__45188));
    InMux I__10470 (
            .O(N__45188),
            .I(N__45185));
    LocalMux I__10469 (
            .O(N__45185),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    InMux I__10468 (
            .O(N__45182),
            .I(N__45179));
    LocalMux I__10467 (
            .O(N__45179),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ));
    InMux I__10466 (
            .O(N__45176),
            .I(N__45172));
    InMux I__10465 (
            .O(N__45175),
            .I(N__45169));
    LocalMux I__10464 (
            .O(N__45172),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    LocalMux I__10463 (
            .O(N__45169),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    CascadeMux I__10462 (
            .O(N__45164),
            .I(N__45161));
    InMux I__10461 (
            .O(N__45161),
            .I(N__45158));
    LocalMux I__10460 (
            .O(N__45158),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    InMux I__10459 (
            .O(N__45155),
            .I(N__45152));
    LocalMux I__10458 (
            .O(N__45152),
            .I(N__45149));
    Odrv12 I__10457 (
            .O(N__45149),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ));
    InMux I__10456 (
            .O(N__45146),
            .I(N__45142));
    InMux I__10455 (
            .O(N__45145),
            .I(N__45139));
    LocalMux I__10454 (
            .O(N__45142),
            .I(N__45136));
    LocalMux I__10453 (
            .O(N__45139),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__10452 (
            .O(N__45136),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    CascadeMux I__10451 (
            .O(N__45131),
            .I(N__45128));
    InMux I__10450 (
            .O(N__45128),
            .I(N__45125));
    LocalMux I__10449 (
            .O(N__45125),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    InMux I__10448 (
            .O(N__45122),
            .I(N__45118));
    InMux I__10447 (
            .O(N__45121),
            .I(N__45115));
    LocalMux I__10446 (
            .O(N__45118),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    LocalMux I__10445 (
            .O(N__45115),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__10444 (
            .O(N__45110),
            .I(N__45107));
    LocalMux I__10443 (
            .O(N__45107),
            .I(N__45104));
    Odrv4 I__10442 (
            .O(N__45104),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ));
    CascadeMux I__10441 (
            .O(N__45101),
            .I(N__45098));
    InMux I__10440 (
            .O(N__45098),
            .I(N__45095));
    LocalMux I__10439 (
            .O(N__45095),
            .I(N__45092));
    Odrv4 I__10438 (
            .O(N__45092),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    InMux I__10437 (
            .O(N__45089),
            .I(N__45085));
    InMux I__10436 (
            .O(N__45088),
            .I(N__45082));
    LocalMux I__10435 (
            .O(N__45085),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    LocalMux I__10434 (
            .O(N__45082),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__10433 (
            .O(N__45077),
            .I(N__45073));
    InMux I__10432 (
            .O(N__45076),
            .I(N__45069));
    LocalMux I__10431 (
            .O(N__45073),
            .I(N__45066));
    InMux I__10430 (
            .O(N__45072),
            .I(N__45063));
    LocalMux I__10429 (
            .O(N__45069),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    Odrv4 I__10428 (
            .O(N__45066),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    LocalMux I__10427 (
            .O(N__45063),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    InMux I__10426 (
            .O(N__45056),
            .I(N__45052));
    InMux I__10425 (
            .O(N__45055),
            .I(N__45049));
    LocalMux I__10424 (
            .O(N__45052),
            .I(N__45045));
    LocalMux I__10423 (
            .O(N__45049),
            .I(N__45042));
    InMux I__10422 (
            .O(N__45048),
            .I(N__45039));
    Span4Mux_v I__10421 (
            .O(N__45045),
            .I(N__45036));
    Span4Mux_h I__10420 (
            .O(N__45042),
            .I(N__45033));
    LocalMux I__10419 (
            .O(N__45039),
            .I(N__45030));
    Span4Mux_v I__10418 (
            .O(N__45036),
            .I(N__45026));
    Span4Mux_v I__10417 (
            .O(N__45033),
            .I(N__45023));
    Span12Mux_v I__10416 (
            .O(N__45030),
            .I(N__45020));
    InMux I__10415 (
            .O(N__45029),
            .I(N__45017));
    Odrv4 I__10414 (
            .O(N__45026),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    Odrv4 I__10413 (
            .O(N__45023),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    Odrv12 I__10412 (
            .O(N__45020),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    LocalMux I__10411 (
            .O(N__45017),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__10410 (
            .O(N__45008),
            .I(N__45005));
    LocalMux I__10409 (
            .O(N__45005),
            .I(N__44999));
    InMux I__10408 (
            .O(N__45004),
            .I(N__44996));
    InMux I__10407 (
            .O(N__45003),
            .I(N__44993));
    InMux I__10406 (
            .O(N__45002),
            .I(N__44990));
    Span4Mux_h I__10405 (
            .O(N__44999),
            .I(N__44987));
    LocalMux I__10404 (
            .O(N__44996),
            .I(N__44982));
    LocalMux I__10403 (
            .O(N__44993),
            .I(N__44982));
    LocalMux I__10402 (
            .O(N__44990),
            .I(N__44979));
    Span4Mux_v I__10401 (
            .O(N__44987),
            .I(N__44976));
    Span4Mux_v I__10400 (
            .O(N__44982),
            .I(N__44971));
    Span4Mux_h I__10399 (
            .O(N__44979),
            .I(N__44971));
    Odrv4 I__10398 (
            .O(N__44976),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    Odrv4 I__10397 (
            .O(N__44971),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    InMux I__10396 (
            .O(N__44966),
            .I(N__44961));
    InMux I__10395 (
            .O(N__44965),
            .I(N__44958));
    InMux I__10394 (
            .O(N__44964),
            .I(N__44955));
    LocalMux I__10393 (
            .O(N__44961),
            .I(N__44952));
    LocalMux I__10392 (
            .O(N__44958),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    LocalMux I__10391 (
            .O(N__44955),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    Odrv4 I__10390 (
            .O(N__44952),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    InMux I__10389 (
            .O(N__44945),
            .I(N__44942));
    LocalMux I__10388 (
            .O(N__44942),
            .I(N__44938));
    InMux I__10387 (
            .O(N__44941),
            .I(N__44934));
    Span4Mux_h I__10386 (
            .O(N__44938),
            .I(N__44931));
    InMux I__10385 (
            .O(N__44937),
            .I(N__44928));
    LocalMux I__10384 (
            .O(N__44934),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    Odrv4 I__10383 (
            .O(N__44931),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    LocalMux I__10382 (
            .O(N__44928),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    InMux I__10381 (
            .O(N__44921),
            .I(N__44916));
    InMux I__10380 (
            .O(N__44920),
            .I(N__44912));
    InMux I__10379 (
            .O(N__44919),
            .I(N__44909));
    LocalMux I__10378 (
            .O(N__44916),
            .I(N__44906));
    InMux I__10377 (
            .O(N__44915),
            .I(N__44903));
    LocalMux I__10376 (
            .O(N__44912),
            .I(N__44898));
    LocalMux I__10375 (
            .O(N__44909),
            .I(N__44898));
    Span4Mux_v I__10374 (
            .O(N__44906),
            .I(N__44893));
    LocalMux I__10373 (
            .O(N__44903),
            .I(N__44893));
    Span4Mux_v I__10372 (
            .O(N__44898),
            .I(N__44890));
    Span4Mux_h I__10371 (
            .O(N__44893),
            .I(N__44887));
    Odrv4 I__10370 (
            .O(N__44890),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    Odrv4 I__10369 (
            .O(N__44887),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    InMux I__10368 (
            .O(N__44882),
            .I(N__44879));
    LocalMux I__10367 (
            .O(N__44879),
            .I(N__44874));
    InMux I__10366 (
            .O(N__44878),
            .I(N__44871));
    InMux I__10365 (
            .O(N__44877),
            .I(N__44868));
    Span4Mux_h I__10364 (
            .O(N__44874),
            .I(N__44865));
    LocalMux I__10363 (
            .O(N__44871),
            .I(N__44862));
    LocalMux I__10362 (
            .O(N__44868),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    Odrv4 I__10361 (
            .O(N__44865),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    Odrv12 I__10360 (
            .O(N__44862),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    InMux I__10359 (
            .O(N__44855),
            .I(N__44850));
    InMux I__10358 (
            .O(N__44854),
            .I(N__44846));
    InMux I__10357 (
            .O(N__44853),
            .I(N__44843));
    LocalMux I__10356 (
            .O(N__44850),
            .I(N__44840));
    InMux I__10355 (
            .O(N__44849),
            .I(N__44837));
    LocalMux I__10354 (
            .O(N__44846),
            .I(N__44834));
    LocalMux I__10353 (
            .O(N__44843),
            .I(N__44831));
    Span4Mux_v I__10352 (
            .O(N__44840),
            .I(N__44826));
    LocalMux I__10351 (
            .O(N__44837),
            .I(N__44826));
    Span4Mux_v I__10350 (
            .O(N__44834),
            .I(N__44823));
    Span4Mux_v I__10349 (
            .O(N__44831),
            .I(N__44818));
    Span4Mux_h I__10348 (
            .O(N__44826),
            .I(N__44818));
    Odrv4 I__10347 (
            .O(N__44823),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    Odrv4 I__10346 (
            .O(N__44818),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    InMux I__10345 (
            .O(N__44813),
            .I(N__44810));
    LocalMux I__10344 (
            .O(N__44810),
            .I(N__44806));
    InMux I__10343 (
            .O(N__44809),
            .I(N__44802));
    Span4Mux_h I__10342 (
            .O(N__44806),
            .I(N__44799));
    InMux I__10341 (
            .O(N__44805),
            .I(N__44796));
    LocalMux I__10340 (
            .O(N__44802),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    Odrv4 I__10339 (
            .O(N__44799),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    LocalMux I__10338 (
            .O(N__44796),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    InMux I__10337 (
            .O(N__44789),
            .I(N__44784));
    InMux I__10336 (
            .O(N__44788),
            .I(N__44781));
    InMux I__10335 (
            .O(N__44787),
            .I(N__44778));
    LocalMux I__10334 (
            .O(N__44784),
            .I(N__44773));
    LocalMux I__10333 (
            .O(N__44781),
            .I(N__44773));
    LocalMux I__10332 (
            .O(N__44778),
            .I(N__44770));
    Span4Mux_h I__10331 (
            .O(N__44773),
            .I(N__44767));
    Span4Mux_h I__10330 (
            .O(N__44770),
            .I(N__44763));
    Span4Mux_v I__10329 (
            .O(N__44767),
            .I(N__44760));
    InMux I__10328 (
            .O(N__44766),
            .I(N__44757));
    Odrv4 I__10327 (
            .O(N__44763),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    Odrv4 I__10326 (
            .O(N__44760),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    LocalMux I__10325 (
            .O(N__44757),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    CascadeMux I__10324 (
            .O(N__44750),
            .I(N__44747));
    InMux I__10323 (
            .O(N__44747),
            .I(N__44741));
    InMux I__10322 (
            .O(N__44746),
            .I(N__44741));
    LocalMux I__10321 (
            .O(N__44741),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ));
    CascadeMux I__10320 (
            .O(N__44738),
            .I(N__44735));
    InMux I__10319 (
            .O(N__44735),
            .I(N__44730));
    InMux I__10318 (
            .O(N__44734),
            .I(N__44727));
    CascadeMux I__10317 (
            .O(N__44733),
            .I(N__44724));
    LocalMux I__10316 (
            .O(N__44730),
            .I(N__44721));
    LocalMux I__10315 (
            .O(N__44727),
            .I(N__44718));
    InMux I__10314 (
            .O(N__44724),
            .I(N__44715));
    Span12Mux_h I__10313 (
            .O(N__44721),
            .I(N__44712));
    Span4Mux_h I__10312 (
            .O(N__44718),
            .I(N__44709));
    LocalMux I__10311 (
            .O(N__44715),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv12 I__10310 (
            .O(N__44712),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__10309 (
            .O(N__44709),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__10308 (
            .O(N__44702),
            .I(N__44699));
    LocalMux I__10307 (
            .O(N__44699),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__10306 (
            .O(N__44696),
            .I(N__44693));
    InMux I__10305 (
            .O(N__44693),
            .I(N__44690));
    LocalMux I__10304 (
            .O(N__44690),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    InMux I__10303 (
            .O(N__44687),
            .I(N__44683));
    InMux I__10302 (
            .O(N__44686),
            .I(N__44680));
    LocalMux I__10301 (
            .O(N__44683),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__10300 (
            .O(N__44680),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    CascadeMux I__10299 (
            .O(N__44675),
            .I(N__44672));
    InMux I__10298 (
            .O(N__44672),
            .I(N__44669));
    LocalMux I__10297 (
            .O(N__44669),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ));
    InMux I__10296 (
            .O(N__44666),
            .I(N__44663));
    LocalMux I__10295 (
            .O(N__44663),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    CascadeMux I__10294 (
            .O(N__44660),
            .I(N__44657));
    InMux I__10293 (
            .O(N__44657),
            .I(N__44654));
    LocalMux I__10292 (
            .O(N__44654),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ));
    InMux I__10291 (
            .O(N__44651),
            .I(N__44647));
    InMux I__10290 (
            .O(N__44650),
            .I(N__44644));
    LocalMux I__10289 (
            .O(N__44647),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__10288 (
            .O(N__44644),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__10287 (
            .O(N__44639),
            .I(N__44636));
    LocalMux I__10286 (
            .O(N__44636),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    InMux I__10285 (
            .O(N__44633),
            .I(N__44628));
    CascadeMux I__10284 (
            .O(N__44632),
            .I(N__44624));
    InMux I__10283 (
            .O(N__44631),
            .I(N__44621));
    LocalMux I__10282 (
            .O(N__44628),
            .I(N__44618));
    InMux I__10281 (
            .O(N__44627),
            .I(N__44613));
    InMux I__10280 (
            .O(N__44624),
            .I(N__44613));
    LocalMux I__10279 (
            .O(N__44621),
            .I(N__44606));
    Span4Mux_h I__10278 (
            .O(N__44618),
            .I(N__44606));
    LocalMux I__10277 (
            .O(N__44613),
            .I(N__44606));
    Odrv4 I__10276 (
            .O(N__44606),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    IoInMux I__10275 (
            .O(N__44603),
            .I(N__44600));
    LocalMux I__10274 (
            .O(N__44600),
            .I(N__44597));
    Span4Mux_s1_v I__10273 (
            .O(N__44597),
            .I(N__44594));
    Span4Mux_v I__10272 (
            .O(N__44594),
            .I(N__44591));
    Span4Mux_v I__10271 (
            .O(N__44591),
            .I(N__44587));
    InMux I__10270 (
            .O(N__44590),
            .I(N__44584));
    Odrv4 I__10269 (
            .O(N__44587),
            .I(T12_c));
    LocalMux I__10268 (
            .O(N__44584),
            .I(T12_c));
    InMux I__10267 (
            .O(N__44579),
            .I(N__44572));
    InMux I__10266 (
            .O(N__44578),
            .I(N__44572));
    InMux I__10265 (
            .O(N__44577),
            .I(N__44569));
    LocalMux I__10264 (
            .O(N__44572),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    LocalMux I__10263 (
            .O(N__44569),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    InMux I__10262 (
            .O(N__44564),
            .I(N__44560));
    InMux I__10261 (
            .O(N__44563),
            .I(N__44557));
    LocalMux I__10260 (
            .O(N__44560),
            .I(N__44554));
    LocalMux I__10259 (
            .O(N__44557),
            .I(N__44551));
    Span4Mux_h I__10258 (
            .O(N__44554),
            .I(N__44546));
    Span4Mux_v I__10257 (
            .O(N__44551),
            .I(N__44546));
    Odrv4 I__10256 (
            .O(N__44546),
            .I(\phase_controller_inst1.state_RNI7NN7Z0Z_0 ));
    InMux I__10255 (
            .O(N__44543),
            .I(N__44540));
    LocalMux I__10254 (
            .O(N__44540),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ));
    InMux I__10253 (
            .O(N__44537),
            .I(N__44534));
    LocalMux I__10252 (
            .O(N__44534),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ));
    CascadeMux I__10251 (
            .O(N__44531),
            .I(N__44528));
    InMux I__10250 (
            .O(N__44528),
            .I(N__44525));
    LocalMux I__10249 (
            .O(N__44525),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ));
    InMux I__10248 (
            .O(N__44522),
            .I(N__44519));
    LocalMux I__10247 (
            .O(N__44519),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ));
    InMux I__10246 (
            .O(N__44516),
            .I(N__44513));
    LocalMux I__10245 (
            .O(N__44513),
            .I(N__44510));
    Span4Mux_v I__10244 (
            .O(N__44510),
            .I(N__44506));
    InMux I__10243 (
            .O(N__44509),
            .I(N__44503));
    Odrv4 I__10242 (
            .O(N__44506),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    LocalMux I__10241 (
            .O(N__44503),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    InMux I__10240 (
            .O(N__44498),
            .I(N__44495));
    LocalMux I__10239 (
            .O(N__44495),
            .I(N__44492));
    Span4Mux_v I__10238 (
            .O(N__44492),
            .I(N__44488));
    InMux I__10237 (
            .O(N__44491),
            .I(N__44485));
    Odrv4 I__10236 (
            .O(N__44488),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    LocalMux I__10235 (
            .O(N__44485),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    CascadeMux I__10234 (
            .O(N__44480),
            .I(N__44477));
    InMux I__10233 (
            .O(N__44477),
            .I(N__44473));
    CascadeMux I__10232 (
            .O(N__44476),
            .I(N__44470));
    LocalMux I__10231 (
            .O(N__44473),
            .I(N__44467));
    InMux I__10230 (
            .O(N__44470),
            .I(N__44464));
    Odrv4 I__10229 (
            .O(N__44467),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    LocalMux I__10228 (
            .O(N__44464),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    InMux I__10227 (
            .O(N__44459),
            .I(N__44456));
    LocalMux I__10226 (
            .O(N__44456),
            .I(N__44452));
    InMux I__10225 (
            .O(N__44455),
            .I(N__44449));
    Odrv4 I__10224 (
            .O(N__44452),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    LocalMux I__10223 (
            .O(N__44449),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    InMux I__10222 (
            .O(N__44444),
            .I(N__44441));
    LocalMux I__10221 (
            .O(N__44441),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    InMux I__10220 (
            .O(N__44438),
            .I(N__44435));
    LocalMux I__10219 (
            .O(N__44435),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ));
    CascadeMux I__10218 (
            .O(N__44432),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9_cascade_ ));
    InMux I__10217 (
            .O(N__44429),
            .I(N__44426));
    LocalMux I__10216 (
            .O(N__44426),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ));
    InMux I__10215 (
            .O(N__44423),
            .I(N__44420));
    LocalMux I__10214 (
            .O(N__44420),
            .I(N__44416));
    InMux I__10213 (
            .O(N__44419),
            .I(N__44413));
    Span12Mux_v I__10212 (
            .O(N__44416),
            .I(N__44408));
    LocalMux I__10211 (
            .O(N__44413),
            .I(N__44408));
    Span12Mux_h I__10210 (
            .O(N__44408),
            .I(N__44405));
    Odrv12 I__10209 (
            .O(N__44405),
            .I(\pwm_generator_inst.O_10 ));
    CascadeMux I__10208 (
            .O(N__44402),
            .I(N__44399));
    InMux I__10207 (
            .O(N__44399),
            .I(N__44396));
    LocalMux I__10206 (
            .O(N__44396),
            .I(N__44391));
    InMux I__10205 (
            .O(N__44395),
            .I(N__44388));
    InMux I__10204 (
            .O(N__44394),
            .I(N__44385));
    Span4Mux_h I__10203 (
            .O(N__44391),
            .I(N__44382));
    LocalMux I__10202 (
            .O(N__44388),
            .I(N__44379));
    LocalMux I__10201 (
            .O(N__44385),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    Odrv4 I__10200 (
            .O(N__44382),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    Odrv4 I__10199 (
            .O(N__44379),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    InMux I__10198 (
            .O(N__44372),
            .I(N__44368));
    InMux I__10197 (
            .O(N__44371),
            .I(N__44364));
    LocalMux I__10196 (
            .O(N__44368),
            .I(N__44361));
    InMux I__10195 (
            .O(N__44367),
            .I(N__44358));
    LocalMux I__10194 (
            .O(N__44364),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    Odrv4 I__10193 (
            .O(N__44361),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    LocalMux I__10192 (
            .O(N__44358),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    InMux I__10191 (
            .O(N__44351),
            .I(N__44346));
    InMux I__10190 (
            .O(N__44350),
            .I(N__44342));
    InMux I__10189 (
            .O(N__44349),
            .I(N__44339));
    LocalMux I__10188 (
            .O(N__44346),
            .I(N__44336));
    InMux I__10187 (
            .O(N__44345),
            .I(N__44333));
    LocalMux I__10186 (
            .O(N__44342),
            .I(N__44330));
    LocalMux I__10185 (
            .O(N__44339),
            .I(N__44327));
    Span4Mux_h I__10184 (
            .O(N__44336),
            .I(N__44324));
    LocalMux I__10183 (
            .O(N__44333),
            .I(N__44321));
    Span12Mux_s7_v I__10182 (
            .O(N__44330),
            .I(N__44318));
    Span12Mux_v I__10181 (
            .O(N__44327),
            .I(N__44315));
    Span4Mux_v I__10180 (
            .O(N__44324),
            .I(N__44310));
    Span4Mux_h I__10179 (
            .O(N__44321),
            .I(N__44310));
    Odrv12 I__10178 (
            .O(N__44318),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    Odrv12 I__10177 (
            .O(N__44315),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    Odrv4 I__10176 (
            .O(N__44310),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    InMux I__10175 (
            .O(N__44303),
            .I(N__44299));
    InMux I__10174 (
            .O(N__44302),
            .I(N__44294));
    LocalMux I__10173 (
            .O(N__44299),
            .I(N__44291));
    InMux I__10172 (
            .O(N__44298),
            .I(N__44288));
    InMux I__10171 (
            .O(N__44297),
            .I(N__44285));
    LocalMux I__10170 (
            .O(N__44294),
            .I(N__44282));
    Span4Mux_v I__10169 (
            .O(N__44291),
            .I(N__44279));
    LocalMux I__10168 (
            .O(N__44288),
            .I(N__44276));
    LocalMux I__10167 (
            .O(N__44285),
            .I(N__44273));
    Span4Mux_v I__10166 (
            .O(N__44282),
            .I(N__44268));
    Span4Mux_h I__10165 (
            .O(N__44279),
            .I(N__44268));
    Span4Mux_v I__10164 (
            .O(N__44276),
            .I(N__44263));
    Span4Mux_h I__10163 (
            .O(N__44273),
            .I(N__44263));
    Odrv4 I__10162 (
            .O(N__44268),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    Odrv4 I__10161 (
            .O(N__44263),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    InMux I__10160 (
            .O(N__44258),
            .I(N__44254));
    InMux I__10159 (
            .O(N__44257),
            .I(N__44250));
    LocalMux I__10158 (
            .O(N__44254),
            .I(N__44247));
    InMux I__10157 (
            .O(N__44253),
            .I(N__44244));
    LocalMux I__10156 (
            .O(N__44250),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    Odrv4 I__10155 (
            .O(N__44247),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    LocalMux I__10154 (
            .O(N__44244),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    CascadeMux I__10153 (
            .O(N__44237),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28_cascade_));
    InMux I__10152 (
            .O(N__44234),
            .I(N__44226));
    InMux I__10151 (
            .O(N__44233),
            .I(N__44226));
    InMux I__10150 (
            .O(N__44232),
            .I(N__44223));
    InMux I__10149 (
            .O(N__44231),
            .I(N__44220));
    LocalMux I__10148 (
            .O(N__44226),
            .I(N__44217));
    LocalMux I__10147 (
            .O(N__44223),
            .I(N__44214));
    LocalMux I__10146 (
            .O(N__44220),
            .I(N__44211));
    Span4Mux_h I__10145 (
            .O(N__44217),
            .I(N__44208));
    Span4Mux_h I__10144 (
            .O(N__44214),
            .I(N__44203));
    Span4Mux_v I__10143 (
            .O(N__44211),
            .I(N__44203));
    Odrv4 I__10142 (
            .O(N__44208),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    Odrv4 I__10141 (
            .O(N__44203),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__10140 (
            .O(N__44198),
            .I(N__44193));
    InMux I__10139 (
            .O(N__44197),
            .I(N__44188));
    InMux I__10138 (
            .O(N__44196),
            .I(N__44188));
    LocalMux I__10137 (
            .O(N__44193),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ));
    LocalMux I__10136 (
            .O(N__44188),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ));
    CascadeMux I__10135 (
            .O(N__44183),
            .I(N__44180));
    InMux I__10134 (
            .O(N__44180),
            .I(N__44174));
    InMux I__10133 (
            .O(N__44179),
            .I(N__44174));
    LocalMux I__10132 (
            .O(N__44174),
            .I(N__44171));
    Span4Mux_h I__10131 (
            .O(N__44171),
            .I(N__44168));
    Odrv4 I__10130 (
            .O(N__44168),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ));
    CascadeMux I__10129 (
            .O(N__44165),
            .I(N__44160));
    InMux I__10128 (
            .O(N__44164),
            .I(N__44157));
    InMux I__10127 (
            .O(N__44163),
            .I(N__44152));
    InMux I__10126 (
            .O(N__44160),
            .I(N__44152));
    LocalMux I__10125 (
            .O(N__44157),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ));
    LocalMux I__10124 (
            .O(N__44152),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ));
    InMux I__10123 (
            .O(N__44147),
            .I(N__44141));
    InMux I__10122 (
            .O(N__44146),
            .I(N__44141));
    LocalMux I__10121 (
            .O(N__44141),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ));
    CascadeMux I__10120 (
            .O(N__44138),
            .I(N__44133));
    InMux I__10119 (
            .O(N__44137),
            .I(N__44126));
    InMux I__10118 (
            .O(N__44136),
            .I(N__44126));
    InMux I__10117 (
            .O(N__44133),
            .I(N__44126));
    LocalMux I__10116 (
            .O(N__44126),
            .I(N__44123));
    Span4Mux_h I__10115 (
            .O(N__44123),
            .I(N__44120));
    Odrv4 I__10114 (
            .O(N__44120),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ));
    CEMux I__10113 (
            .O(N__44117),
            .I(N__44113));
    CEMux I__10112 (
            .O(N__44116),
            .I(N__44109));
    LocalMux I__10111 (
            .O(N__44113),
            .I(N__44105));
    CEMux I__10110 (
            .O(N__44112),
            .I(N__44102));
    LocalMux I__10109 (
            .O(N__44109),
            .I(N__44099));
    CEMux I__10108 (
            .O(N__44108),
            .I(N__44096));
    Span4Mux_h I__10107 (
            .O(N__44105),
            .I(N__44092));
    LocalMux I__10106 (
            .O(N__44102),
            .I(N__44089));
    Span4Mux_v I__10105 (
            .O(N__44099),
            .I(N__44086));
    LocalMux I__10104 (
            .O(N__44096),
            .I(N__44083));
    CEMux I__10103 (
            .O(N__44095),
            .I(N__44080));
    Span4Mux_v I__10102 (
            .O(N__44092),
            .I(N__44075));
    Span4Mux_h I__10101 (
            .O(N__44089),
            .I(N__44075));
    Span4Mux_h I__10100 (
            .O(N__44086),
            .I(N__44072));
    Span4Mux_h I__10099 (
            .O(N__44083),
            .I(N__44069));
    LocalMux I__10098 (
            .O(N__44080),
            .I(N__44066));
    Odrv4 I__10097 (
            .O(N__44075),
            .I(\delay_measurement_inst.delay_tr_timer.N_200_i ));
    Odrv4 I__10096 (
            .O(N__44072),
            .I(\delay_measurement_inst.delay_tr_timer.N_200_i ));
    Odrv4 I__10095 (
            .O(N__44069),
            .I(\delay_measurement_inst.delay_tr_timer.N_200_i ));
    Odrv12 I__10094 (
            .O(N__44066),
            .I(\delay_measurement_inst.delay_tr_timer.N_200_i ));
    InMux I__10093 (
            .O(N__44057),
            .I(N__44052));
    InMux I__10092 (
            .O(N__44056),
            .I(N__44049));
    CascadeMux I__10091 (
            .O(N__44055),
            .I(N__44046));
    LocalMux I__10090 (
            .O(N__44052),
            .I(N__44043));
    LocalMux I__10089 (
            .O(N__44049),
            .I(N__44039));
    InMux I__10088 (
            .O(N__44046),
            .I(N__44036));
    Span12Mux_v I__10087 (
            .O(N__44043),
            .I(N__44033));
    InMux I__10086 (
            .O(N__44042),
            .I(N__44030));
    Span12Mux_s11_v I__10085 (
            .O(N__44039),
            .I(N__44027));
    LocalMux I__10084 (
            .O(N__44036),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv12 I__10083 (
            .O(N__44033),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__10082 (
            .O(N__44030),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv12 I__10081 (
            .O(N__44027),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    InMux I__10080 (
            .O(N__44018),
            .I(N__44013));
    InMux I__10079 (
            .O(N__44017),
            .I(N__44010));
    InMux I__10078 (
            .O(N__44016),
            .I(N__44007));
    LocalMux I__10077 (
            .O(N__44013),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    LocalMux I__10076 (
            .O(N__44010),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    LocalMux I__10075 (
            .O(N__44007),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    InMux I__10074 (
            .O(N__44000),
            .I(N__43996));
    InMux I__10073 (
            .O(N__43999),
            .I(N__43992));
    LocalMux I__10072 (
            .O(N__43996),
            .I(N__43989));
    InMux I__10071 (
            .O(N__43995),
            .I(N__43986));
    LocalMux I__10070 (
            .O(N__43992),
            .I(N__43978));
    Span4Mux_v I__10069 (
            .O(N__43989),
            .I(N__43978));
    LocalMux I__10068 (
            .O(N__43986),
            .I(N__43978));
    InMux I__10067 (
            .O(N__43985),
            .I(N__43975));
    Odrv4 I__10066 (
            .O(N__43978),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__10065 (
            .O(N__43975),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    InMux I__10064 (
            .O(N__43970),
            .I(N__43967));
    LocalMux I__10063 (
            .O(N__43967),
            .I(N__43961));
    InMux I__10062 (
            .O(N__43966),
            .I(N__43958));
    InMux I__10061 (
            .O(N__43965),
            .I(N__43955));
    InMux I__10060 (
            .O(N__43964),
            .I(N__43952));
    Span4Mux_v I__10059 (
            .O(N__43961),
            .I(N__43949));
    LocalMux I__10058 (
            .O(N__43958),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    LocalMux I__10057 (
            .O(N__43955),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    LocalMux I__10056 (
            .O(N__43952),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    Odrv4 I__10055 (
            .O(N__43949),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    CEMux I__10054 (
            .O(N__43940),
            .I(N__43935));
    CEMux I__10053 (
            .O(N__43939),
            .I(N__43931));
    CEMux I__10052 (
            .O(N__43938),
            .I(N__43928));
    LocalMux I__10051 (
            .O(N__43935),
            .I(N__43925));
    CEMux I__10050 (
            .O(N__43934),
            .I(N__43922));
    LocalMux I__10049 (
            .O(N__43931),
            .I(N__43919));
    LocalMux I__10048 (
            .O(N__43928),
            .I(N__43916));
    Span4Mux_v I__10047 (
            .O(N__43925),
            .I(N__43911));
    LocalMux I__10046 (
            .O(N__43922),
            .I(N__43911));
    Span4Mux_h I__10045 (
            .O(N__43919),
            .I(N__43908));
    Span4Mux_h I__10044 (
            .O(N__43916),
            .I(N__43905));
    Span4Mux_h I__10043 (
            .O(N__43911),
            .I(N__43902));
    Odrv4 I__10042 (
            .O(N__43908),
            .I(\delay_measurement_inst.delay_tr_timer.N_201_i ));
    Odrv4 I__10041 (
            .O(N__43905),
            .I(\delay_measurement_inst.delay_tr_timer.N_201_i ));
    Odrv4 I__10040 (
            .O(N__43902),
            .I(\delay_measurement_inst.delay_tr_timer.N_201_i ));
    InMux I__10039 (
            .O(N__43895),
            .I(bfn_17_14_0_));
    InMux I__10038 (
            .O(N__43892),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ));
    InMux I__10037 (
            .O(N__43889),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ));
    InMux I__10036 (
            .O(N__43886),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ));
    InMux I__10035 (
            .O(N__43883),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ));
    InMux I__10034 (
            .O(N__43880),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ));
    InMux I__10033 (
            .O(N__43877),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ));
    InMux I__10032 (
            .O(N__43874),
            .I(N__43870));
    InMux I__10031 (
            .O(N__43873),
            .I(N__43865));
    LocalMux I__10030 (
            .O(N__43870),
            .I(N__43862));
    InMux I__10029 (
            .O(N__43869),
            .I(N__43859));
    InMux I__10028 (
            .O(N__43868),
            .I(N__43856));
    LocalMux I__10027 (
            .O(N__43865),
            .I(N__43853));
    Span4Mux_h I__10026 (
            .O(N__43862),
            .I(N__43848));
    LocalMux I__10025 (
            .O(N__43859),
            .I(N__43848));
    LocalMux I__10024 (
            .O(N__43856),
            .I(N__43845));
    Span4Mux_h I__10023 (
            .O(N__43853),
            .I(N__43842));
    Span4Mux_v I__10022 (
            .O(N__43848),
            .I(N__43839));
    Odrv12 I__10021 (
            .O(N__43845),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    Odrv4 I__10020 (
            .O(N__43842),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    Odrv4 I__10019 (
            .O(N__43839),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__10018 (
            .O(N__43832),
            .I(N__43829));
    LocalMux I__10017 (
            .O(N__43829),
            .I(N__43825));
    InMux I__10016 (
            .O(N__43828),
            .I(N__43821));
    Span4Mux_v I__10015 (
            .O(N__43825),
            .I(N__43818));
    InMux I__10014 (
            .O(N__43824),
            .I(N__43815));
    LocalMux I__10013 (
            .O(N__43821),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    Odrv4 I__10012 (
            .O(N__43818),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    LocalMux I__10011 (
            .O(N__43815),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    InMux I__10010 (
            .O(N__43808),
            .I(N__43805));
    LocalMux I__10009 (
            .O(N__43805),
            .I(N__43802));
    Span4Mux_v I__10008 (
            .O(N__43802),
            .I(N__43798));
    InMux I__10007 (
            .O(N__43801),
            .I(N__43795));
    Odrv4 I__10006 (
            .O(N__43798),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    LocalMux I__10005 (
            .O(N__43795),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    InMux I__10004 (
            .O(N__43790),
            .I(N__43785));
    InMux I__10003 (
            .O(N__43789),
            .I(N__43780));
    InMux I__10002 (
            .O(N__43788),
            .I(N__43780));
    LocalMux I__10001 (
            .O(N__43785),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    LocalMux I__10000 (
            .O(N__43780),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__9999 (
            .O(N__43775),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ));
    CascadeMux I__9998 (
            .O(N__43772),
            .I(N__43767));
    CascadeMux I__9997 (
            .O(N__43771),
            .I(N__43764));
    InMux I__9996 (
            .O(N__43770),
            .I(N__43761));
    InMux I__9995 (
            .O(N__43767),
            .I(N__43756));
    InMux I__9994 (
            .O(N__43764),
            .I(N__43756));
    LocalMux I__9993 (
            .O(N__43761),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__9992 (
            .O(N__43756),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__9991 (
            .O(N__43751),
            .I(bfn_17_13_0_));
    InMux I__9990 (
            .O(N__43748),
            .I(N__43741));
    InMux I__9989 (
            .O(N__43747),
            .I(N__43741));
    InMux I__9988 (
            .O(N__43746),
            .I(N__43738));
    LocalMux I__9987 (
            .O(N__43741),
            .I(N__43735));
    LocalMux I__9986 (
            .O(N__43738),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv12 I__9985 (
            .O(N__43735),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__9984 (
            .O(N__43730),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ));
    CascadeMux I__9983 (
            .O(N__43727),
            .I(N__43724));
    InMux I__9982 (
            .O(N__43724),
            .I(N__43717));
    InMux I__9981 (
            .O(N__43723),
            .I(N__43717));
    InMux I__9980 (
            .O(N__43722),
            .I(N__43714));
    LocalMux I__9979 (
            .O(N__43717),
            .I(N__43711));
    LocalMux I__9978 (
            .O(N__43714),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv12 I__9977 (
            .O(N__43711),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__9976 (
            .O(N__43706),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ));
    InMux I__9975 (
            .O(N__43703),
            .I(N__43696));
    InMux I__9974 (
            .O(N__43702),
            .I(N__43696));
    InMux I__9973 (
            .O(N__43701),
            .I(N__43693));
    LocalMux I__9972 (
            .O(N__43696),
            .I(N__43690));
    LocalMux I__9971 (
            .O(N__43693),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ));
    Odrv4 I__9970 (
            .O(N__43690),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ));
    InMux I__9969 (
            .O(N__43685),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ));
    CascadeMux I__9968 (
            .O(N__43682),
            .I(N__43678));
    InMux I__9967 (
            .O(N__43681),
            .I(N__43672));
    InMux I__9966 (
            .O(N__43678),
            .I(N__43672));
    InMux I__9965 (
            .O(N__43677),
            .I(N__43669));
    LocalMux I__9964 (
            .O(N__43672),
            .I(N__43666));
    LocalMux I__9963 (
            .O(N__43669),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ));
    Odrv4 I__9962 (
            .O(N__43666),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ));
    InMux I__9961 (
            .O(N__43661),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__9960 (
            .O(N__43658),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ));
    InMux I__9959 (
            .O(N__43655),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ));
    InMux I__9958 (
            .O(N__43652),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ));
    InMux I__9957 (
            .O(N__43649),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__9956 (
            .O(N__43646),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__9955 (
            .O(N__43643),
            .I(bfn_17_12_0_));
    InMux I__9954 (
            .O(N__43640),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__9953 (
            .O(N__43637),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__9952 (
            .O(N__43634),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__9951 (
            .O(N__43631),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__9950 (
            .O(N__43628),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__9949 (
            .O(N__43625),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ));
    InMux I__9948 (
            .O(N__43622),
            .I(N__43619));
    LocalMux I__9947 (
            .O(N__43619),
            .I(N__43614));
    InMux I__9946 (
            .O(N__43618),
            .I(N__43611));
    InMux I__9945 (
            .O(N__43617),
            .I(N__43608));
    Span4Mux_v I__9944 (
            .O(N__43614),
            .I(N__43605));
    LocalMux I__9943 (
            .O(N__43611),
            .I(N__43600));
    LocalMux I__9942 (
            .O(N__43608),
            .I(N__43600));
    Span4Mux_h I__9941 (
            .O(N__43605),
            .I(N__43597));
    Odrv12 I__9940 (
            .O(N__43600),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    Odrv4 I__9939 (
            .O(N__43597),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    InMux I__9938 (
            .O(N__43592),
            .I(N__43589));
    LocalMux I__9937 (
            .O(N__43589),
            .I(N__43585));
    InMux I__9936 (
            .O(N__43588),
            .I(N__43582));
    Span4Mux_v I__9935 (
            .O(N__43585),
            .I(N__43575));
    LocalMux I__9934 (
            .O(N__43582),
            .I(N__43575));
    InMux I__9933 (
            .O(N__43581),
            .I(N__43570));
    InMux I__9932 (
            .O(N__43580),
            .I(N__43570));
    Odrv4 I__9931 (
            .O(N__43575),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    LocalMux I__9930 (
            .O(N__43570),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    InMux I__9929 (
            .O(N__43565),
            .I(N__43561));
    InMux I__9928 (
            .O(N__43564),
            .I(N__43556));
    LocalMux I__9927 (
            .O(N__43561),
            .I(N__43553));
    InMux I__9926 (
            .O(N__43560),
            .I(N__43550));
    CascadeMux I__9925 (
            .O(N__43559),
            .I(N__43547));
    LocalMux I__9924 (
            .O(N__43556),
            .I(N__43544));
    Span4Mux_v I__9923 (
            .O(N__43553),
            .I(N__43539));
    LocalMux I__9922 (
            .O(N__43550),
            .I(N__43539));
    InMux I__9921 (
            .O(N__43547),
            .I(N__43536));
    Span4Mux_h I__9920 (
            .O(N__43544),
            .I(N__43533));
    Span4Mux_v I__9919 (
            .O(N__43539),
            .I(N__43530));
    LocalMux I__9918 (
            .O(N__43536),
            .I(N__43527));
    Odrv4 I__9917 (
            .O(N__43533),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    Odrv4 I__9916 (
            .O(N__43530),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    Odrv12 I__9915 (
            .O(N__43527),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    InMux I__9914 (
            .O(N__43520),
            .I(N__43515));
    InMux I__9913 (
            .O(N__43519),
            .I(N__43512));
    InMux I__9912 (
            .O(N__43518),
            .I(N__43509));
    LocalMux I__9911 (
            .O(N__43515),
            .I(N__43506));
    LocalMux I__9910 (
            .O(N__43512),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    LocalMux I__9909 (
            .O(N__43509),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    Odrv4 I__9908 (
            .O(N__43506),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    InMux I__9907 (
            .O(N__43499),
            .I(N__43494));
    InMux I__9906 (
            .O(N__43498),
            .I(N__43491));
    InMux I__9905 (
            .O(N__43497),
            .I(N__43488));
    LocalMux I__9904 (
            .O(N__43494),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    LocalMux I__9903 (
            .O(N__43491),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    LocalMux I__9902 (
            .O(N__43488),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    InMux I__9901 (
            .O(N__43481),
            .I(N__43477));
    InMux I__9900 (
            .O(N__43480),
            .I(N__43474));
    LocalMux I__9899 (
            .O(N__43477),
            .I(N__43469));
    LocalMux I__9898 (
            .O(N__43474),
            .I(N__43466));
    InMux I__9897 (
            .O(N__43473),
            .I(N__43463));
    InMux I__9896 (
            .O(N__43472),
            .I(N__43460));
    Span4Mux_h I__9895 (
            .O(N__43469),
            .I(N__43457));
    Span4Mux_v I__9894 (
            .O(N__43466),
            .I(N__43454));
    LocalMux I__9893 (
            .O(N__43463),
            .I(N__43449));
    LocalMux I__9892 (
            .O(N__43460),
            .I(N__43449));
    Odrv4 I__9891 (
            .O(N__43457),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    Odrv4 I__9890 (
            .O(N__43454),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    Odrv12 I__9889 (
            .O(N__43449),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    InMux I__9888 (
            .O(N__43442),
            .I(N__43439));
    LocalMux I__9887 (
            .O(N__43439),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ));
    InMux I__9886 (
            .O(N__43436),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ));
    CascadeMux I__9885 (
            .O(N__43433),
            .I(N__43430));
    InMux I__9884 (
            .O(N__43430),
            .I(N__43427));
    LocalMux I__9883 (
            .O(N__43427),
            .I(N__43424));
    Odrv4 I__9882 (
            .O(N__43424),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28 ));
    InMux I__9881 (
            .O(N__43421),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__9880 (
            .O(N__43418),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__9879 (
            .O(N__43415),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ));
    InMux I__9878 (
            .O(N__43412),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__9877 (
            .O(N__43409),
            .I(N__43406));
    LocalMux I__9876 (
            .O(N__43406),
            .I(N__43402));
    InMux I__9875 (
            .O(N__43405),
            .I(N__43398));
    Span4Mux_h I__9874 (
            .O(N__43402),
            .I(N__43395));
    InMux I__9873 (
            .O(N__43401),
            .I(N__43392));
    LocalMux I__9872 (
            .O(N__43398),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    Odrv4 I__9871 (
            .O(N__43395),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    LocalMux I__9870 (
            .O(N__43392),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    InMux I__9869 (
            .O(N__43385),
            .I(N__43380));
    InMux I__9868 (
            .O(N__43384),
            .I(N__43377));
    InMux I__9867 (
            .O(N__43383),
            .I(N__43374));
    LocalMux I__9866 (
            .O(N__43380),
            .I(N__43371));
    LocalMux I__9865 (
            .O(N__43377),
            .I(N__43368));
    LocalMux I__9864 (
            .O(N__43374),
            .I(N__43365));
    Span4Mux_h I__9863 (
            .O(N__43371),
            .I(N__43362));
    Span4Mux_h I__9862 (
            .O(N__43368),
            .I(N__43359));
    Span4Mux_v I__9861 (
            .O(N__43365),
            .I(N__43355));
    Span4Mux_v I__9860 (
            .O(N__43362),
            .I(N__43352));
    Span4Mux_v I__9859 (
            .O(N__43359),
            .I(N__43349));
    InMux I__9858 (
            .O(N__43358),
            .I(N__43346));
    Odrv4 I__9857 (
            .O(N__43355),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    Odrv4 I__9856 (
            .O(N__43352),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    Odrv4 I__9855 (
            .O(N__43349),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    LocalMux I__9854 (
            .O(N__43346),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    InMux I__9853 (
            .O(N__43337),
            .I(N__43334));
    LocalMux I__9852 (
            .O(N__43334),
            .I(N__43330));
    InMux I__9851 (
            .O(N__43333),
            .I(N__43327));
    Odrv4 I__9850 (
            .O(N__43330),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    LocalMux I__9849 (
            .O(N__43327),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    CascadeMux I__9848 (
            .O(N__43322),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18_cascade_));
    InMux I__9847 (
            .O(N__43319),
            .I(N__43312));
    InMux I__9846 (
            .O(N__43318),
            .I(N__43312));
    InMux I__9845 (
            .O(N__43317),
            .I(N__43309));
    LocalMux I__9844 (
            .O(N__43312),
            .I(N__43306));
    LocalMux I__9843 (
            .O(N__43309),
            .I(N__43303));
    Span4Mux_h I__9842 (
            .O(N__43306),
            .I(N__43300));
    Span12Mux_v I__9841 (
            .O(N__43303),
            .I(N__43296));
    Span4Mux_v I__9840 (
            .O(N__43300),
            .I(N__43293));
    InMux I__9839 (
            .O(N__43299),
            .I(N__43290));
    Odrv12 I__9838 (
            .O(N__43296),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    Odrv4 I__9837 (
            .O(N__43293),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    LocalMux I__9836 (
            .O(N__43290),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    InMux I__9835 (
            .O(N__43283),
            .I(N__43277));
    InMux I__9834 (
            .O(N__43282),
            .I(N__43277));
    LocalMux I__9833 (
            .O(N__43277),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    InMux I__9832 (
            .O(N__43274),
            .I(N__43269));
    InMux I__9831 (
            .O(N__43273),
            .I(N__43266));
    InMux I__9830 (
            .O(N__43272),
            .I(N__43263));
    LocalMux I__9829 (
            .O(N__43269),
            .I(N__43260));
    LocalMux I__9828 (
            .O(N__43266),
            .I(N__43257));
    LocalMux I__9827 (
            .O(N__43263),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20));
    Odrv4 I__9826 (
            .O(N__43260),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20));
    Odrv4 I__9825 (
            .O(N__43257),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20));
    InMux I__9824 (
            .O(N__43250),
            .I(N__43246));
    InMux I__9823 (
            .O(N__43249),
            .I(N__43242));
    LocalMux I__9822 (
            .O(N__43246),
            .I(N__43239));
    InMux I__9821 (
            .O(N__43245),
            .I(N__43236));
    LocalMux I__9820 (
            .O(N__43242),
            .I(N__43233));
    Span4Mux_h I__9819 (
            .O(N__43239),
            .I(N__43229));
    LocalMux I__9818 (
            .O(N__43236),
            .I(N__43224));
    Span4Mux_h I__9817 (
            .O(N__43233),
            .I(N__43224));
    CascadeMux I__9816 (
            .O(N__43232),
            .I(N__43221));
    Span4Mux_v I__9815 (
            .O(N__43229),
            .I(N__43218));
    Span4Mux_v I__9814 (
            .O(N__43224),
            .I(N__43215));
    InMux I__9813 (
            .O(N__43221),
            .I(N__43212));
    Odrv4 I__9812 (
            .O(N__43218),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    Odrv4 I__9811 (
            .O(N__43215),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    LocalMux I__9810 (
            .O(N__43212),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__9809 (
            .O(N__43205),
            .I(N__43199));
    InMux I__9808 (
            .O(N__43204),
            .I(N__43199));
    LocalMux I__9807 (
            .O(N__43199),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ));
    CascadeMux I__9806 (
            .O(N__43196),
            .I(N__43193));
    InMux I__9805 (
            .O(N__43193),
            .I(N__43187));
    InMux I__9804 (
            .O(N__43192),
            .I(N__43187));
    LocalMux I__9803 (
            .O(N__43187),
            .I(N__43184));
    Span4Mux_v I__9802 (
            .O(N__43184),
            .I(N__43181));
    Odrv4 I__9801 (
            .O(N__43181),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ));
    InMux I__9800 (
            .O(N__43178),
            .I(N__43174));
    InMux I__9799 (
            .O(N__43177),
            .I(N__43170));
    LocalMux I__9798 (
            .O(N__43174),
            .I(N__43167));
    InMux I__9797 (
            .O(N__43173),
            .I(N__43164));
    LocalMux I__9796 (
            .O(N__43170),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    Odrv4 I__9795 (
            .O(N__43167),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    LocalMux I__9794 (
            .O(N__43164),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    InMux I__9793 (
            .O(N__43157),
            .I(N__43152));
    InMux I__9792 (
            .O(N__43156),
            .I(N__43149));
    InMux I__9791 (
            .O(N__43155),
            .I(N__43146));
    LocalMux I__9790 (
            .O(N__43152),
            .I(N__43142));
    LocalMux I__9789 (
            .O(N__43149),
            .I(N__43139));
    LocalMux I__9788 (
            .O(N__43146),
            .I(N__43136));
    InMux I__9787 (
            .O(N__43145),
            .I(N__43133));
    Odrv4 I__9786 (
            .O(N__43142),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    Odrv4 I__9785 (
            .O(N__43139),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    Odrv4 I__9784 (
            .O(N__43136),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    LocalMux I__9783 (
            .O(N__43133),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    InMux I__9782 (
            .O(N__43124),
            .I(N__43118));
    InMux I__9781 (
            .O(N__43123),
            .I(N__43118));
    LocalMux I__9780 (
            .O(N__43118),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    CascadeMux I__9779 (
            .O(N__43115),
            .I(N__43112));
    InMux I__9778 (
            .O(N__43112),
            .I(N__43106));
    InMux I__9777 (
            .O(N__43111),
            .I(N__43106));
    LocalMux I__9776 (
            .O(N__43106),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    CascadeMux I__9775 (
            .O(N__43103),
            .I(N__43100));
    InMux I__9774 (
            .O(N__43100),
            .I(N__43097));
    LocalMux I__9773 (
            .O(N__43097),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ));
    CascadeMux I__9772 (
            .O(N__43094),
            .I(N__43090));
    InMux I__9771 (
            .O(N__43093),
            .I(N__43087));
    InMux I__9770 (
            .O(N__43090),
            .I(N__43084));
    LocalMux I__9769 (
            .O(N__43087),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    LocalMux I__9768 (
            .O(N__43084),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    InMux I__9767 (
            .O(N__43079),
            .I(N__43076));
    LocalMux I__9766 (
            .O(N__43076),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ));
    InMux I__9765 (
            .O(N__43073),
            .I(N__43070));
    LocalMux I__9764 (
            .O(N__43070),
            .I(N__43064));
    InMux I__9763 (
            .O(N__43069),
            .I(N__43061));
    InMux I__9762 (
            .O(N__43068),
            .I(N__43058));
    InMux I__9761 (
            .O(N__43067),
            .I(N__43054));
    Span12Mux_s2_v I__9760 (
            .O(N__43064),
            .I(N__43047));
    LocalMux I__9759 (
            .O(N__43061),
            .I(N__43047));
    LocalMux I__9758 (
            .O(N__43058),
            .I(N__43047));
    InMux I__9757 (
            .O(N__43057),
            .I(N__43044));
    LocalMux I__9756 (
            .O(N__43054),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv12 I__9755 (
            .O(N__43047),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__9754 (
            .O(N__43044),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    IoInMux I__9753 (
            .O(N__43037),
            .I(N__43034));
    LocalMux I__9752 (
            .O(N__43034),
            .I(N__43031));
    IoSpan4Mux I__9751 (
            .O(N__43031),
            .I(N__43028));
    Odrv4 I__9750 (
            .O(N__43028),
            .I(s2_phy_c));
    InMux I__9749 (
            .O(N__43025),
            .I(N__43021));
    InMux I__9748 (
            .O(N__43024),
            .I(N__43018));
    LocalMux I__9747 (
            .O(N__43021),
            .I(N__43013));
    LocalMux I__9746 (
            .O(N__43018),
            .I(N__43013));
    Span4Mux_s3_v I__9745 (
            .O(N__43013),
            .I(N__43010));
    Sp12to4 I__9744 (
            .O(N__43010),
            .I(N__43007));
    Span12Mux_s6_h I__9743 (
            .O(N__43007),
            .I(N__43003));
    InMux I__9742 (
            .O(N__43006),
            .I(N__43000));
    Span12Mux_v I__9741 (
            .O(N__43003),
            .I(N__42996));
    LocalMux I__9740 (
            .O(N__43000),
            .I(N__42993));
    InMux I__9739 (
            .O(N__42999),
            .I(N__42990));
    Span12Mux_v I__9738 (
            .O(N__42996),
            .I(N__42987));
    Span4Mux_v I__9737 (
            .O(N__42993),
            .I(N__42984));
    LocalMux I__9736 (
            .O(N__42990),
            .I(N__42981));
    Span12Mux_h I__9735 (
            .O(N__42987),
            .I(N__42978));
    Span4Mux_h I__9734 (
            .O(N__42984),
            .I(N__42973));
    Span4Mux_v I__9733 (
            .O(N__42981),
            .I(N__42973));
    Odrv12 I__9732 (
            .O(N__42978),
            .I(start_stop_c));
    Odrv4 I__9731 (
            .O(N__42973),
            .I(start_stop_c));
    CascadeMux I__9730 (
            .O(N__42968),
            .I(N__42963));
    InMux I__9729 (
            .O(N__42967),
            .I(N__42959));
    InMux I__9728 (
            .O(N__42966),
            .I(N__42956));
    InMux I__9727 (
            .O(N__42963),
            .I(N__42953));
    InMux I__9726 (
            .O(N__42962),
            .I(N__42950));
    LocalMux I__9725 (
            .O(N__42959),
            .I(N__42947));
    LocalMux I__9724 (
            .O(N__42956),
            .I(N__42942));
    LocalMux I__9723 (
            .O(N__42953),
            .I(N__42942));
    LocalMux I__9722 (
            .O(N__42950),
            .I(N__42936));
    Span4Mux_h I__9721 (
            .O(N__42947),
            .I(N__42936));
    Span4Mux_v I__9720 (
            .O(N__42942),
            .I(N__42933));
    InMux I__9719 (
            .O(N__42941),
            .I(N__42930));
    Span4Mux_v I__9718 (
            .O(N__42936),
            .I(N__42926));
    Span4Mux_v I__9717 (
            .O(N__42933),
            .I(N__42921));
    LocalMux I__9716 (
            .O(N__42930),
            .I(N__42921));
    InMux I__9715 (
            .O(N__42929),
            .I(N__42918));
    Span4Mux_v I__9714 (
            .O(N__42926),
            .I(N__42913));
    Span4Mux_h I__9713 (
            .O(N__42921),
            .I(N__42913));
    LocalMux I__9712 (
            .O(N__42918),
            .I(phase_controller_inst1_state_4));
    Odrv4 I__9711 (
            .O(N__42913),
            .I(phase_controller_inst1_state_4));
    CascadeMux I__9710 (
            .O(N__42908),
            .I(N__42904));
    InMux I__9709 (
            .O(N__42907),
            .I(N__42901));
    InMux I__9708 (
            .O(N__42904),
            .I(N__42898));
    LocalMux I__9707 (
            .O(N__42901),
            .I(N__42895));
    LocalMux I__9706 (
            .O(N__42898),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    Odrv12 I__9705 (
            .O(N__42895),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    InMux I__9704 (
            .O(N__42890),
            .I(N__42884));
    InMux I__9703 (
            .O(N__42889),
            .I(N__42884));
    LocalMux I__9702 (
            .O(N__42884),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    InMux I__9701 (
            .O(N__42881),
            .I(N__42875));
    InMux I__9700 (
            .O(N__42880),
            .I(N__42875));
    LocalMux I__9699 (
            .O(N__42875),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    CascadeMux I__9698 (
            .O(N__42872),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ));
    InMux I__9697 (
            .O(N__42869),
            .I(N__42863));
    InMux I__9696 (
            .O(N__42868),
            .I(N__42863));
    LocalMux I__9695 (
            .O(N__42863),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    InMux I__9694 (
            .O(N__42860),
            .I(N__42854));
    InMux I__9693 (
            .O(N__42859),
            .I(N__42854));
    LocalMux I__9692 (
            .O(N__42854),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    InMux I__9691 (
            .O(N__42851),
            .I(N__42845));
    InMux I__9690 (
            .O(N__42850),
            .I(N__42845));
    LocalMux I__9689 (
            .O(N__42845),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    InMux I__9688 (
            .O(N__42842),
            .I(N__42836));
    InMux I__9687 (
            .O(N__42841),
            .I(N__42836));
    LocalMux I__9686 (
            .O(N__42836),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    InMux I__9685 (
            .O(N__42833),
            .I(N__42827));
    InMux I__9684 (
            .O(N__42832),
            .I(N__42827));
    LocalMux I__9683 (
            .O(N__42827),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    InMux I__9682 (
            .O(N__42824),
            .I(N__42820));
    InMux I__9681 (
            .O(N__42823),
            .I(N__42817));
    LocalMux I__9680 (
            .O(N__42820),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    LocalMux I__9679 (
            .O(N__42817),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    CascadeMux I__9678 (
            .O(N__42812),
            .I(N__42809));
    InMux I__9677 (
            .O(N__42809),
            .I(N__42805));
    InMux I__9676 (
            .O(N__42808),
            .I(N__42802));
    LocalMux I__9675 (
            .O(N__42805),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    LocalMux I__9674 (
            .O(N__42802),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    CascadeMux I__9673 (
            .O(N__42797),
            .I(N__42794));
    InMux I__9672 (
            .O(N__42794),
            .I(N__42791));
    LocalMux I__9671 (
            .O(N__42791),
            .I(N__42787));
    InMux I__9670 (
            .O(N__42790),
            .I(N__42784));
    Odrv4 I__9669 (
            .O(N__42787),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    LocalMux I__9668 (
            .O(N__42784),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    InMux I__9667 (
            .O(N__42779),
            .I(N__42776));
    LocalMux I__9666 (
            .O(N__42776),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ));
    InMux I__9665 (
            .O(N__42773),
            .I(N__42769));
    InMux I__9664 (
            .O(N__42772),
            .I(N__42766));
    LocalMux I__9663 (
            .O(N__42769),
            .I(N__42763));
    LocalMux I__9662 (
            .O(N__42766),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    Odrv4 I__9661 (
            .O(N__42763),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    CascadeMux I__9660 (
            .O(N__42758),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_ ));
    CascadeMux I__9659 (
            .O(N__42755),
            .I(N__42751));
    InMux I__9658 (
            .O(N__42754),
            .I(N__42748));
    InMux I__9657 (
            .O(N__42751),
            .I(N__42745));
    LocalMux I__9656 (
            .O(N__42748),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    LocalMux I__9655 (
            .O(N__42745),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    InMux I__9654 (
            .O(N__42740),
            .I(N__42734));
    InMux I__9653 (
            .O(N__42739),
            .I(N__42734));
    LocalMux I__9652 (
            .O(N__42734),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    InMux I__9651 (
            .O(N__42731),
            .I(N__42725));
    InMux I__9650 (
            .O(N__42730),
            .I(N__42725));
    LocalMux I__9649 (
            .O(N__42725),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    ClkMux I__9648 (
            .O(N__42722),
            .I(N__42716));
    ClkMux I__9647 (
            .O(N__42721),
            .I(N__42716));
    GlobalMux I__9646 (
            .O(N__42716),
            .I(N__42713));
    gio2CtrlBuf I__9645 (
            .O(N__42713),
            .I(delay_tr_input_c_g));
    CascadeMux I__9644 (
            .O(N__42710),
            .I(N__42705));
    InMux I__9643 (
            .O(N__42709),
            .I(N__42700));
    InMux I__9642 (
            .O(N__42708),
            .I(N__42700));
    InMux I__9641 (
            .O(N__42705),
            .I(N__42696));
    LocalMux I__9640 (
            .O(N__42700),
            .I(N__42693));
    InMux I__9639 (
            .O(N__42699),
            .I(N__42690));
    LocalMux I__9638 (
            .O(N__42696),
            .I(N__42687));
    Span4Mux_v I__9637 (
            .O(N__42693),
            .I(N__42684));
    LocalMux I__9636 (
            .O(N__42690),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv4 I__9635 (
            .O(N__42687),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv4 I__9634 (
            .O(N__42684),
            .I(\phase_controller_inst1.hc_time_passed ));
    InMux I__9633 (
            .O(N__42677),
            .I(N__42674));
    LocalMux I__9632 (
            .O(N__42674),
            .I(N__42671));
    Odrv4 I__9631 (
            .O(N__42671),
            .I(\phase_controller_inst1.start_timer_tr_RNOZ0Z_0 ));
    InMux I__9630 (
            .O(N__42668),
            .I(N__42664));
    InMux I__9629 (
            .O(N__42667),
            .I(N__42661));
    LocalMux I__9628 (
            .O(N__42664),
            .I(\phase_controller_inst1.state_RNIE87FZ0Z_2 ));
    LocalMux I__9627 (
            .O(N__42661),
            .I(\phase_controller_inst1.state_RNIE87FZ0Z_2 ));
    IoInMux I__9626 (
            .O(N__42656),
            .I(N__42653));
    LocalMux I__9625 (
            .O(N__42653),
            .I(N__42649));
    InMux I__9624 (
            .O(N__42652),
            .I(N__42646));
    Odrv12 I__9623 (
            .O(N__42649),
            .I(T45_c));
    LocalMux I__9622 (
            .O(N__42646),
            .I(T45_c));
    CascadeMux I__9621 (
            .O(N__42641),
            .I(N__42638));
    InMux I__9620 (
            .O(N__42638),
            .I(N__42635));
    LocalMux I__9619 (
            .O(N__42635),
            .I(N__42630));
    InMux I__9618 (
            .O(N__42634),
            .I(N__42627));
    InMux I__9617 (
            .O(N__42633),
            .I(N__42624));
    Span4Mux_v I__9616 (
            .O(N__42630),
            .I(N__42619));
    LocalMux I__9615 (
            .O(N__42627),
            .I(N__42619));
    LocalMux I__9614 (
            .O(N__42624),
            .I(N__42616));
    Span4Mux_v I__9613 (
            .O(N__42619),
            .I(N__42613));
    Span4Mux_h I__9612 (
            .O(N__42616),
            .I(N__42610));
    Span4Mux_h I__9611 (
            .O(N__42613),
            .I(N__42607));
    Span4Mux_h I__9610 (
            .O(N__42610),
            .I(N__42604));
    Span4Mux_v I__9609 (
            .O(N__42607),
            .I(N__42601));
    Span4Mux_v I__9608 (
            .O(N__42604),
            .I(N__42598));
    Odrv4 I__9607 (
            .O(N__42601),
            .I(il_min_comp1_D2));
    Odrv4 I__9606 (
            .O(N__42598),
            .I(il_min_comp1_D2));
    IoInMux I__9605 (
            .O(N__42593),
            .I(N__42590));
    LocalMux I__9604 (
            .O(N__42590),
            .I(N__42587));
    Span12Mux_s7_v I__9603 (
            .O(N__42587),
            .I(N__42583));
    InMux I__9602 (
            .O(N__42586),
            .I(N__42580));
    Odrv12 I__9601 (
            .O(N__42583),
            .I(T23_c));
    LocalMux I__9600 (
            .O(N__42580),
            .I(T23_c));
    InMux I__9599 (
            .O(N__42575),
            .I(N__42572));
    LocalMux I__9598 (
            .O(N__42572),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ));
    CascadeMux I__9597 (
            .O(N__42569),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18_cascade_ ));
    InMux I__9596 (
            .O(N__42566),
            .I(N__42563));
    LocalMux I__9595 (
            .O(N__42563),
            .I(N__42560));
    Span4Mux_h I__9594 (
            .O(N__42560),
            .I(N__42557));
    Odrv4 I__9593 (
            .O(N__42557),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ));
    InMux I__9592 (
            .O(N__42554),
            .I(N__42549));
    InMux I__9591 (
            .O(N__42553),
            .I(N__42546));
    InMux I__9590 (
            .O(N__42552),
            .I(N__42543));
    LocalMux I__9589 (
            .O(N__42549),
            .I(N__42540));
    LocalMux I__9588 (
            .O(N__42546),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    LocalMux I__9587 (
            .O(N__42543),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    Odrv12 I__9586 (
            .O(N__42540),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    InMux I__9585 (
            .O(N__42533),
            .I(N__42530));
    LocalMux I__9584 (
            .O(N__42530),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ));
    InMux I__9583 (
            .O(N__42527),
            .I(N__42524));
    LocalMux I__9582 (
            .O(N__42524),
            .I(N__42519));
    InMux I__9581 (
            .O(N__42523),
            .I(N__42516));
    InMux I__9580 (
            .O(N__42522),
            .I(N__42513));
    Span4Mux_h I__9579 (
            .O(N__42519),
            .I(N__42507));
    LocalMux I__9578 (
            .O(N__42516),
            .I(N__42507));
    LocalMux I__9577 (
            .O(N__42513),
            .I(N__42504));
    InMux I__9576 (
            .O(N__42512),
            .I(N__42501));
    Odrv4 I__9575 (
            .O(N__42507),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    Odrv4 I__9574 (
            .O(N__42504),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    LocalMux I__9573 (
            .O(N__42501),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    InMux I__9572 (
            .O(N__42494),
            .I(N__42491));
    LocalMux I__9571 (
            .O(N__42491),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ));
    InMux I__9570 (
            .O(N__42488),
            .I(N__42483));
    InMux I__9569 (
            .O(N__42487),
            .I(N__42480));
    InMux I__9568 (
            .O(N__42486),
            .I(N__42477));
    LocalMux I__9567 (
            .O(N__42483),
            .I(N__42474));
    LocalMux I__9566 (
            .O(N__42480),
            .I(N__42470));
    LocalMux I__9565 (
            .O(N__42477),
            .I(N__42465));
    Span4Mux_h I__9564 (
            .O(N__42474),
            .I(N__42465));
    InMux I__9563 (
            .O(N__42473),
            .I(N__42462));
    Odrv12 I__9562 (
            .O(N__42470),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    Odrv4 I__9561 (
            .O(N__42465),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    LocalMux I__9560 (
            .O(N__42462),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    InMux I__9559 (
            .O(N__42455),
            .I(N__42452));
    LocalMux I__9558 (
            .O(N__42452),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ));
    InMux I__9557 (
            .O(N__42449),
            .I(N__42446));
    LocalMux I__9556 (
            .O(N__42446),
            .I(N__42442));
    InMux I__9555 (
            .O(N__42445),
            .I(N__42438));
    Span4Mux_h I__9554 (
            .O(N__42442),
            .I(N__42435));
    InMux I__9553 (
            .O(N__42441),
            .I(N__42432));
    LocalMux I__9552 (
            .O(N__42438),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    Odrv4 I__9551 (
            .O(N__42435),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    LocalMux I__9550 (
            .O(N__42432),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    InMux I__9549 (
            .O(N__42425),
            .I(N__42422));
    LocalMux I__9548 (
            .O(N__42422),
            .I(N__42419));
    Span4Mux_h I__9547 (
            .O(N__42419),
            .I(N__42414));
    InMux I__9546 (
            .O(N__42418),
            .I(N__42408));
    InMux I__9545 (
            .O(N__42417),
            .I(N__42408));
    Span4Mux_v I__9544 (
            .O(N__42414),
            .I(N__42405));
    InMux I__9543 (
            .O(N__42413),
            .I(N__42402));
    LocalMux I__9542 (
            .O(N__42408),
            .I(N__42399));
    Odrv4 I__9541 (
            .O(N__42405),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    LocalMux I__9540 (
            .O(N__42402),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    Odrv4 I__9539 (
            .O(N__42399),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__9538 (
            .O(N__42392),
            .I(N__42389));
    LocalMux I__9537 (
            .O(N__42389),
            .I(N__42385));
    CascadeMux I__9536 (
            .O(N__42388),
            .I(N__42381));
    Sp12to4 I__9535 (
            .O(N__42385),
            .I(N__42377));
    InMux I__9534 (
            .O(N__42384),
            .I(N__42374));
    InMux I__9533 (
            .O(N__42381),
            .I(N__42371));
    InMux I__9532 (
            .O(N__42380),
            .I(N__42368));
    Span12Mux_s11_v I__9531 (
            .O(N__42377),
            .I(N__42365));
    LocalMux I__9530 (
            .O(N__42374),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    LocalMux I__9529 (
            .O(N__42371),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    LocalMux I__9528 (
            .O(N__42368),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv12 I__9527 (
            .O(N__42365),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    InMux I__9526 (
            .O(N__42356),
            .I(N__42352));
    InMux I__9525 (
            .O(N__42355),
            .I(N__42349));
    LocalMux I__9524 (
            .O(N__42352),
            .I(N__42345));
    LocalMux I__9523 (
            .O(N__42349),
            .I(N__42341));
    InMux I__9522 (
            .O(N__42348),
            .I(N__42337));
    Span4Mux_h I__9521 (
            .O(N__42345),
            .I(N__42334));
    InMux I__9520 (
            .O(N__42344),
            .I(N__42331));
    Span4Mux_v I__9519 (
            .O(N__42341),
            .I(N__42328));
    CascadeMux I__9518 (
            .O(N__42340),
            .I(N__42325));
    LocalMux I__9517 (
            .O(N__42337),
            .I(N__42322));
    Span4Mux_v I__9516 (
            .O(N__42334),
            .I(N__42319));
    LocalMux I__9515 (
            .O(N__42331),
            .I(N__42316));
    Span4Mux_v I__9514 (
            .O(N__42328),
            .I(N__42313));
    InMux I__9513 (
            .O(N__42325),
            .I(N__42310));
    Span12Mux_h I__9512 (
            .O(N__42322),
            .I(N__42307));
    Span4Mux_v I__9511 (
            .O(N__42319),
            .I(N__42302));
    Span4Mux_h I__9510 (
            .O(N__42316),
            .I(N__42302));
    Span4Mux_h I__9509 (
            .O(N__42313),
            .I(N__42299));
    LocalMux I__9508 (
            .O(N__42310),
            .I(N__42294));
    Span12Mux_v I__9507 (
            .O(N__42307),
            .I(N__42294));
    Odrv4 I__9506 (
            .O(N__42302),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    Odrv4 I__9505 (
            .O(N__42299),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    Odrv12 I__9504 (
            .O(N__42294),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    CascadeMux I__9503 (
            .O(N__42287),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ));
    InMux I__9502 (
            .O(N__42284),
            .I(N__42281));
    LocalMux I__9501 (
            .O(N__42281),
            .I(N__42278));
    Span4Mux_h I__9500 (
            .O(N__42278),
            .I(N__42274));
    InMux I__9499 (
            .O(N__42277),
            .I(N__42271));
    Odrv4 I__9498 (
            .O(N__42274),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    LocalMux I__9497 (
            .O(N__42271),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    InMux I__9496 (
            .O(N__42266),
            .I(N__42263));
    LocalMux I__9495 (
            .O(N__42263),
            .I(N__42259));
    InMux I__9494 (
            .O(N__42262),
            .I(N__42255));
    Span4Mux_h I__9493 (
            .O(N__42259),
            .I(N__42252));
    InMux I__9492 (
            .O(N__42258),
            .I(N__42249));
    LocalMux I__9491 (
            .O(N__42255),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    Odrv4 I__9490 (
            .O(N__42252),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    LocalMux I__9489 (
            .O(N__42249),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    InMux I__9488 (
            .O(N__42242),
            .I(N__42236));
    InMux I__9487 (
            .O(N__42241),
            .I(N__42236));
    LocalMux I__9486 (
            .O(N__42236),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ));
    InMux I__9485 (
            .O(N__42233),
            .I(N__42227));
    InMux I__9484 (
            .O(N__42232),
            .I(N__42227));
    LocalMux I__9483 (
            .O(N__42227),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    InMux I__9482 (
            .O(N__42224),
            .I(N__42221));
    LocalMux I__9481 (
            .O(N__42221),
            .I(N__42217));
    InMux I__9480 (
            .O(N__42220),
            .I(N__42213));
    Span4Mux_h I__9479 (
            .O(N__42217),
            .I(N__42210));
    InMux I__9478 (
            .O(N__42216),
            .I(N__42207));
    LocalMux I__9477 (
            .O(N__42213),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    Odrv4 I__9476 (
            .O(N__42210),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    LocalMux I__9475 (
            .O(N__42207),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    InMux I__9474 (
            .O(N__42200),
            .I(N__42194));
    InMux I__9473 (
            .O(N__42199),
            .I(N__42194));
    LocalMux I__9472 (
            .O(N__42194),
            .I(N__42189));
    InMux I__9471 (
            .O(N__42193),
            .I(N__42186));
    InMux I__9470 (
            .O(N__42192),
            .I(N__42183));
    Span4Mux_h I__9469 (
            .O(N__42189),
            .I(N__42180));
    LocalMux I__9468 (
            .O(N__42186),
            .I(N__42175));
    LocalMux I__9467 (
            .O(N__42183),
            .I(N__42175));
    Odrv4 I__9466 (
            .O(N__42180),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    Odrv4 I__9465 (
            .O(N__42175),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    InMux I__9464 (
            .O(N__42170),
            .I(N__42166));
    InMux I__9463 (
            .O(N__42169),
            .I(N__42161));
    LocalMux I__9462 (
            .O(N__42166),
            .I(N__42158));
    InMux I__9461 (
            .O(N__42165),
            .I(N__42155));
    CascadeMux I__9460 (
            .O(N__42164),
            .I(N__42152));
    LocalMux I__9459 (
            .O(N__42161),
            .I(N__42145));
    Span4Mux_h I__9458 (
            .O(N__42158),
            .I(N__42145));
    LocalMux I__9457 (
            .O(N__42155),
            .I(N__42145));
    InMux I__9456 (
            .O(N__42152),
            .I(N__42142));
    Odrv4 I__9455 (
            .O(N__42145),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    LocalMux I__9454 (
            .O(N__42142),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    CascadeMux I__9453 (
            .O(N__42137),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_ ));
    CascadeMux I__9452 (
            .O(N__42134),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ));
    InMux I__9451 (
            .O(N__42131),
            .I(N__42128));
    LocalMux I__9450 (
            .O(N__42128),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ));
    CascadeMux I__9449 (
            .O(N__42125),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ));
    InMux I__9448 (
            .O(N__42122),
            .I(N__42119));
    LocalMux I__9447 (
            .O(N__42119),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ));
    InMux I__9446 (
            .O(N__42116),
            .I(N__42112));
    InMux I__9445 (
            .O(N__42115),
            .I(N__42109));
    LocalMux I__9444 (
            .O(N__42112),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    LocalMux I__9443 (
            .O(N__42109),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    InMux I__9442 (
            .O(N__42104),
            .I(N__42098));
    InMux I__9441 (
            .O(N__42103),
            .I(N__42091));
    InMux I__9440 (
            .O(N__42102),
            .I(N__42091));
    InMux I__9439 (
            .O(N__42101),
            .I(N__42091));
    LocalMux I__9438 (
            .O(N__42098),
            .I(N__42086));
    LocalMux I__9437 (
            .O(N__42091),
            .I(N__42086));
    Span4Mux_h I__9436 (
            .O(N__42086),
            .I(N__42083));
    Odrv4 I__9435 (
            .O(N__42083),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    CascadeMux I__9434 (
            .O(N__42080),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10_cascade_));
    CascadeMux I__9433 (
            .O(N__42077),
            .I(N__42073));
    InMux I__9432 (
            .O(N__42076),
            .I(N__42066));
    InMux I__9431 (
            .O(N__42073),
            .I(N__42066));
    InMux I__9430 (
            .O(N__42072),
            .I(N__42061));
    InMux I__9429 (
            .O(N__42071),
            .I(N__42061));
    LocalMux I__9428 (
            .O(N__42066),
            .I(N__42058));
    LocalMux I__9427 (
            .O(N__42061),
            .I(N__42053));
    Span4Mux_h I__9426 (
            .O(N__42058),
            .I(N__42053));
    Odrv4 I__9425 (
            .O(N__42053),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    InMux I__9424 (
            .O(N__42050),
            .I(N__42046));
    InMux I__9423 (
            .O(N__42049),
            .I(N__42043));
    LocalMux I__9422 (
            .O(N__42046),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    LocalMux I__9421 (
            .O(N__42043),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    CascadeMux I__9420 (
            .O(N__42038),
            .I(N__42035));
    InMux I__9419 (
            .O(N__42035),
            .I(N__42032));
    LocalMux I__9418 (
            .O(N__42032),
            .I(N__42029));
    Odrv4 I__9417 (
            .O(N__42029),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt26 ));
    InMux I__9416 (
            .O(N__42026),
            .I(N__42020));
    InMux I__9415 (
            .O(N__42025),
            .I(N__42020));
    LocalMux I__9414 (
            .O(N__42020),
            .I(N__42016));
    InMux I__9413 (
            .O(N__42019),
            .I(N__42013));
    Span4Mux_h I__9412 (
            .O(N__42016),
            .I(N__42010));
    LocalMux I__9411 (
            .O(N__42013),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ));
    Odrv4 I__9410 (
            .O(N__42010),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ));
    CascadeMux I__9409 (
            .O(N__42005),
            .I(N__42001));
    CascadeMux I__9408 (
            .O(N__42004),
            .I(N__41998));
    InMux I__9407 (
            .O(N__42001),
            .I(N__41995));
    InMux I__9406 (
            .O(N__41998),
            .I(N__41992));
    LocalMux I__9405 (
            .O(N__41995),
            .I(N__41987));
    LocalMux I__9404 (
            .O(N__41992),
            .I(N__41987));
    Span4Mux_h I__9403 (
            .O(N__41987),
            .I(N__41983));
    InMux I__9402 (
            .O(N__41986),
            .I(N__41980));
    Span4Mux_h I__9401 (
            .O(N__41983),
            .I(N__41977));
    LocalMux I__9400 (
            .O(N__41980),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ));
    Odrv4 I__9399 (
            .O(N__41977),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ));
    InMux I__9398 (
            .O(N__41972),
            .I(N__41968));
    InMux I__9397 (
            .O(N__41971),
            .I(N__41965));
    LocalMux I__9396 (
            .O(N__41968),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ));
    LocalMux I__9395 (
            .O(N__41965),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ));
    InMux I__9394 (
            .O(N__41960),
            .I(N__41957));
    LocalMux I__9393 (
            .O(N__41957),
            .I(N__41954));
    Odrv4 I__9392 (
            .O(N__41954),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ));
    InMux I__9391 (
            .O(N__41951),
            .I(N__41948));
    LocalMux I__9390 (
            .O(N__41948),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15 ));
    InMux I__9389 (
            .O(N__41945),
            .I(N__41939));
    InMux I__9388 (
            .O(N__41944),
            .I(N__41936));
    CascadeMux I__9387 (
            .O(N__41943),
            .I(N__41933));
    InMux I__9386 (
            .O(N__41942),
            .I(N__41930));
    LocalMux I__9385 (
            .O(N__41939),
            .I(N__41927));
    LocalMux I__9384 (
            .O(N__41936),
            .I(N__41924));
    InMux I__9383 (
            .O(N__41933),
            .I(N__41921));
    LocalMux I__9382 (
            .O(N__41930),
            .I(N__41914));
    Span4Mux_v I__9381 (
            .O(N__41927),
            .I(N__41914));
    Span4Mux_h I__9380 (
            .O(N__41924),
            .I(N__41914));
    LocalMux I__9379 (
            .O(N__41921),
            .I(N__41911));
    Span4Mux_h I__9378 (
            .O(N__41914),
            .I(N__41906));
    Span4Mux_v I__9377 (
            .O(N__41911),
            .I(N__41906));
    Odrv4 I__9376 (
            .O(N__41906),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    InMux I__9375 (
            .O(N__41903),
            .I(N__41875));
    InMux I__9374 (
            .O(N__41902),
            .I(N__41868));
    InMux I__9373 (
            .O(N__41901),
            .I(N__41868));
    InMux I__9372 (
            .O(N__41900),
            .I(N__41868));
    InMux I__9371 (
            .O(N__41899),
            .I(N__41865));
    InMux I__9370 (
            .O(N__41898),
            .I(N__41862));
    InMux I__9369 (
            .O(N__41897),
            .I(N__41844));
    InMux I__9368 (
            .O(N__41896),
            .I(N__41844));
    InMux I__9367 (
            .O(N__41895),
            .I(N__41841));
    InMux I__9366 (
            .O(N__41894),
            .I(N__41834));
    InMux I__9365 (
            .O(N__41893),
            .I(N__41834));
    InMux I__9364 (
            .O(N__41892),
            .I(N__41834));
    InMux I__9363 (
            .O(N__41891),
            .I(N__41829));
    InMux I__9362 (
            .O(N__41890),
            .I(N__41826));
    InMux I__9361 (
            .O(N__41889),
            .I(N__41822));
    InMux I__9360 (
            .O(N__41888),
            .I(N__41817));
    InMux I__9359 (
            .O(N__41887),
            .I(N__41811));
    InMux I__9358 (
            .O(N__41886),
            .I(N__41806));
    InMux I__9357 (
            .O(N__41885),
            .I(N__41806));
    InMux I__9356 (
            .O(N__41884),
            .I(N__41803));
    InMux I__9355 (
            .O(N__41883),
            .I(N__41796));
    InMux I__9354 (
            .O(N__41882),
            .I(N__41796));
    InMux I__9353 (
            .O(N__41881),
            .I(N__41796));
    InMux I__9352 (
            .O(N__41880),
            .I(N__41776));
    InMux I__9351 (
            .O(N__41879),
            .I(N__41765));
    InMux I__9350 (
            .O(N__41878),
            .I(N__41762));
    LocalMux I__9349 (
            .O(N__41875),
            .I(N__41757));
    LocalMux I__9348 (
            .O(N__41868),
            .I(N__41757));
    LocalMux I__9347 (
            .O(N__41865),
            .I(N__41752));
    LocalMux I__9346 (
            .O(N__41862),
            .I(N__41752));
    InMux I__9345 (
            .O(N__41861),
            .I(N__41749));
    InMux I__9344 (
            .O(N__41860),
            .I(N__41744));
    InMux I__9343 (
            .O(N__41859),
            .I(N__41744));
    InMux I__9342 (
            .O(N__41858),
            .I(N__41733));
    InMux I__9341 (
            .O(N__41857),
            .I(N__41733));
    InMux I__9340 (
            .O(N__41856),
            .I(N__41733));
    InMux I__9339 (
            .O(N__41855),
            .I(N__41733));
    InMux I__9338 (
            .O(N__41854),
            .I(N__41728));
    InMux I__9337 (
            .O(N__41853),
            .I(N__41728));
    InMux I__9336 (
            .O(N__41852),
            .I(N__41723));
    InMux I__9335 (
            .O(N__41851),
            .I(N__41723));
    InMux I__9334 (
            .O(N__41850),
            .I(N__41718));
    InMux I__9333 (
            .O(N__41849),
            .I(N__41718));
    LocalMux I__9332 (
            .O(N__41844),
            .I(N__41711));
    LocalMux I__9331 (
            .O(N__41841),
            .I(N__41711));
    LocalMux I__9330 (
            .O(N__41834),
            .I(N__41711));
    InMux I__9329 (
            .O(N__41833),
            .I(N__41706));
    InMux I__9328 (
            .O(N__41832),
            .I(N__41706));
    LocalMux I__9327 (
            .O(N__41829),
            .I(N__41701));
    LocalMux I__9326 (
            .O(N__41826),
            .I(N__41701));
    InMux I__9325 (
            .O(N__41825),
            .I(N__41698));
    LocalMux I__9324 (
            .O(N__41822),
            .I(N__41695));
    InMux I__9323 (
            .O(N__41821),
            .I(N__41690));
    InMux I__9322 (
            .O(N__41820),
            .I(N__41690));
    LocalMux I__9321 (
            .O(N__41817),
            .I(N__41687));
    InMux I__9320 (
            .O(N__41816),
            .I(N__41684));
    InMux I__9319 (
            .O(N__41815),
            .I(N__41679));
    InMux I__9318 (
            .O(N__41814),
            .I(N__41679));
    LocalMux I__9317 (
            .O(N__41811),
            .I(N__41676));
    LocalMux I__9316 (
            .O(N__41806),
            .I(N__41669));
    LocalMux I__9315 (
            .O(N__41803),
            .I(N__41669));
    LocalMux I__9314 (
            .O(N__41796),
            .I(N__41669));
    InMux I__9313 (
            .O(N__41795),
            .I(N__41648));
    InMux I__9312 (
            .O(N__41794),
            .I(N__41635));
    InMux I__9311 (
            .O(N__41793),
            .I(N__41635));
    InMux I__9310 (
            .O(N__41792),
            .I(N__41635));
    InMux I__9309 (
            .O(N__41791),
            .I(N__41635));
    InMux I__9308 (
            .O(N__41790),
            .I(N__41635));
    InMux I__9307 (
            .O(N__41789),
            .I(N__41635));
    InMux I__9306 (
            .O(N__41788),
            .I(N__41628));
    InMux I__9305 (
            .O(N__41787),
            .I(N__41628));
    InMux I__9304 (
            .O(N__41786),
            .I(N__41628));
    InMux I__9303 (
            .O(N__41785),
            .I(N__41623));
    InMux I__9302 (
            .O(N__41784),
            .I(N__41623));
    InMux I__9301 (
            .O(N__41783),
            .I(N__41620));
    InMux I__9300 (
            .O(N__41782),
            .I(N__41613));
    InMux I__9299 (
            .O(N__41781),
            .I(N__41613));
    InMux I__9298 (
            .O(N__41780),
            .I(N__41613));
    InMux I__9297 (
            .O(N__41779),
            .I(N__41610));
    LocalMux I__9296 (
            .O(N__41776),
            .I(N__41607));
    InMux I__9295 (
            .O(N__41775),
            .I(N__41596));
    InMux I__9294 (
            .O(N__41774),
            .I(N__41596));
    InMux I__9293 (
            .O(N__41773),
            .I(N__41596));
    InMux I__9292 (
            .O(N__41772),
            .I(N__41596));
    InMux I__9291 (
            .O(N__41771),
            .I(N__41596));
    InMux I__9290 (
            .O(N__41770),
            .I(N__41589));
    InMux I__9289 (
            .O(N__41769),
            .I(N__41589));
    InMux I__9288 (
            .O(N__41768),
            .I(N__41589));
    LocalMux I__9287 (
            .O(N__41765),
            .I(N__41584));
    LocalMux I__9286 (
            .O(N__41762),
            .I(N__41584));
    Span4Mux_v I__9285 (
            .O(N__41757),
            .I(N__41577));
    Span4Mux_v I__9284 (
            .O(N__41752),
            .I(N__41577));
    LocalMux I__9283 (
            .O(N__41749),
            .I(N__41577));
    LocalMux I__9282 (
            .O(N__41744),
            .I(N__41574));
    InMux I__9281 (
            .O(N__41743),
            .I(N__41569));
    InMux I__9280 (
            .O(N__41742),
            .I(N__41569));
    LocalMux I__9279 (
            .O(N__41733),
            .I(N__41562));
    LocalMux I__9278 (
            .O(N__41728),
            .I(N__41562));
    LocalMux I__9277 (
            .O(N__41723),
            .I(N__41562));
    LocalMux I__9276 (
            .O(N__41718),
            .I(N__41551));
    Span4Mux_h I__9275 (
            .O(N__41711),
            .I(N__41551));
    LocalMux I__9274 (
            .O(N__41706),
            .I(N__41551));
    Span4Mux_s3_v I__9273 (
            .O(N__41701),
            .I(N__41551));
    LocalMux I__9272 (
            .O(N__41698),
            .I(N__41551));
    Span4Mux_h I__9271 (
            .O(N__41695),
            .I(N__41548));
    LocalMux I__9270 (
            .O(N__41690),
            .I(N__41543));
    Span4Mux_v I__9269 (
            .O(N__41687),
            .I(N__41543));
    LocalMux I__9268 (
            .O(N__41684),
            .I(N__41534));
    LocalMux I__9267 (
            .O(N__41679),
            .I(N__41534));
    Span4Mux_v I__9266 (
            .O(N__41676),
            .I(N__41534));
    Span4Mux_v I__9265 (
            .O(N__41669),
            .I(N__41534));
    InMux I__9264 (
            .O(N__41668),
            .I(N__41531));
    InMux I__9263 (
            .O(N__41667),
            .I(N__41524));
    InMux I__9262 (
            .O(N__41666),
            .I(N__41524));
    InMux I__9261 (
            .O(N__41665),
            .I(N__41524));
    InMux I__9260 (
            .O(N__41664),
            .I(N__41513));
    InMux I__9259 (
            .O(N__41663),
            .I(N__41513));
    InMux I__9258 (
            .O(N__41662),
            .I(N__41513));
    InMux I__9257 (
            .O(N__41661),
            .I(N__41513));
    InMux I__9256 (
            .O(N__41660),
            .I(N__41513));
    InMux I__9255 (
            .O(N__41659),
            .I(N__41500));
    InMux I__9254 (
            .O(N__41658),
            .I(N__41500));
    InMux I__9253 (
            .O(N__41657),
            .I(N__41500));
    InMux I__9252 (
            .O(N__41656),
            .I(N__41500));
    InMux I__9251 (
            .O(N__41655),
            .I(N__41500));
    InMux I__9250 (
            .O(N__41654),
            .I(N__41500));
    InMux I__9249 (
            .O(N__41653),
            .I(N__41497));
    InMux I__9248 (
            .O(N__41652),
            .I(N__41492));
    InMux I__9247 (
            .O(N__41651),
            .I(N__41492));
    LocalMux I__9246 (
            .O(N__41648),
            .I(N__41485));
    LocalMux I__9245 (
            .O(N__41635),
            .I(N__41485));
    LocalMux I__9244 (
            .O(N__41628),
            .I(N__41485));
    LocalMux I__9243 (
            .O(N__41623),
            .I(N__41482));
    LocalMux I__9242 (
            .O(N__41620),
            .I(N__41477));
    LocalMux I__9241 (
            .O(N__41613),
            .I(N__41477));
    LocalMux I__9240 (
            .O(N__41610),
            .I(N__41474));
    Span12Mux_s7_v I__9239 (
            .O(N__41607),
            .I(N__41471));
    LocalMux I__9238 (
            .O(N__41596),
            .I(N__41462));
    LocalMux I__9237 (
            .O(N__41589),
            .I(N__41462));
    Span4Mux_h I__9236 (
            .O(N__41584),
            .I(N__41462));
    Span4Mux_h I__9235 (
            .O(N__41577),
            .I(N__41462));
    Span4Mux_v I__9234 (
            .O(N__41574),
            .I(N__41447));
    LocalMux I__9233 (
            .O(N__41569),
            .I(N__41447));
    Span4Mux_v I__9232 (
            .O(N__41562),
            .I(N__41447));
    Span4Mux_v I__9231 (
            .O(N__41551),
            .I(N__41447));
    Span4Mux_v I__9230 (
            .O(N__41548),
            .I(N__41447));
    Span4Mux_h I__9229 (
            .O(N__41543),
            .I(N__41447));
    Span4Mux_h I__9228 (
            .O(N__41534),
            .I(N__41447));
    LocalMux I__9227 (
            .O(N__41531),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__9226 (
            .O(N__41524),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__9225 (
            .O(N__41513),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__9224 (
            .O(N__41500),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__9223 (
            .O(N__41497),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__9222 (
            .O(N__41492),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__9221 (
            .O(N__41485),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__9220 (
            .O(N__41482),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__9219 (
            .O(N__41477),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv12 I__9218 (
            .O(N__41474),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv12 I__9217 (
            .O(N__41471),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__9216 (
            .O(N__41462),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__9215 (
            .O(N__41447),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    InMux I__9214 (
            .O(N__41420),
            .I(N__41416));
    InMux I__9213 (
            .O(N__41419),
            .I(N__41412));
    LocalMux I__9212 (
            .O(N__41416),
            .I(N__41409));
    InMux I__9211 (
            .O(N__41415),
            .I(N__41406));
    LocalMux I__9210 (
            .O(N__41412),
            .I(N__41403));
    Span12Mux_h I__9209 (
            .O(N__41409),
            .I(N__41400));
    LocalMux I__9208 (
            .O(N__41406),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    Odrv12 I__9207 (
            .O(N__41403),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    Odrv12 I__9206 (
            .O(N__41400),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    InMux I__9205 (
            .O(N__41393),
            .I(N__41390));
    LocalMux I__9204 (
            .O(N__41390),
            .I(N__41387));
    Span4Mux_h I__9203 (
            .O(N__41387),
            .I(N__41383));
    InMux I__9202 (
            .O(N__41386),
            .I(N__41380));
    Odrv4 I__9201 (
            .O(N__41383),
            .I(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ));
    LocalMux I__9200 (
            .O(N__41380),
            .I(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ));
    InMux I__9199 (
            .O(N__41375),
            .I(N__41372));
    LocalMux I__9198 (
            .O(N__41372),
            .I(N__41368));
    InMux I__9197 (
            .O(N__41371),
            .I(N__41364));
    Span4Mux_h I__9196 (
            .O(N__41368),
            .I(N__41361));
    InMux I__9195 (
            .O(N__41367),
            .I(N__41358));
    LocalMux I__9194 (
            .O(N__41364),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    Odrv4 I__9193 (
            .O(N__41361),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    LocalMux I__9192 (
            .O(N__41358),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    InMux I__9191 (
            .O(N__41351),
            .I(N__41345));
    InMux I__9190 (
            .O(N__41350),
            .I(N__41345));
    LocalMux I__9189 (
            .O(N__41345),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ));
    CascadeMux I__9188 (
            .O(N__41342),
            .I(N__41339));
    InMux I__9187 (
            .O(N__41339),
            .I(N__41333));
    InMux I__9186 (
            .O(N__41338),
            .I(N__41333));
    LocalMux I__9185 (
            .O(N__41333),
            .I(N__41330));
    Odrv4 I__9184 (
            .O(N__41330),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ));
    CascadeMux I__9183 (
            .O(N__41327),
            .I(N__41324));
    InMux I__9182 (
            .O(N__41324),
            .I(N__41321));
    LocalMux I__9181 (
            .O(N__41321),
            .I(N__41318));
    Odrv4 I__9180 (
            .O(N__41318),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__9179 (
            .O(N__41315),
            .I(N__41311));
    CascadeMux I__9178 (
            .O(N__41314),
            .I(N__41308));
    InMux I__9177 (
            .O(N__41311),
            .I(N__41305));
    InMux I__9176 (
            .O(N__41308),
            .I(N__41301));
    LocalMux I__9175 (
            .O(N__41305),
            .I(N__41298));
    InMux I__9174 (
            .O(N__41304),
            .I(N__41294));
    LocalMux I__9173 (
            .O(N__41301),
            .I(N__41291));
    Span12Mux_v I__9172 (
            .O(N__41298),
            .I(N__41288));
    InMux I__9171 (
            .O(N__41297),
            .I(N__41285));
    LocalMux I__9170 (
            .O(N__41294),
            .I(N__41280));
    Span4Mux_v I__9169 (
            .O(N__41291),
            .I(N__41280));
    Odrv12 I__9168 (
            .O(N__41288),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    LocalMux I__9167 (
            .O(N__41285),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__9166 (
            .O(N__41280),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    InMux I__9165 (
            .O(N__41273),
            .I(bfn_15_26_0_));
    CascadeMux I__9164 (
            .O(N__41270),
            .I(N__41266));
    InMux I__9163 (
            .O(N__41269),
            .I(N__41263));
    InMux I__9162 (
            .O(N__41266),
            .I(N__41260));
    LocalMux I__9161 (
            .O(N__41263),
            .I(N__41255));
    LocalMux I__9160 (
            .O(N__41260),
            .I(N__41252));
    InMux I__9159 (
            .O(N__41259),
            .I(N__41249));
    InMux I__9158 (
            .O(N__41258),
            .I(N__41246));
    Span12Mux_h I__9157 (
            .O(N__41255),
            .I(N__41239));
    Sp12to4 I__9156 (
            .O(N__41252),
            .I(N__41239));
    LocalMux I__9155 (
            .O(N__41249),
            .I(N__41239));
    LocalMux I__9154 (
            .O(N__41246),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv12 I__9153 (
            .O(N__41239),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    InMux I__9152 (
            .O(N__41234),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    CascadeMux I__9151 (
            .O(N__41231),
            .I(N__41228));
    InMux I__9150 (
            .O(N__41228),
            .I(N__41225));
    LocalMux I__9149 (
            .O(N__41225),
            .I(N__41221));
    InMux I__9148 (
            .O(N__41224),
            .I(N__41218));
    Span4Mux_v I__9147 (
            .O(N__41221),
            .I(N__41215));
    LocalMux I__9146 (
            .O(N__41218),
            .I(N__41212));
    Sp12to4 I__9145 (
            .O(N__41215),
            .I(N__41208));
    Span4Mux_h I__9144 (
            .O(N__41212),
            .I(N__41204));
    InMux I__9143 (
            .O(N__41211),
            .I(N__41201));
    Span12Mux_h I__9142 (
            .O(N__41208),
            .I(N__41198));
    InMux I__9141 (
            .O(N__41207),
            .I(N__41195));
    Span4Mux_v I__9140 (
            .O(N__41204),
            .I(N__41192));
    LocalMux I__9139 (
            .O(N__41201),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv12 I__9138 (
            .O(N__41198),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    LocalMux I__9137 (
            .O(N__41195),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__9136 (
            .O(N__41192),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    InMux I__9135 (
            .O(N__41183),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    InMux I__9134 (
            .O(N__41180),
            .I(N__41176));
    InMux I__9133 (
            .O(N__41179),
            .I(N__41173));
    LocalMux I__9132 (
            .O(N__41176),
            .I(N__41170));
    LocalMux I__9131 (
            .O(N__41173),
            .I(N__41165));
    Span12Mux_v I__9130 (
            .O(N__41170),
            .I(N__41162));
    InMux I__9129 (
            .O(N__41169),
            .I(N__41159));
    InMux I__9128 (
            .O(N__41168),
            .I(N__41156));
    Span4Mux_v I__9127 (
            .O(N__41165),
            .I(N__41153));
    Odrv12 I__9126 (
            .O(N__41162),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__9125 (
            .O(N__41159),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__9124 (
            .O(N__41156),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__9123 (
            .O(N__41153),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    InMux I__9122 (
            .O(N__41144),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ));
    CascadeMux I__9121 (
            .O(N__41141),
            .I(N__41137));
    InMux I__9120 (
            .O(N__41140),
            .I(N__41133));
    InMux I__9119 (
            .O(N__41137),
            .I(N__41130));
    InMux I__9118 (
            .O(N__41136),
            .I(N__41127));
    LocalMux I__9117 (
            .O(N__41133),
            .I(N__41124));
    LocalMux I__9116 (
            .O(N__41130),
            .I(N__41121));
    LocalMux I__9115 (
            .O(N__41127),
            .I(N__41115));
    Span4Mux_v I__9114 (
            .O(N__41124),
            .I(N__41115));
    Span12Mux_v I__9113 (
            .O(N__41121),
            .I(N__41112));
    InMux I__9112 (
            .O(N__41120),
            .I(N__41109));
    Span4Mux_v I__9111 (
            .O(N__41115),
            .I(N__41106));
    Odrv12 I__9110 (
            .O(N__41112),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    LocalMux I__9109 (
            .O(N__41109),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv4 I__9108 (
            .O(N__41106),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    InMux I__9107 (
            .O(N__41099),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    InMux I__9106 (
            .O(N__41096),
            .I(N__41093));
    LocalMux I__9105 (
            .O(N__41093),
            .I(N__41089));
    InMux I__9104 (
            .O(N__41092),
            .I(N__41085));
    Span12Mux_s10_h I__9103 (
            .O(N__41089),
            .I(N__41082));
    CascadeMux I__9102 (
            .O(N__41088),
            .I(N__41079));
    LocalMux I__9101 (
            .O(N__41085),
            .I(N__41075));
    Span12Mux_h I__9100 (
            .O(N__41082),
            .I(N__41072));
    InMux I__9099 (
            .O(N__41079),
            .I(N__41069));
    InMux I__9098 (
            .O(N__41078),
            .I(N__41066));
    Span4Mux_v I__9097 (
            .O(N__41075),
            .I(N__41063));
    Odrv12 I__9096 (
            .O(N__41072),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    LocalMux I__9095 (
            .O(N__41069),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    LocalMux I__9094 (
            .O(N__41066),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__9093 (
            .O(N__41063),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    InMux I__9092 (
            .O(N__41054),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    InMux I__9091 (
            .O(N__41051),
            .I(N__41047));
    CascadeMux I__9090 (
            .O(N__41050),
            .I(N__41043));
    LocalMux I__9089 (
            .O(N__41047),
            .I(N__41037));
    InMux I__9088 (
            .O(N__41046),
            .I(N__41028));
    InMux I__9087 (
            .O(N__41043),
            .I(N__41025));
    InMux I__9086 (
            .O(N__41042),
            .I(N__41022));
    InMux I__9085 (
            .O(N__41041),
            .I(N__41017));
    InMux I__9084 (
            .O(N__41040),
            .I(N__41017));
    Sp12to4 I__9083 (
            .O(N__41037),
            .I(N__41014));
    InMux I__9082 (
            .O(N__41036),
            .I(N__40992));
    InMux I__9081 (
            .O(N__41035),
            .I(N__40989));
    InMux I__9080 (
            .O(N__41034),
            .I(N__40980));
    InMux I__9079 (
            .O(N__41033),
            .I(N__40980));
    InMux I__9078 (
            .O(N__41032),
            .I(N__40980));
    InMux I__9077 (
            .O(N__41031),
            .I(N__40980));
    LocalMux I__9076 (
            .O(N__41028),
            .I(N__40977));
    LocalMux I__9075 (
            .O(N__41025),
            .I(N__40972));
    LocalMux I__9074 (
            .O(N__41022),
            .I(N__40972));
    LocalMux I__9073 (
            .O(N__41017),
            .I(N__40968));
    Span12Mux_v I__9072 (
            .O(N__41014),
            .I(N__40965));
    InMux I__9071 (
            .O(N__41013),
            .I(N__40962));
    InMux I__9070 (
            .O(N__41012),
            .I(N__40959));
    InMux I__9069 (
            .O(N__41011),
            .I(N__40956));
    InMux I__9068 (
            .O(N__41010),
            .I(N__40949));
    InMux I__9067 (
            .O(N__41009),
            .I(N__40949));
    InMux I__9066 (
            .O(N__41008),
            .I(N__40949));
    InMux I__9065 (
            .O(N__41007),
            .I(N__40946));
    InMux I__9064 (
            .O(N__41006),
            .I(N__40931));
    InMux I__9063 (
            .O(N__41005),
            .I(N__40931));
    InMux I__9062 (
            .O(N__41004),
            .I(N__40931));
    InMux I__9061 (
            .O(N__41003),
            .I(N__40931));
    InMux I__9060 (
            .O(N__41002),
            .I(N__40931));
    InMux I__9059 (
            .O(N__41001),
            .I(N__40931));
    InMux I__9058 (
            .O(N__41000),
            .I(N__40931));
    InMux I__9057 (
            .O(N__40999),
            .I(N__40920));
    InMux I__9056 (
            .O(N__40998),
            .I(N__40920));
    InMux I__9055 (
            .O(N__40997),
            .I(N__40920));
    InMux I__9054 (
            .O(N__40996),
            .I(N__40920));
    InMux I__9053 (
            .O(N__40995),
            .I(N__40920));
    LocalMux I__9052 (
            .O(N__40992),
            .I(N__40917));
    LocalMux I__9051 (
            .O(N__40989),
            .I(N__40908));
    LocalMux I__9050 (
            .O(N__40980),
            .I(N__40908));
    Span4Mux_h I__9049 (
            .O(N__40977),
            .I(N__40908));
    Span4Mux_h I__9048 (
            .O(N__40972),
            .I(N__40908));
    InMux I__9047 (
            .O(N__40971),
            .I(N__40905));
    Span12Mux_s4_h I__9046 (
            .O(N__40968),
            .I(N__40898));
    Span12Mux_h I__9045 (
            .O(N__40965),
            .I(N__40898));
    LocalMux I__9044 (
            .O(N__40962),
            .I(N__40898));
    LocalMux I__9043 (
            .O(N__40959),
            .I(N__40895));
    LocalMux I__9042 (
            .O(N__40956),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__9041 (
            .O(N__40949),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__9040 (
            .O(N__40946),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__9039 (
            .O(N__40931),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__9038 (
            .O(N__40920),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__9037 (
            .O(N__40917),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__9036 (
            .O(N__40908),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__9035 (
            .O(N__40905),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv12 I__9034 (
            .O(N__40898),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__9033 (
            .O(N__40895),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    CascadeMux I__9032 (
            .O(N__40874),
            .I(N__40863));
    CascadeMux I__9031 (
            .O(N__40873),
            .I(N__40859));
    CascadeMux I__9030 (
            .O(N__40872),
            .I(N__40855));
    CascadeMux I__9029 (
            .O(N__40871),
            .I(N__40851));
    CascadeMux I__9028 (
            .O(N__40870),
            .I(N__40847));
    CascadeMux I__9027 (
            .O(N__40869),
            .I(N__40843));
    CascadeMux I__9026 (
            .O(N__40868),
            .I(N__40839));
    CascadeMux I__9025 (
            .O(N__40867),
            .I(N__40834));
    InMux I__9024 (
            .O(N__40866),
            .I(N__40818));
    InMux I__9023 (
            .O(N__40863),
            .I(N__40818));
    InMux I__9022 (
            .O(N__40862),
            .I(N__40818));
    InMux I__9021 (
            .O(N__40859),
            .I(N__40818));
    InMux I__9020 (
            .O(N__40858),
            .I(N__40818));
    InMux I__9019 (
            .O(N__40855),
            .I(N__40818));
    InMux I__9018 (
            .O(N__40854),
            .I(N__40818));
    InMux I__9017 (
            .O(N__40851),
            .I(N__40801));
    InMux I__9016 (
            .O(N__40850),
            .I(N__40801));
    InMux I__9015 (
            .O(N__40847),
            .I(N__40801));
    InMux I__9014 (
            .O(N__40846),
            .I(N__40801));
    InMux I__9013 (
            .O(N__40843),
            .I(N__40801));
    InMux I__9012 (
            .O(N__40842),
            .I(N__40801));
    InMux I__9011 (
            .O(N__40839),
            .I(N__40801));
    InMux I__9010 (
            .O(N__40838),
            .I(N__40801));
    InMux I__9009 (
            .O(N__40837),
            .I(N__40794));
    InMux I__9008 (
            .O(N__40834),
            .I(N__40794));
    InMux I__9007 (
            .O(N__40833),
            .I(N__40794));
    LocalMux I__9006 (
            .O(N__40818),
            .I(N__40787));
    LocalMux I__9005 (
            .O(N__40801),
            .I(N__40787));
    LocalMux I__9004 (
            .O(N__40794),
            .I(N__40787));
    Span4Mux_v I__9003 (
            .O(N__40787),
            .I(N__40784));
    Odrv4 I__9002 (
            .O(N__40784),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    InMux I__9001 (
            .O(N__40781),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    InMux I__9000 (
            .O(N__40778),
            .I(N__40775));
    LocalMux I__8999 (
            .O(N__40775),
            .I(N__40771));
    InMux I__8998 (
            .O(N__40774),
            .I(N__40768));
    Odrv4 I__8997 (
            .O(N__40771),
            .I(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ));
    LocalMux I__8996 (
            .O(N__40768),
            .I(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ));
    CascadeMux I__8995 (
            .O(N__40763),
            .I(N__40760));
    InMux I__8994 (
            .O(N__40760),
            .I(N__40756));
    InMux I__8993 (
            .O(N__40759),
            .I(N__40753));
    LocalMux I__8992 (
            .O(N__40756),
            .I(N__40750));
    LocalMux I__8991 (
            .O(N__40753),
            .I(N__40744));
    Span4Mux_v I__8990 (
            .O(N__40750),
            .I(N__40744));
    InMux I__8989 (
            .O(N__40749),
            .I(N__40741));
    Odrv4 I__8988 (
            .O(N__40744),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    LocalMux I__8987 (
            .O(N__40741),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    CascadeMux I__8986 (
            .O(N__40736),
            .I(N__40732));
    CascadeMux I__8985 (
            .O(N__40735),
            .I(N__40729));
    InMux I__8984 (
            .O(N__40732),
            .I(N__40726));
    InMux I__8983 (
            .O(N__40729),
            .I(N__40722));
    LocalMux I__8982 (
            .O(N__40726),
            .I(N__40719));
    CascadeMux I__8981 (
            .O(N__40725),
            .I(N__40716));
    LocalMux I__8980 (
            .O(N__40722),
            .I(N__40713));
    Span4Mux_h I__8979 (
            .O(N__40719),
            .I(N__40710));
    InMux I__8978 (
            .O(N__40716),
            .I(N__40706));
    Span4Mux_v I__8977 (
            .O(N__40713),
            .I(N__40703));
    Sp12to4 I__8976 (
            .O(N__40710),
            .I(N__40700));
    InMux I__8975 (
            .O(N__40709),
            .I(N__40697));
    LocalMux I__8974 (
            .O(N__40706),
            .I(N__40694));
    Span4Mux_v I__8973 (
            .O(N__40703),
            .I(N__40691));
    Span12Mux_v I__8972 (
            .O(N__40700),
            .I(N__40688));
    LocalMux I__8971 (
            .O(N__40697),
            .I(N__40683));
    Span4Mux_v I__8970 (
            .O(N__40694),
            .I(N__40683));
    Odrv4 I__8969 (
            .O(N__40691),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv12 I__8968 (
            .O(N__40688),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__8967 (
            .O(N__40683),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    InMux I__8966 (
            .O(N__40676),
            .I(bfn_15_25_0_));
    InMux I__8965 (
            .O(N__40673),
            .I(N__40670));
    LocalMux I__8964 (
            .O(N__40670),
            .I(N__40666));
    InMux I__8963 (
            .O(N__40669),
            .I(N__40662));
    Span12Mux_s7_v I__8962 (
            .O(N__40666),
            .I(N__40658));
    InMux I__8961 (
            .O(N__40665),
            .I(N__40655));
    LocalMux I__8960 (
            .O(N__40662),
            .I(N__40652));
    InMux I__8959 (
            .O(N__40661),
            .I(N__40649));
    Span12Mux_h I__8958 (
            .O(N__40658),
            .I(N__40646));
    LocalMux I__8957 (
            .O(N__40655),
            .I(N__40643));
    Span4Mux_v I__8956 (
            .O(N__40652),
            .I(N__40640));
    LocalMux I__8955 (
            .O(N__40649),
            .I(N__40637));
    Odrv12 I__8954 (
            .O(N__40646),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__8953 (
            .O(N__40643),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__8952 (
            .O(N__40640),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__8951 (
            .O(N__40637),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    InMux I__8950 (
            .O(N__40628),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    CascadeMux I__8949 (
            .O(N__40625),
            .I(N__40622));
    InMux I__8948 (
            .O(N__40622),
            .I(N__40619));
    LocalMux I__8947 (
            .O(N__40619),
            .I(N__40616));
    Span4Mux_v I__8946 (
            .O(N__40616),
            .I(N__40611));
    InMux I__8945 (
            .O(N__40615),
            .I(N__40608));
    InMux I__8944 (
            .O(N__40614),
            .I(N__40605));
    Sp12to4 I__8943 (
            .O(N__40611),
            .I(N__40599));
    LocalMux I__8942 (
            .O(N__40608),
            .I(N__40599));
    LocalMux I__8941 (
            .O(N__40605),
            .I(N__40596));
    InMux I__8940 (
            .O(N__40604),
            .I(N__40593));
    Span12Mux_h I__8939 (
            .O(N__40599),
            .I(N__40590));
    Span4Mux_v I__8938 (
            .O(N__40596),
            .I(N__40587));
    LocalMux I__8937 (
            .O(N__40593),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv12 I__8936 (
            .O(N__40590),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__8935 (
            .O(N__40587),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    InMux I__8934 (
            .O(N__40580),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    InMux I__8933 (
            .O(N__40577),
            .I(N__40574));
    LocalMux I__8932 (
            .O(N__40574),
            .I(N__40570));
    InMux I__8931 (
            .O(N__40573),
            .I(N__40567));
    Span4Mux_v I__8930 (
            .O(N__40570),
            .I(N__40564));
    LocalMux I__8929 (
            .O(N__40567),
            .I(N__40561));
    Sp12to4 I__8928 (
            .O(N__40564),
            .I(N__40557));
    Span4Mux_h I__8927 (
            .O(N__40561),
            .I(N__40554));
    InMux I__8926 (
            .O(N__40560),
            .I(N__40551));
    Span12Mux_h I__8925 (
            .O(N__40557),
            .I(N__40543));
    Sp12to4 I__8924 (
            .O(N__40554),
            .I(N__40543));
    LocalMux I__8923 (
            .O(N__40551),
            .I(N__40543));
    InMux I__8922 (
            .O(N__40550),
            .I(N__40540));
    Span12Mux_v I__8921 (
            .O(N__40543),
            .I(N__40537));
    LocalMux I__8920 (
            .O(N__40540),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv12 I__8919 (
            .O(N__40537),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    InMux I__8918 (
            .O(N__40532),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ));
    CascadeMux I__8917 (
            .O(N__40529),
            .I(N__40525));
    CascadeMux I__8916 (
            .O(N__40528),
            .I(N__40522));
    InMux I__8915 (
            .O(N__40525),
            .I(N__40519));
    InMux I__8914 (
            .O(N__40522),
            .I(N__40516));
    LocalMux I__8913 (
            .O(N__40519),
            .I(N__40511));
    LocalMux I__8912 (
            .O(N__40516),
            .I(N__40508));
    InMux I__8911 (
            .O(N__40515),
            .I(N__40505));
    InMux I__8910 (
            .O(N__40514),
            .I(N__40502));
    Span4Mux_v I__8909 (
            .O(N__40511),
            .I(N__40499));
    Span12Mux_h I__8908 (
            .O(N__40508),
            .I(N__40494));
    LocalMux I__8907 (
            .O(N__40505),
            .I(N__40494));
    LocalMux I__8906 (
            .O(N__40502),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv4 I__8905 (
            .O(N__40499),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv12 I__8904 (
            .O(N__40494),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    InMux I__8903 (
            .O(N__40487),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    InMux I__8902 (
            .O(N__40484),
            .I(N__40481));
    LocalMux I__8901 (
            .O(N__40481),
            .I(N__40478));
    Sp12to4 I__8900 (
            .O(N__40478),
            .I(N__40474));
    InMux I__8899 (
            .O(N__40477),
            .I(N__40470));
    Span12Mux_v I__8898 (
            .O(N__40474),
            .I(N__40466));
    InMux I__8897 (
            .O(N__40473),
            .I(N__40463));
    LocalMux I__8896 (
            .O(N__40470),
            .I(N__40460));
    InMux I__8895 (
            .O(N__40469),
            .I(N__40457));
    Span12Mux_h I__8894 (
            .O(N__40466),
            .I(N__40454));
    LocalMux I__8893 (
            .O(N__40463),
            .I(N__40451));
    Span4Mux_v I__8892 (
            .O(N__40460),
            .I(N__40448));
    LocalMux I__8891 (
            .O(N__40457),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv12 I__8890 (
            .O(N__40454),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv12 I__8889 (
            .O(N__40451),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__8888 (
            .O(N__40448),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    InMux I__8887 (
            .O(N__40439),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    CascadeMux I__8886 (
            .O(N__40436),
            .I(N__40433));
    InMux I__8885 (
            .O(N__40433),
            .I(N__40430));
    LocalMux I__8884 (
            .O(N__40430),
            .I(N__40427));
    Span4Mux_v I__8883 (
            .O(N__40427),
            .I(N__40424));
    Span4Mux_h I__8882 (
            .O(N__40424),
            .I(N__40421));
    Span4Mux_h I__8881 (
            .O(N__40421),
            .I(N__40417));
    InMux I__8880 (
            .O(N__40420),
            .I(N__40414));
    Span4Mux_h I__8879 (
            .O(N__40417),
            .I(N__40407));
    LocalMux I__8878 (
            .O(N__40414),
            .I(N__40407));
    InMux I__8877 (
            .O(N__40413),
            .I(N__40404));
    InMux I__8876 (
            .O(N__40412),
            .I(N__40401));
    Span4Mux_v I__8875 (
            .O(N__40407),
            .I(N__40396));
    LocalMux I__8874 (
            .O(N__40404),
            .I(N__40396));
    LocalMux I__8873 (
            .O(N__40401),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__8872 (
            .O(N__40396),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    InMux I__8871 (
            .O(N__40391),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    InMux I__8870 (
            .O(N__40388),
            .I(N__40385));
    LocalMux I__8869 (
            .O(N__40385),
            .I(N__40380));
    InMux I__8868 (
            .O(N__40384),
            .I(N__40376));
    InMux I__8867 (
            .O(N__40383),
            .I(N__40373));
    Sp12to4 I__8866 (
            .O(N__40380),
            .I(N__40370));
    CascadeMux I__8865 (
            .O(N__40379),
            .I(N__40367));
    LocalMux I__8864 (
            .O(N__40376),
            .I(N__40362));
    LocalMux I__8863 (
            .O(N__40373),
            .I(N__40362));
    Span12Mux_v I__8862 (
            .O(N__40370),
            .I(N__40359));
    InMux I__8861 (
            .O(N__40367),
            .I(N__40356));
    Span4Mux_v I__8860 (
            .O(N__40362),
            .I(N__40353));
    Odrv12 I__8859 (
            .O(N__40359),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    LocalMux I__8858 (
            .O(N__40356),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__8857 (
            .O(N__40353),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    InMux I__8856 (
            .O(N__40346),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ));
    InMux I__8855 (
            .O(N__40343),
            .I(N__40340));
    LocalMux I__8854 (
            .O(N__40340),
            .I(N__40337));
    Odrv4 I__8853 (
            .O(N__40337),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    CascadeMux I__8852 (
            .O(N__40334),
            .I(N__40331));
    InMux I__8851 (
            .O(N__40331),
            .I(N__40328));
    LocalMux I__8850 (
            .O(N__40328),
            .I(N__40324));
    InMux I__8849 (
            .O(N__40327),
            .I(N__40320));
    Span4Mux_v I__8848 (
            .O(N__40324),
            .I(N__40317));
    InMux I__8847 (
            .O(N__40323),
            .I(N__40314));
    LocalMux I__8846 (
            .O(N__40320),
            .I(N__40311));
    Span4Mux_h I__8845 (
            .O(N__40317),
            .I(N__40308));
    LocalMux I__8844 (
            .O(N__40314),
            .I(N__40303));
    Span4Mux_v I__8843 (
            .O(N__40311),
            .I(N__40303));
    Sp12to4 I__8842 (
            .O(N__40308),
            .I(N__40299));
    Span4Mux_v I__8841 (
            .O(N__40303),
            .I(N__40296));
    InMux I__8840 (
            .O(N__40302),
            .I(N__40293));
    Span12Mux_h I__8839 (
            .O(N__40299),
            .I(N__40290));
    Odrv4 I__8838 (
            .O(N__40296),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    LocalMux I__8837 (
            .O(N__40293),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv12 I__8836 (
            .O(N__40290),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    InMux I__8835 (
            .O(N__40283),
            .I(bfn_15_24_0_));
    InMux I__8834 (
            .O(N__40280),
            .I(N__40277));
    LocalMux I__8833 (
            .O(N__40277),
            .I(N__40274));
    Odrv12 I__8832 (
            .O(N__40274),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    CascadeMux I__8831 (
            .O(N__40271),
            .I(N__40268));
    InMux I__8830 (
            .O(N__40268),
            .I(N__40265));
    LocalMux I__8829 (
            .O(N__40265),
            .I(N__40262));
    Span4Mux_v I__8828 (
            .O(N__40262),
            .I(N__40258));
    CascadeMux I__8827 (
            .O(N__40261),
            .I(N__40255));
    Span4Mux_v I__8826 (
            .O(N__40258),
            .I(N__40251));
    InMux I__8825 (
            .O(N__40255),
            .I(N__40247));
    InMux I__8824 (
            .O(N__40254),
            .I(N__40244));
    Span4Mux_v I__8823 (
            .O(N__40251),
            .I(N__40241));
    InMux I__8822 (
            .O(N__40250),
            .I(N__40238));
    LocalMux I__8821 (
            .O(N__40247),
            .I(N__40235));
    LocalMux I__8820 (
            .O(N__40244),
            .I(N__40232));
    Sp12to4 I__8819 (
            .O(N__40241),
            .I(N__40229));
    LocalMux I__8818 (
            .O(N__40238),
            .I(N__40222));
    Span4Mux_v I__8817 (
            .O(N__40235),
            .I(N__40222));
    Span4Mux_h I__8816 (
            .O(N__40232),
            .I(N__40222));
    Odrv12 I__8815 (
            .O(N__40229),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv4 I__8814 (
            .O(N__40222),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    InMux I__8813 (
            .O(N__40217),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    InMux I__8812 (
            .O(N__40214),
            .I(N__40211));
    LocalMux I__8811 (
            .O(N__40211),
            .I(N__40208));
    Span12Mux_h I__8810 (
            .O(N__40208),
            .I(N__40205));
    Odrv12 I__8809 (
            .O(N__40205),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    CascadeMux I__8808 (
            .O(N__40202),
            .I(N__40199));
    InMux I__8807 (
            .O(N__40199),
            .I(N__40195));
    CascadeMux I__8806 (
            .O(N__40198),
            .I(N__40191));
    LocalMux I__8805 (
            .O(N__40195),
            .I(N__40188));
    InMux I__8804 (
            .O(N__40194),
            .I(N__40185));
    InMux I__8803 (
            .O(N__40191),
            .I(N__40182));
    Sp12to4 I__8802 (
            .O(N__40188),
            .I(N__40178));
    LocalMux I__8801 (
            .O(N__40185),
            .I(N__40175));
    LocalMux I__8800 (
            .O(N__40182),
            .I(N__40172));
    InMux I__8799 (
            .O(N__40181),
            .I(N__40169));
    Span12Mux_h I__8798 (
            .O(N__40178),
            .I(N__40166));
    Span4Mux_v I__8797 (
            .O(N__40175),
            .I(N__40161));
    Span4Mux_v I__8796 (
            .O(N__40172),
            .I(N__40161));
    LocalMux I__8795 (
            .O(N__40169),
            .I(N__40158));
    Odrv12 I__8794 (
            .O(N__40166),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__8793 (
            .O(N__40161),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__8792 (
            .O(N__40158),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    InMux I__8791 (
            .O(N__40151),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    InMux I__8790 (
            .O(N__40148),
            .I(N__40145));
    LocalMux I__8789 (
            .O(N__40145),
            .I(N__40142));
    Sp12to4 I__8788 (
            .O(N__40142),
            .I(N__40139));
    Odrv12 I__8787 (
            .O(N__40139),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    CascadeMux I__8786 (
            .O(N__40136),
            .I(N__40133));
    InMux I__8785 (
            .O(N__40133),
            .I(N__40130));
    LocalMux I__8784 (
            .O(N__40130),
            .I(N__40125));
    InMux I__8783 (
            .O(N__40129),
            .I(N__40122));
    InMux I__8782 (
            .O(N__40128),
            .I(N__40119));
    Span4Mux_v I__8781 (
            .O(N__40125),
            .I(N__40115));
    LocalMux I__8780 (
            .O(N__40122),
            .I(N__40112));
    LocalMux I__8779 (
            .O(N__40119),
            .I(N__40109));
    CascadeMux I__8778 (
            .O(N__40118),
            .I(N__40106));
    Sp12to4 I__8777 (
            .O(N__40115),
            .I(N__40103));
    Span4Mux_v I__8776 (
            .O(N__40112),
            .I(N__40098));
    Span4Mux_v I__8775 (
            .O(N__40109),
            .I(N__40098));
    InMux I__8774 (
            .O(N__40106),
            .I(N__40095));
    Span12Mux_h I__8773 (
            .O(N__40103),
            .I(N__40092));
    Odrv4 I__8772 (
            .O(N__40098),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    LocalMux I__8771 (
            .O(N__40095),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv12 I__8770 (
            .O(N__40092),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    InMux I__8769 (
            .O(N__40085),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ));
    InMux I__8768 (
            .O(N__40082),
            .I(N__40077));
    CascadeMux I__8767 (
            .O(N__40081),
            .I(N__40074));
    InMux I__8766 (
            .O(N__40080),
            .I(N__40071));
    LocalMux I__8765 (
            .O(N__40077),
            .I(N__40068));
    InMux I__8764 (
            .O(N__40074),
            .I(N__40064));
    LocalMux I__8763 (
            .O(N__40071),
            .I(N__40061));
    Span12Mux_v I__8762 (
            .O(N__40068),
            .I(N__40058));
    InMux I__8761 (
            .O(N__40067),
            .I(N__40055));
    LocalMux I__8760 (
            .O(N__40064),
            .I(N__40050));
    Span4Mux_v I__8759 (
            .O(N__40061),
            .I(N__40050));
    Odrv12 I__8758 (
            .O(N__40058),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    LocalMux I__8757 (
            .O(N__40055),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__8756 (
            .O(N__40050),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    CascadeMux I__8755 (
            .O(N__40043),
            .I(N__40040));
    InMux I__8754 (
            .O(N__40040),
            .I(N__40037));
    LocalMux I__8753 (
            .O(N__40037),
            .I(N__40034));
    Odrv12 I__8752 (
            .O(N__40034),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ));
    InMux I__8751 (
            .O(N__40031),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    CascadeMux I__8750 (
            .O(N__40028),
            .I(N__40025));
    InMux I__8749 (
            .O(N__40025),
            .I(N__40022));
    LocalMux I__8748 (
            .O(N__40022),
            .I(N__40017));
    InMux I__8747 (
            .O(N__40021),
            .I(N__40013));
    InMux I__8746 (
            .O(N__40020),
            .I(N__40010));
    Sp12to4 I__8745 (
            .O(N__40017),
            .I(N__40007));
    InMux I__8744 (
            .O(N__40016),
            .I(N__40004));
    LocalMux I__8743 (
            .O(N__40013),
            .I(N__40001));
    LocalMux I__8742 (
            .O(N__40010),
            .I(N__39994));
    Span12Mux_h I__8741 (
            .O(N__40007),
            .I(N__39994));
    LocalMux I__8740 (
            .O(N__40004),
            .I(N__39994));
    Span4Mux_v I__8739 (
            .O(N__40001),
            .I(N__39991));
    Odrv12 I__8738 (
            .O(N__39994),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__8737 (
            .O(N__39991),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    InMux I__8736 (
            .O(N__39986),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    InMux I__8735 (
            .O(N__39983),
            .I(N__39980));
    LocalMux I__8734 (
            .O(N__39980),
            .I(N__39976));
    InMux I__8733 (
            .O(N__39979),
            .I(N__39973));
    Sp12to4 I__8732 (
            .O(N__39976),
            .I(N__39970));
    LocalMux I__8731 (
            .O(N__39973),
            .I(N__39967));
    Span12Mux_v I__8730 (
            .O(N__39970),
            .I(N__39962));
    Span4Mux_h I__8729 (
            .O(N__39967),
            .I(N__39959));
    InMux I__8728 (
            .O(N__39966),
            .I(N__39956));
    InMux I__8727 (
            .O(N__39965),
            .I(N__39953));
    Span12Mux_h I__8726 (
            .O(N__39962),
            .I(N__39946));
    Sp12to4 I__8725 (
            .O(N__39959),
            .I(N__39946));
    LocalMux I__8724 (
            .O(N__39956),
            .I(N__39946));
    LocalMux I__8723 (
            .O(N__39953),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv12 I__8722 (
            .O(N__39946),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    InMux I__8721 (
            .O(N__39941),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    CascadeMux I__8720 (
            .O(N__39938),
            .I(N__39935));
    InMux I__8719 (
            .O(N__39935),
            .I(N__39932));
    LocalMux I__8718 (
            .O(N__39932),
            .I(N__39929));
    Span4Mux_v I__8717 (
            .O(N__39929),
            .I(N__39926));
    Span4Mux_h I__8716 (
            .O(N__39926),
            .I(N__39922));
    InMux I__8715 (
            .O(N__39925),
            .I(N__39917));
    Sp12to4 I__8714 (
            .O(N__39922),
            .I(N__39914));
    InMux I__8713 (
            .O(N__39921),
            .I(N__39911));
    InMux I__8712 (
            .O(N__39920),
            .I(N__39908));
    LocalMux I__8711 (
            .O(N__39917),
            .I(N__39901));
    Span12Mux_h I__8710 (
            .O(N__39914),
            .I(N__39901));
    LocalMux I__8709 (
            .O(N__39911),
            .I(N__39901));
    LocalMux I__8708 (
            .O(N__39908),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv12 I__8707 (
            .O(N__39901),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    InMux I__8706 (
            .O(N__39896),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ));
    InMux I__8705 (
            .O(N__39893),
            .I(N__39889));
    InMux I__8704 (
            .O(N__39892),
            .I(N__39886));
    LocalMux I__8703 (
            .O(N__39889),
            .I(N__39881));
    LocalMux I__8702 (
            .O(N__39886),
            .I(N__39881));
    Odrv12 I__8701 (
            .O(N__39881),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    CascadeMux I__8700 (
            .O(N__39878),
            .I(N__39874));
    CascadeMux I__8699 (
            .O(N__39877),
            .I(N__39870));
    InMux I__8698 (
            .O(N__39874),
            .I(N__39867));
    InMux I__8697 (
            .O(N__39873),
            .I(N__39864));
    InMux I__8696 (
            .O(N__39870),
            .I(N__39861));
    LocalMux I__8695 (
            .O(N__39867),
            .I(N__39858));
    LocalMux I__8694 (
            .O(N__39864),
            .I(N__39854));
    LocalMux I__8693 (
            .O(N__39861),
            .I(N__39851));
    Span4Mux_v I__8692 (
            .O(N__39858),
            .I(N__39848));
    CascadeMux I__8691 (
            .O(N__39857),
            .I(N__39845));
    Span4Mux_v I__8690 (
            .O(N__39854),
            .I(N__39842));
    Span4Mux_v I__8689 (
            .O(N__39851),
            .I(N__39839));
    Span4Mux_h I__8688 (
            .O(N__39848),
            .I(N__39836));
    InMux I__8687 (
            .O(N__39845),
            .I(N__39832));
    Sp12to4 I__8686 (
            .O(N__39842),
            .I(N__39825));
    Sp12to4 I__8685 (
            .O(N__39839),
            .I(N__39825));
    Sp12to4 I__8684 (
            .O(N__39836),
            .I(N__39825));
    InMux I__8683 (
            .O(N__39835),
            .I(N__39822));
    LocalMux I__8682 (
            .O(N__39832),
            .I(N__39819));
    Span12Mux_h I__8681 (
            .O(N__39825),
            .I(N__39816));
    LocalMux I__8680 (
            .O(N__39822),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__8679 (
            .O(N__39819),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv12 I__8678 (
            .O(N__39816),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    InMux I__8677 (
            .O(N__39809),
            .I(N__39806));
    LocalMux I__8676 (
            .O(N__39806),
            .I(N__39803));
    Odrv12 I__8675 (
            .O(N__39803),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ));
    CascadeMux I__8674 (
            .O(N__39800),
            .I(N__39797));
    InMux I__8673 (
            .O(N__39797),
            .I(N__39793));
    InMux I__8672 (
            .O(N__39796),
            .I(N__39790));
    LocalMux I__8671 (
            .O(N__39793),
            .I(N__39787));
    LocalMux I__8670 (
            .O(N__39790),
            .I(N__39781));
    Span12Mux_h I__8669 (
            .O(N__39787),
            .I(N__39781));
    InMux I__8668 (
            .O(N__39786),
            .I(N__39778));
    Odrv12 I__8667 (
            .O(N__39781),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    LocalMux I__8666 (
            .O(N__39778),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    InMux I__8665 (
            .O(N__39773),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ));
    InMux I__8664 (
            .O(N__39770),
            .I(N__39767));
    LocalMux I__8663 (
            .O(N__39767),
            .I(N__39764));
    Span4Mux_v I__8662 (
            .O(N__39764),
            .I(N__39761));
    Odrv4 I__8661 (
            .O(N__39761),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ));
    CascadeMux I__8660 (
            .O(N__39758),
            .I(N__39755));
    InMux I__8659 (
            .O(N__39755),
            .I(N__39752));
    LocalMux I__8658 (
            .O(N__39752),
            .I(N__39749));
    Span4Mux_v I__8657 (
            .O(N__39749),
            .I(N__39744));
    InMux I__8656 (
            .O(N__39748),
            .I(N__39741));
    InMux I__8655 (
            .O(N__39747),
            .I(N__39738));
    Span4Mux_h I__8654 (
            .O(N__39744),
            .I(N__39735));
    LocalMux I__8653 (
            .O(N__39741),
            .I(N__39730));
    LocalMux I__8652 (
            .O(N__39738),
            .I(N__39730));
    Sp12to4 I__8651 (
            .O(N__39735),
            .I(N__39726));
    Span12Mux_v I__8650 (
            .O(N__39730),
            .I(N__39723));
    InMux I__8649 (
            .O(N__39729),
            .I(N__39720));
    Span12Mux_v I__8648 (
            .O(N__39726),
            .I(N__39717));
    Odrv12 I__8647 (
            .O(N__39723),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    LocalMux I__8646 (
            .O(N__39720),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv12 I__8645 (
            .O(N__39717),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    InMux I__8644 (
            .O(N__39710),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ));
    InMux I__8643 (
            .O(N__39707),
            .I(N__39704));
    LocalMux I__8642 (
            .O(N__39704),
            .I(N__39701));
    Span4Mux_h I__8641 (
            .O(N__39701),
            .I(N__39698));
    Odrv4 I__8640 (
            .O(N__39698),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    CascadeMux I__8639 (
            .O(N__39695),
            .I(N__39691));
    InMux I__8638 (
            .O(N__39694),
            .I(N__39687));
    InMux I__8637 (
            .O(N__39691),
            .I(N__39684));
    InMux I__8636 (
            .O(N__39690),
            .I(N__39681));
    LocalMux I__8635 (
            .O(N__39687),
            .I(N__39678));
    LocalMux I__8634 (
            .O(N__39684),
            .I(N__39675));
    LocalMux I__8633 (
            .O(N__39681),
            .I(N__39670));
    Span4Mux_v I__8632 (
            .O(N__39678),
            .I(N__39670));
    Span4Mux_v I__8631 (
            .O(N__39675),
            .I(N__39667));
    Sp12to4 I__8630 (
            .O(N__39670),
            .I(N__39661));
    Sp12to4 I__8629 (
            .O(N__39667),
            .I(N__39661));
    InMux I__8628 (
            .O(N__39666),
            .I(N__39658));
    Span12Mux_h I__8627 (
            .O(N__39661),
            .I(N__39655));
    LocalMux I__8626 (
            .O(N__39658),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv12 I__8625 (
            .O(N__39655),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    InMux I__8624 (
            .O(N__39650),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ));
    InMux I__8623 (
            .O(N__39647),
            .I(N__39642));
    InMux I__8622 (
            .O(N__39646),
            .I(N__39639));
    InMux I__8621 (
            .O(N__39645),
            .I(N__39635));
    LocalMux I__8620 (
            .O(N__39642),
            .I(N__39632));
    LocalMux I__8619 (
            .O(N__39639),
            .I(N__39629));
    InMux I__8618 (
            .O(N__39638),
            .I(N__39626));
    LocalMux I__8617 (
            .O(N__39635),
            .I(N__39621));
    Span4Mux_v I__8616 (
            .O(N__39632),
            .I(N__39621));
    Span12Mux_v I__8615 (
            .O(N__39629),
            .I(N__39618));
    LocalMux I__8614 (
            .O(N__39626),
            .I(N__39615));
    Span4Mux_v I__8613 (
            .O(N__39621),
            .I(N__39612));
    Odrv12 I__8612 (
            .O(N__39618),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__8611 (
            .O(N__39615),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__8610 (
            .O(N__39612),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    CascadeMux I__8609 (
            .O(N__39605),
            .I(N__39602));
    InMux I__8608 (
            .O(N__39602),
            .I(N__39599));
    LocalMux I__8607 (
            .O(N__39599),
            .I(N__39596));
    Odrv4 I__8606 (
            .O(N__39596),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    InMux I__8605 (
            .O(N__39593),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    InMux I__8604 (
            .O(N__39590),
            .I(N__39587));
    LocalMux I__8603 (
            .O(N__39587),
            .I(N__39584));
    Odrv4 I__8602 (
            .O(N__39584),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    CascadeMux I__8601 (
            .O(N__39581),
            .I(N__39577));
    CascadeMux I__8600 (
            .O(N__39580),
            .I(N__39574));
    InMux I__8599 (
            .O(N__39577),
            .I(N__39570));
    InMux I__8598 (
            .O(N__39574),
            .I(N__39567));
    InMux I__8597 (
            .O(N__39573),
            .I(N__39564));
    LocalMux I__8596 (
            .O(N__39570),
            .I(N__39561));
    LocalMux I__8595 (
            .O(N__39567),
            .I(N__39558));
    LocalMux I__8594 (
            .O(N__39564),
            .I(N__39550));
    Sp12to4 I__8593 (
            .O(N__39561),
            .I(N__39550));
    Span12Mux_h I__8592 (
            .O(N__39558),
            .I(N__39550));
    InMux I__8591 (
            .O(N__39557),
            .I(N__39547));
    Odrv12 I__8590 (
            .O(N__39550),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    LocalMux I__8589 (
            .O(N__39547),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    InMux I__8588 (
            .O(N__39542),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    InMux I__8587 (
            .O(N__39539),
            .I(N__39536));
    LocalMux I__8586 (
            .O(N__39536),
            .I(N__39533));
    Odrv12 I__8585 (
            .O(N__39533),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    CascadeMux I__8584 (
            .O(N__39530),
            .I(N__39527));
    InMux I__8583 (
            .O(N__39527),
            .I(N__39524));
    LocalMux I__8582 (
            .O(N__39524),
            .I(N__39520));
    InMux I__8581 (
            .O(N__39523),
            .I(N__39516));
    Sp12to4 I__8580 (
            .O(N__39520),
            .I(N__39513));
    InMux I__8579 (
            .O(N__39519),
            .I(N__39509));
    LocalMux I__8578 (
            .O(N__39516),
            .I(N__39506));
    Span12Mux_v I__8577 (
            .O(N__39513),
            .I(N__39503));
    InMux I__8576 (
            .O(N__39512),
            .I(N__39500));
    LocalMux I__8575 (
            .O(N__39509),
            .I(N__39495));
    Span12Mux_s11_v I__8574 (
            .O(N__39506),
            .I(N__39495));
    Odrv12 I__8573 (
            .O(N__39503),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    LocalMux I__8572 (
            .O(N__39500),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv12 I__8571 (
            .O(N__39495),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    InMux I__8570 (
            .O(N__39488),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    InMux I__8569 (
            .O(N__39485),
            .I(N__39482));
    LocalMux I__8568 (
            .O(N__39482),
            .I(N__39479));
    Odrv4 I__8567 (
            .O(N__39479),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    CascadeMux I__8566 (
            .O(N__39476),
            .I(N__39473));
    InMux I__8565 (
            .O(N__39473),
            .I(N__39468));
    InMux I__8564 (
            .O(N__39472),
            .I(N__39465));
    InMux I__8563 (
            .O(N__39471),
            .I(N__39462));
    LocalMux I__8562 (
            .O(N__39468),
            .I(N__39459));
    LocalMux I__8561 (
            .O(N__39465),
            .I(N__39453));
    LocalMux I__8560 (
            .O(N__39462),
            .I(N__39453));
    Span12Mux_v I__8559 (
            .O(N__39459),
            .I(N__39450));
    InMux I__8558 (
            .O(N__39458),
            .I(N__39447));
    Span12Mux_v I__8557 (
            .O(N__39453),
            .I(N__39444));
    Odrv12 I__8556 (
            .O(N__39450),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    LocalMux I__8555 (
            .O(N__39447),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv12 I__8554 (
            .O(N__39444),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    InMux I__8553 (
            .O(N__39437),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ));
    InMux I__8552 (
            .O(N__39434),
            .I(N__39430));
    InMux I__8551 (
            .O(N__39433),
            .I(N__39427));
    LocalMux I__8550 (
            .O(N__39430),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    LocalMux I__8549 (
            .O(N__39427),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CascadeMux I__8548 (
            .O(N__39422),
            .I(N__39419));
    InMux I__8547 (
            .O(N__39419),
            .I(N__39414));
    InMux I__8546 (
            .O(N__39418),
            .I(N__39411));
    InMux I__8545 (
            .O(N__39417),
            .I(N__39408));
    LocalMux I__8544 (
            .O(N__39414),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    LocalMux I__8543 (
            .O(N__39411),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    LocalMux I__8542 (
            .O(N__39408),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__8541 (
            .O(N__39401),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__8540 (
            .O(N__39398),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__8539 (
            .O(N__39395),
            .I(N__39392));
    LocalMux I__8538 (
            .O(N__39392),
            .I(\phase_controller_inst1.start_timer_hc_0_sqmuxa ));
    InMux I__8537 (
            .O(N__39389),
            .I(N__39385));
    InMux I__8536 (
            .O(N__39388),
            .I(N__39382));
    LocalMux I__8535 (
            .O(N__39385),
            .I(N__39379));
    LocalMux I__8534 (
            .O(N__39382),
            .I(N__39376));
    Span4Mux_s3_h I__8533 (
            .O(N__39379),
            .I(N__39373));
    Span12Mux_h I__8532 (
            .O(N__39376),
            .I(N__39370));
    Span4Mux_h I__8531 (
            .O(N__39373),
            .I(N__39367));
    Odrv12 I__8530 (
            .O(N__39370),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    Odrv4 I__8529 (
            .O(N__39367),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    IoInMux I__8528 (
            .O(N__39362),
            .I(N__39359));
    LocalMux I__8527 (
            .O(N__39359),
            .I(N__39356));
    IoSpan4Mux I__8526 (
            .O(N__39356),
            .I(N__39353));
    Sp12to4 I__8525 (
            .O(N__39353),
            .I(N__39348));
    InMux I__8524 (
            .O(N__39352),
            .I(N__39345));
    InMux I__8523 (
            .O(N__39351),
            .I(N__39342));
    Odrv12 I__8522 (
            .O(N__39348),
            .I(s1_phy_c));
    LocalMux I__8521 (
            .O(N__39345),
            .I(s1_phy_c));
    LocalMux I__8520 (
            .O(N__39342),
            .I(s1_phy_c));
    InMux I__8519 (
            .O(N__39335),
            .I(N__39329));
    InMux I__8518 (
            .O(N__39334),
            .I(N__39324));
    InMux I__8517 (
            .O(N__39333),
            .I(N__39324));
    InMux I__8516 (
            .O(N__39332),
            .I(N__39321));
    LocalMux I__8515 (
            .O(N__39329),
            .I(N__39318));
    LocalMux I__8514 (
            .O(N__39324),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__8513 (
            .O(N__39321),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    Odrv4 I__8512 (
            .O(N__39318),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    InMux I__8511 (
            .O(N__39311),
            .I(N__39303));
    InMux I__8510 (
            .O(N__39310),
            .I(N__39300));
    InMux I__8509 (
            .O(N__39309),
            .I(N__39295));
    InMux I__8508 (
            .O(N__39308),
            .I(N__39295));
    InMux I__8507 (
            .O(N__39307),
            .I(N__39289));
    InMux I__8506 (
            .O(N__39306),
            .I(N__39289));
    LocalMux I__8505 (
            .O(N__39303),
            .I(N__39282));
    LocalMux I__8504 (
            .O(N__39300),
            .I(N__39282));
    LocalMux I__8503 (
            .O(N__39295),
            .I(N__39282));
    InMux I__8502 (
            .O(N__39294),
            .I(N__39279));
    LocalMux I__8501 (
            .O(N__39289),
            .I(state_3));
    Odrv4 I__8500 (
            .O(N__39282),
            .I(state_3));
    LocalMux I__8499 (
            .O(N__39279),
            .I(state_3));
    IoInMux I__8498 (
            .O(N__39272),
            .I(N__39269));
    LocalMux I__8497 (
            .O(N__39269),
            .I(N__39266));
    Span4Mux_s1_v I__8496 (
            .O(N__39266),
            .I(N__39263));
    Span4Mux_h I__8495 (
            .O(N__39263),
            .I(N__39260));
    Span4Mux_v I__8494 (
            .O(N__39260),
            .I(N__39256));
    InMux I__8493 (
            .O(N__39259),
            .I(N__39253));
    Odrv4 I__8492 (
            .O(N__39256),
            .I(T01_c));
    LocalMux I__8491 (
            .O(N__39253),
            .I(T01_c));
    CascadeMux I__8490 (
            .O(N__39248),
            .I(N__39245));
    InMux I__8489 (
            .O(N__39245),
            .I(N__39240));
    InMux I__8488 (
            .O(N__39244),
            .I(N__39237));
    InMux I__8487 (
            .O(N__39243),
            .I(N__39234));
    LocalMux I__8486 (
            .O(N__39240),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    LocalMux I__8485 (
            .O(N__39237),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    LocalMux I__8484 (
            .O(N__39234),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__8483 (
            .O(N__39227),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__8482 (
            .O(N__39224),
            .I(N__39221));
    InMux I__8481 (
            .O(N__39221),
            .I(N__39216));
    InMux I__8480 (
            .O(N__39220),
            .I(N__39213));
    InMux I__8479 (
            .O(N__39219),
            .I(N__39210));
    LocalMux I__8478 (
            .O(N__39216),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    LocalMux I__8477 (
            .O(N__39213),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    LocalMux I__8476 (
            .O(N__39210),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__8475 (
            .O(N__39203),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__8474 (
            .O(N__39200),
            .I(N__39197));
    InMux I__8473 (
            .O(N__39197),
            .I(N__39192));
    InMux I__8472 (
            .O(N__39196),
            .I(N__39189));
    InMux I__8471 (
            .O(N__39195),
            .I(N__39186));
    LocalMux I__8470 (
            .O(N__39192),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    LocalMux I__8469 (
            .O(N__39189),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    LocalMux I__8468 (
            .O(N__39186),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__8467 (
            .O(N__39179),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__8466 (
            .O(N__39176),
            .I(N__39173));
    InMux I__8465 (
            .O(N__39173),
            .I(N__39168));
    InMux I__8464 (
            .O(N__39172),
            .I(N__39165));
    InMux I__8463 (
            .O(N__39171),
            .I(N__39162));
    LocalMux I__8462 (
            .O(N__39168),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__8461 (
            .O(N__39165),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__8460 (
            .O(N__39162),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__8459 (
            .O(N__39155),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__8458 (
            .O(N__39152),
            .I(N__39149));
    InMux I__8457 (
            .O(N__39149),
            .I(N__39144));
    InMux I__8456 (
            .O(N__39148),
            .I(N__39141));
    InMux I__8455 (
            .O(N__39147),
            .I(N__39138));
    LocalMux I__8454 (
            .O(N__39144),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__8453 (
            .O(N__39141),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__8452 (
            .O(N__39138),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__8451 (
            .O(N__39131),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__8450 (
            .O(N__39128),
            .I(N__39125));
    InMux I__8449 (
            .O(N__39125),
            .I(N__39120));
    InMux I__8448 (
            .O(N__39124),
            .I(N__39117));
    InMux I__8447 (
            .O(N__39123),
            .I(N__39114));
    LocalMux I__8446 (
            .O(N__39120),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__8445 (
            .O(N__39117),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__8444 (
            .O(N__39114),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__8443 (
            .O(N__39107),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__8442 (
            .O(N__39104),
            .I(N__39101));
    InMux I__8441 (
            .O(N__39101),
            .I(N__39096));
    InMux I__8440 (
            .O(N__39100),
            .I(N__39093));
    InMux I__8439 (
            .O(N__39099),
            .I(N__39090));
    LocalMux I__8438 (
            .O(N__39096),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__8437 (
            .O(N__39093),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__8436 (
            .O(N__39090),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__8435 (
            .O(N__39083),
            .I(bfn_15_17_0_));
    CascadeMux I__8434 (
            .O(N__39080),
            .I(N__39077));
    InMux I__8433 (
            .O(N__39077),
            .I(N__39072));
    InMux I__8432 (
            .O(N__39076),
            .I(N__39069));
    InMux I__8431 (
            .O(N__39075),
            .I(N__39066));
    LocalMux I__8430 (
            .O(N__39072),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__8429 (
            .O(N__39069),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__8428 (
            .O(N__39066),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    InMux I__8427 (
            .O(N__39059),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__8426 (
            .O(N__39056),
            .I(N__39051));
    InMux I__8425 (
            .O(N__39055),
            .I(N__39046));
    InMux I__8424 (
            .O(N__39054),
            .I(N__39046));
    LocalMux I__8423 (
            .O(N__39051),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    LocalMux I__8422 (
            .O(N__39046),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    CascadeMux I__8421 (
            .O(N__39041),
            .I(N__39037));
    InMux I__8420 (
            .O(N__39040),
            .I(N__39034));
    InMux I__8419 (
            .O(N__39037),
            .I(N__39031));
    LocalMux I__8418 (
            .O(N__39034),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    LocalMux I__8417 (
            .O(N__39031),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    InMux I__8416 (
            .O(N__39026),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__8415 (
            .O(N__39023),
            .I(N__39018));
    InMux I__8414 (
            .O(N__39022),
            .I(N__39013));
    InMux I__8413 (
            .O(N__39021),
            .I(N__39013));
    LocalMux I__8412 (
            .O(N__39018),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    LocalMux I__8411 (
            .O(N__39013),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__8410 (
            .O(N__39008),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__8409 (
            .O(N__39005),
            .I(N__39002));
    InMux I__8408 (
            .O(N__39002),
            .I(N__38997));
    InMux I__8407 (
            .O(N__39001),
            .I(N__38994));
    InMux I__8406 (
            .O(N__39000),
            .I(N__38991));
    LocalMux I__8405 (
            .O(N__38997),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    LocalMux I__8404 (
            .O(N__38994),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    LocalMux I__8403 (
            .O(N__38991),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__8402 (
            .O(N__38984),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__8401 (
            .O(N__38981),
            .I(N__38976));
    CascadeMux I__8400 (
            .O(N__38980),
            .I(N__38973));
    InMux I__8399 (
            .O(N__38979),
            .I(N__38970));
    InMux I__8398 (
            .O(N__38976),
            .I(N__38965));
    InMux I__8397 (
            .O(N__38973),
            .I(N__38965));
    LocalMux I__8396 (
            .O(N__38970),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    LocalMux I__8395 (
            .O(N__38965),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__8394 (
            .O(N__38960),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__8393 (
            .O(N__38957),
            .I(N__38954));
    InMux I__8392 (
            .O(N__38954),
            .I(N__38949));
    InMux I__8391 (
            .O(N__38953),
            .I(N__38946));
    InMux I__8390 (
            .O(N__38952),
            .I(N__38943));
    LocalMux I__8389 (
            .O(N__38949),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__8388 (
            .O(N__38946),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__8387 (
            .O(N__38943),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__8386 (
            .O(N__38936),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__8385 (
            .O(N__38933),
            .I(N__38930));
    InMux I__8384 (
            .O(N__38930),
            .I(N__38925));
    InMux I__8383 (
            .O(N__38929),
            .I(N__38922));
    InMux I__8382 (
            .O(N__38928),
            .I(N__38919));
    LocalMux I__8381 (
            .O(N__38925),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__8380 (
            .O(N__38922),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__8379 (
            .O(N__38919),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__8378 (
            .O(N__38912),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__8377 (
            .O(N__38909),
            .I(N__38906));
    InMux I__8376 (
            .O(N__38906),
            .I(N__38901));
    InMux I__8375 (
            .O(N__38905),
            .I(N__38898));
    InMux I__8374 (
            .O(N__38904),
            .I(N__38895));
    LocalMux I__8373 (
            .O(N__38901),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__8372 (
            .O(N__38898),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__8371 (
            .O(N__38895),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__8370 (
            .O(N__38888),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__8369 (
            .O(N__38885),
            .I(N__38882));
    InMux I__8368 (
            .O(N__38882),
            .I(N__38877));
    InMux I__8367 (
            .O(N__38881),
            .I(N__38874));
    InMux I__8366 (
            .O(N__38880),
            .I(N__38871));
    LocalMux I__8365 (
            .O(N__38877),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__8364 (
            .O(N__38874),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__8363 (
            .O(N__38871),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__8362 (
            .O(N__38864),
            .I(bfn_15_16_0_));
    CascadeMux I__8361 (
            .O(N__38861),
            .I(N__38858));
    InMux I__8360 (
            .O(N__38858),
            .I(N__38853));
    InMux I__8359 (
            .O(N__38857),
            .I(N__38850));
    InMux I__8358 (
            .O(N__38856),
            .I(N__38847));
    LocalMux I__8357 (
            .O(N__38853),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__8356 (
            .O(N__38850),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__8355 (
            .O(N__38847),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__8354 (
            .O(N__38840),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__8353 (
            .O(N__38837),
            .I(N__38834));
    InMux I__8352 (
            .O(N__38834),
            .I(N__38829));
    InMux I__8351 (
            .O(N__38833),
            .I(N__38826));
    InMux I__8350 (
            .O(N__38832),
            .I(N__38823));
    LocalMux I__8349 (
            .O(N__38829),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    LocalMux I__8348 (
            .O(N__38826),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    LocalMux I__8347 (
            .O(N__38823),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__8346 (
            .O(N__38816),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__8345 (
            .O(N__38813),
            .I(N__38810));
    InMux I__8344 (
            .O(N__38810),
            .I(N__38805));
    InMux I__8343 (
            .O(N__38809),
            .I(N__38802));
    InMux I__8342 (
            .O(N__38808),
            .I(N__38799));
    LocalMux I__8341 (
            .O(N__38805),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    LocalMux I__8340 (
            .O(N__38802),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    LocalMux I__8339 (
            .O(N__38799),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__8338 (
            .O(N__38792),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__8337 (
            .O(N__38789),
            .I(N__38786));
    InMux I__8336 (
            .O(N__38786),
            .I(N__38781));
    InMux I__8335 (
            .O(N__38785),
            .I(N__38778));
    InMux I__8334 (
            .O(N__38784),
            .I(N__38775));
    LocalMux I__8333 (
            .O(N__38781),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    LocalMux I__8332 (
            .O(N__38778),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    LocalMux I__8331 (
            .O(N__38775),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__8330 (
            .O(N__38768),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__8329 (
            .O(N__38765),
            .I(N__38762));
    InMux I__8328 (
            .O(N__38762),
            .I(N__38757));
    InMux I__8327 (
            .O(N__38761),
            .I(N__38754));
    InMux I__8326 (
            .O(N__38760),
            .I(N__38751));
    LocalMux I__8325 (
            .O(N__38757),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__8324 (
            .O(N__38754),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__8323 (
            .O(N__38751),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__8322 (
            .O(N__38744),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__8321 (
            .O(N__38741),
            .I(N__38738));
    InMux I__8320 (
            .O(N__38738),
            .I(N__38733));
    InMux I__8319 (
            .O(N__38737),
            .I(N__38730));
    InMux I__8318 (
            .O(N__38736),
            .I(N__38727));
    LocalMux I__8317 (
            .O(N__38733),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__8316 (
            .O(N__38730),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__8315 (
            .O(N__38727),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__8314 (
            .O(N__38720),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__8313 (
            .O(N__38717),
            .I(N__38714));
    InMux I__8312 (
            .O(N__38714),
            .I(N__38709));
    InMux I__8311 (
            .O(N__38713),
            .I(N__38706));
    InMux I__8310 (
            .O(N__38712),
            .I(N__38703));
    LocalMux I__8309 (
            .O(N__38709),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__8308 (
            .O(N__38706),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__8307 (
            .O(N__38703),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__8306 (
            .O(N__38696),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__8305 (
            .O(N__38693),
            .I(N__38690));
    InMux I__8304 (
            .O(N__38690),
            .I(N__38685));
    InMux I__8303 (
            .O(N__38689),
            .I(N__38682));
    InMux I__8302 (
            .O(N__38688),
            .I(N__38679));
    LocalMux I__8301 (
            .O(N__38685),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__8300 (
            .O(N__38682),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__8299 (
            .O(N__38679),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__8298 (
            .O(N__38672),
            .I(bfn_15_15_0_));
    CascadeMux I__8297 (
            .O(N__38669),
            .I(N__38666));
    InMux I__8296 (
            .O(N__38666),
            .I(N__38661));
    InMux I__8295 (
            .O(N__38665),
            .I(N__38658));
    InMux I__8294 (
            .O(N__38664),
            .I(N__38655));
    LocalMux I__8293 (
            .O(N__38661),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__8292 (
            .O(N__38658),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__8291 (
            .O(N__38655),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__8290 (
            .O(N__38648),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__8289 (
            .O(N__38645),
            .I(N__38642));
    InMux I__8288 (
            .O(N__38642),
            .I(N__38636));
    InMux I__8287 (
            .O(N__38641),
            .I(N__38636));
    LocalMux I__8286 (
            .O(N__38636),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ));
    CascadeMux I__8285 (
            .O(N__38633),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12_cascade_));
    InMux I__8284 (
            .O(N__38630),
            .I(N__38627));
    LocalMux I__8283 (
            .O(N__38627),
            .I(N__38624));
    Span4Mux_v I__8282 (
            .O(N__38624),
            .I(N__38621));
    Odrv4 I__8281 (
            .O(N__38621),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ));
    InMux I__8280 (
            .O(N__38618),
            .I(N__38615));
    LocalMux I__8279 (
            .O(N__38615),
            .I(N__38612));
    Span4Mux_v I__8278 (
            .O(N__38612),
            .I(N__38609));
    Odrv4 I__8277 (
            .O(N__38609),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ));
    InMux I__8276 (
            .O(N__38606),
            .I(N__38600));
    InMux I__8275 (
            .O(N__38605),
            .I(N__38600));
    LocalMux I__8274 (
            .O(N__38600),
            .I(N__38597));
    Span4Mux_h I__8273 (
            .O(N__38597),
            .I(N__38594));
    Odrv4 I__8272 (
            .O(N__38594),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ));
    InMux I__8271 (
            .O(N__38591),
            .I(N__38588));
    LocalMux I__8270 (
            .O(N__38588),
            .I(N__38585));
    Span4Mux_h I__8269 (
            .O(N__38585),
            .I(N__38581));
    InMux I__8268 (
            .O(N__38584),
            .I(N__38578));
    Odrv4 I__8267 (
            .O(N__38581),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13));
    LocalMux I__8266 (
            .O(N__38578),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13));
    InMux I__8265 (
            .O(N__38573),
            .I(N__38570));
    LocalMux I__8264 (
            .O(N__38570),
            .I(N__38566));
    CascadeMux I__8263 (
            .O(N__38569),
            .I(N__38563));
    Span4Mux_h I__8262 (
            .O(N__38566),
            .I(N__38559));
    InMux I__8261 (
            .O(N__38563),
            .I(N__38556));
    InMux I__8260 (
            .O(N__38562),
            .I(N__38553));
    Odrv4 I__8259 (
            .O(N__38559),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__8258 (
            .O(N__38556),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__8257 (
            .O(N__38553),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    InMux I__8256 (
            .O(N__38546),
            .I(N__38543));
    LocalMux I__8255 (
            .O(N__38543),
            .I(N__38539));
    CascadeMux I__8254 (
            .O(N__38542),
            .I(N__38536));
    Span4Mux_v I__8253 (
            .O(N__38539),
            .I(N__38532));
    InMux I__8252 (
            .O(N__38536),
            .I(N__38529));
    InMux I__8251 (
            .O(N__38535),
            .I(N__38526));
    Odrv4 I__8250 (
            .O(N__38532),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__8249 (
            .O(N__38529),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__8248 (
            .O(N__38526),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    InMux I__8247 (
            .O(N__38519),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__8246 (
            .O(N__38516),
            .I(N__38513));
    LocalMux I__8245 (
            .O(N__38513),
            .I(N__38510));
    Span4Mux_h I__8244 (
            .O(N__38510),
            .I(N__38507));
    Odrv4 I__8243 (
            .O(N__38507),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt20 ));
    CascadeMux I__8242 (
            .O(N__38504),
            .I(N__38499));
    InMux I__8241 (
            .O(N__38503),
            .I(N__38496));
    InMux I__8240 (
            .O(N__38502),
            .I(N__38491));
    InMux I__8239 (
            .O(N__38499),
            .I(N__38491));
    LocalMux I__8238 (
            .O(N__38496),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ));
    LocalMux I__8237 (
            .O(N__38491),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ));
    CascadeMux I__8236 (
            .O(N__38486),
            .I(N__38481));
    InMux I__8235 (
            .O(N__38485),
            .I(N__38478));
    InMux I__8234 (
            .O(N__38484),
            .I(N__38473));
    InMux I__8233 (
            .O(N__38481),
            .I(N__38473));
    LocalMux I__8232 (
            .O(N__38478),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ));
    LocalMux I__8231 (
            .O(N__38473),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ));
    CascadeMux I__8230 (
            .O(N__38468),
            .I(N__38465));
    InMux I__8229 (
            .O(N__38465),
            .I(N__38462));
    LocalMux I__8228 (
            .O(N__38462),
            .I(N__38459));
    Span4Mux_h I__8227 (
            .O(N__38459),
            .I(N__38456));
    Odrv4 I__8226 (
            .O(N__38456),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ));
    InMux I__8225 (
            .O(N__38453),
            .I(N__38447));
    InMux I__8224 (
            .O(N__38452),
            .I(N__38447));
    LocalMux I__8223 (
            .O(N__38447),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ));
    InMux I__8222 (
            .O(N__38444),
            .I(N__38438));
    InMux I__8221 (
            .O(N__38443),
            .I(N__38438));
    LocalMux I__8220 (
            .O(N__38438),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ));
    InMux I__8219 (
            .O(N__38435),
            .I(N__38432));
    LocalMux I__8218 (
            .O(N__38432),
            .I(N__38429));
    Span4Mux_h I__8217 (
            .O(N__38429),
            .I(N__38426));
    Odrv4 I__8216 (
            .O(N__38426),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ));
    CascadeMux I__8215 (
            .O(N__38423),
            .I(N__38420));
    InMux I__8214 (
            .O(N__38420),
            .I(N__38417));
    LocalMux I__8213 (
            .O(N__38417),
            .I(N__38414));
    Span4Mux_h I__8212 (
            .O(N__38414),
            .I(N__38411));
    Odrv4 I__8211 (
            .O(N__38411),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt22 ));
    InMux I__8210 (
            .O(N__38408),
            .I(N__38403));
    InMux I__8209 (
            .O(N__38407),
            .I(N__38400));
    InMux I__8208 (
            .O(N__38406),
            .I(N__38397));
    LocalMux I__8207 (
            .O(N__38403),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ));
    LocalMux I__8206 (
            .O(N__38400),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ));
    LocalMux I__8205 (
            .O(N__38397),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ));
    CascadeMux I__8204 (
            .O(N__38390),
            .I(N__38386));
    InMux I__8203 (
            .O(N__38389),
            .I(N__38382));
    InMux I__8202 (
            .O(N__38386),
            .I(N__38379));
    InMux I__8201 (
            .O(N__38385),
            .I(N__38376));
    LocalMux I__8200 (
            .O(N__38382),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ));
    LocalMux I__8199 (
            .O(N__38379),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ));
    LocalMux I__8198 (
            .O(N__38376),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ));
    InMux I__8197 (
            .O(N__38369),
            .I(N__38366));
    LocalMux I__8196 (
            .O(N__38366),
            .I(N__38363));
    Odrv4 I__8195 (
            .O(N__38363),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ));
    InMux I__8194 (
            .O(N__38360),
            .I(N__38354));
    InMux I__8193 (
            .O(N__38359),
            .I(N__38354));
    LocalMux I__8192 (
            .O(N__38354),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ));
    InMux I__8191 (
            .O(N__38351),
            .I(N__38348));
    LocalMux I__8190 (
            .O(N__38348),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ));
    InMux I__8189 (
            .O(N__38345),
            .I(N__38342));
    LocalMux I__8188 (
            .O(N__38342),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ));
    CascadeMux I__8187 (
            .O(N__38339),
            .I(N__38336));
    InMux I__8186 (
            .O(N__38336),
            .I(N__38333));
    LocalMux I__8185 (
            .O(N__38333),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__8184 (
            .O(N__38330),
            .I(N__38327));
    InMux I__8183 (
            .O(N__38327),
            .I(N__38324));
    LocalMux I__8182 (
            .O(N__38324),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt24 ));
    InMux I__8181 (
            .O(N__38321),
            .I(N__38315));
    InMux I__8180 (
            .O(N__38320),
            .I(N__38315));
    LocalMux I__8179 (
            .O(N__38315),
            .I(N__38311));
    InMux I__8178 (
            .O(N__38314),
            .I(N__38308));
    Span4Mux_h I__8177 (
            .O(N__38311),
            .I(N__38305));
    LocalMux I__8176 (
            .O(N__38308),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ));
    Odrv4 I__8175 (
            .O(N__38305),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ));
    CascadeMux I__8174 (
            .O(N__38300),
            .I(N__38297));
    InMux I__8173 (
            .O(N__38297),
            .I(N__38291));
    InMux I__8172 (
            .O(N__38296),
            .I(N__38291));
    LocalMux I__8171 (
            .O(N__38291),
            .I(N__38287));
    InMux I__8170 (
            .O(N__38290),
            .I(N__38284));
    Span4Mux_h I__8169 (
            .O(N__38287),
            .I(N__38281));
    LocalMux I__8168 (
            .O(N__38284),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ));
    Odrv4 I__8167 (
            .O(N__38281),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ));
    InMux I__8166 (
            .O(N__38276),
            .I(N__38273));
    LocalMux I__8165 (
            .O(N__38273),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ));
    InMux I__8164 (
            .O(N__38270),
            .I(\pwm_generator_inst.un3_threshold_cry_19 ));
    InMux I__8163 (
            .O(N__38267),
            .I(N__38264));
    LocalMux I__8162 (
            .O(N__38264),
            .I(\pwm_generator_inst.un3_threshold_cry_19_THRU_CO ));
    InMux I__8161 (
            .O(N__38261),
            .I(N__38257));
    InMux I__8160 (
            .O(N__38260),
            .I(N__38253));
    LocalMux I__8159 (
            .O(N__38257),
            .I(N__38250));
    InMux I__8158 (
            .O(N__38256),
            .I(N__38246));
    LocalMux I__8157 (
            .O(N__38253),
            .I(N__38243));
    Span4Mux_v I__8156 (
            .O(N__38250),
            .I(N__38240));
    InMux I__8155 (
            .O(N__38249),
            .I(N__38237));
    LocalMux I__8154 (
            .O(N__38246),
            .I(N__38234));
    Span4Mux_v I__8153 (
            .O(N__38243),
            .I(N__38231));
    Span4Mux_h I__8152 (
            .O(N__38240),
            .I(N__38228));
    LocalMux I__8151 (
            .O(N__38237),
            .I(N__38225));
    Span4Mux_h I__8150 (
            .O(N__38234),
            .I(N__38222));
    Span4Mux_v I__8149 (
            .O(N__38231),
            .I(N__38219));
    Span4Mux_h I__8148 (
            .O(N__38228),
            .I(N__38216));
    Span4Mux_v I__8147 (
            .O(N__38225),
            .I(N__38213));
    Odrv4 I__8146 (
            .O(N__38222),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    Odrv4 I__8145 (
            .O(N__38219),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    Odrv4 I__8144 (
            .O(N__38216),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    Odrv4 I__8143 (
            .O(N__38213),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    InMux I__8142 (
            .O(N__38204),
            .I(N__38201));
    LocalMux I__8141 (
            .O(N__38201),
            .I(N__38197));
    InMux I__8140 (
            .O(N__38200),
            .I(N__38193));
    Span4Mux_h I__8139 (
            .O(N__38197),
            .I(N__38190));
    InMux I__8138 (
            .O(N__38196),
            .I(N__38187));
    LocalMux I__8137 (
            .O(N__38193),
            .I(N__38184));
    Span4Mux_v I__8136 (
            .O(N__38190),
            .I(N__38181));
    LocalMux I__8135 (
            .O(N__38187),
            .I(N__38176));
    Span4Mux_h I__8134 (
            .O(N__38184),
            .I(N__38176));
    Odrv4 I__8133 (
            .O(N__38181),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    Odrv4 I__8132 (
            .O(N__38176),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    CascadeMux I__8131 (
            .O(N__38171),
            .I(N__38168));
    InMux I__8130 (
            .O(N__38168),
            .I(N__38165));
    LocalMux I__8129 (
            .O(N__38165),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ));
    InMux I__8128 (
            .O(N__38162),
            .I(N__38159));
    LocalMux I__8127 (
            .O(N__38159),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ));
    InMux I__8126 (
            .O(N__38156),
            .I(N__38153));
    LocalMux I__8125 (
            .O(N__38153),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ));
    InMux I__8124 (
            .O(N__38150),
            .I(N__38147));
    LocalMux I__8123 (
            .O(N__38147),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__8122 (
            .O(N__38144),
            .I(N__38141));
    InMux I__8121 (
            .O(N__38141),
            .I(N__38138));
    LocalMux I__8120 (
            .O(N__38138),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt18 ));
    InMux I__8119 (
            .O(N__38135),
            .I(N__38129));
    InMux I__8118 (
            .O(N__38134),
            .I(N__38129));
    LocalMux I__8117 (
            .O(N__38129),
            .I(N__38125));
    InMux I__8116 (
            .O(N__38128),
            .I(N__38122));
    Span4Mux_h I__8115 (
            .O(N__38125),
            .I(N__38119));
    LocalMux I__8114 (
            .O(N__38122),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__8113 (
            .O(N__38119),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    CascadeMux I__8112 (
            .O(N__38114),
            .I(N__38110));
    InMux I__8111 (
            .O(N__38113),
            .I(N__38105));
    InMux I__8110 (
            .O(N__38110),
            .I(N__38105));
    LocalMux I__8109 (
            .O(N__38105),
            .I(N__38102));
    Span4Mux_h I__8108 (
            .O(N__38102),
            .I(N__38099));
    Span4Mux_v I__8107 (
            .O(N__38099),
            .I(N__38096));
    Odrv4 I__8106 (
            .O(N__38096),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ));
    CascadeMux I__8105 (
            .O(N__38093),
            .I(N__38089));
    InMux I__8104 (
            .O(N__38092),
            .I(N__38084));
    InMux I__8103 (
            .O(N__38089),
            .I(N__38084));
    LocalMux I__8102 (
            .O(N__38084),
            .I(N__38080));
    InMux I__8101 (
            .O(N__38083),
            .I(N__38077));
    Span4Mux_h I__8100 (
            .O(N__38080),
            .I(N__38074));
    LocalMux I__8099 (
            .O(N__38077),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__8098 (
            .O(N__38074),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__8097 (
            .O(N__38069),
            .I(N__38066));
    LocalMux I__8096 (
            .O(N__38066),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ));
    InMux I__8095 (
            .O(N__38063),
            .I(N__38060));
    LocalMux I__8094 (
            .O(N__38060),
            .I(\pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ));
    InMux I__8093 (
            .O(N__38057),
            .I(N__38054));
    LocalMux I__8092 (
            .O(N__38054),
            .I(\pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ));
    InMux I__8091 (
            .O(N__38051),
            .I(N__38048));
    LocalMux I__8090 (
            .O(N__38048),
            .I(\pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ));
    InMux I__8089 (
            .O(N__38045),
            .I(N__38042));
    LocalMux I__8088 (
            .O(N__38042),
            .I(\pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ));
    InMux I__8087 (
            .O(N__38039),
            .I(N__38036));
    LocalMux I__8086 (
            .O(N__38036),
            .I(\pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ));
    InMux I__8085 (
            .O(N__38033),
            .I(N__38030));
    LocalMux I__8084 (
            .O(N__38030),
            .I(\pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ));
    InMux I__8083 (
            .O(N__38027),
            .I(N__38024));
    LocalMux I__8082 (
            .O(N__38024),
            .I(\pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ));
    InMux I__8081 (
            .O(N__38021),
            .I(N__38018));
    LocalMux I__8080 (
            .O(N__38018),
            .I(\pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ));
    InMux I__8079 (
            .O(N__38015),
            .I(N__38012));
    LocalMux I__8078 (
            .O(N__38012),
            .I(\pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ));
    InMux I__8077 (
            .O(N__38009),
            .I(N__38006));
    LocalMux I__8076 (
            .O(N__38006),
            .I(N__38003));
    Sp12to4 I__8075 (
            .O(N__38003),
            .I(N__38000));
    Span12Mux_s6_v I__8074 (
            .O(N__38000),
            .I(N__37997));
    Odrv12 I__8073 (
            .O(N__37997),
            .I(\pwm_generator_inst.O_14 ));
    InMux I__8072 (
            .O(N__37994),
            .I(\pwm_generator_inst.un3_threshold_cry_2 ));
    InMux I__8071 (
            .O(N__37991),
            .I(N__37988));
    LocalMux I__8070 (
            .O(N__37988),
            .I(\pwm_generator_inst.un3_threshold_axbZ0Z_4 ));
    CascadeMux I__8069 (
            .O(N__37985),
            .I(N__37982));
    InMux I__8068 (
            .O(N__37982),
            .I(N__37979));
    LocalMux I__8067 (
            .O(N__37979),
            .I(N__37975));
    InMux I__8066 (
            .O(N__37978),
            .I(N__37972));
    Odrv4 I__8065 (
            .O(N__37975),
            .I(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ));
    LocalMux I__8064 (
            .O(N__37972),
            .I(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ));
    InMux I__8063 (
            .O(N__37967),
            .I(\pwm_generator_inst.un3_threshold_cry_3 ));
    CascadeMux I__8062 (
            .O(N__37964),
            .I(N__37961));
    InMux I__8061 (
            .O(N__37961),
            .I(N__37958));
    LocalMux I__8060 (
            .O(N__37958),
            .I(N__37955));
    Odrv4 I__8059 (
            .O(N__37955),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ));
    InMux I__8058 (
            .O(N__37952),
            .I(N__37949));
    LocalMux I__8057 (
            .O(N__37949),
            .I(N__37945));
    InMux I__8056 (
            .O(N__37948),
            .I(N__37942));
    Odrv4 I__8055 (
            .O(N__37945),
            .I(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ));
    LocalMux I__8054 (
            .O(N__37942),
            .I(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ));
    InMux I__8053 (
            .O(N__37937),
            .I(\pwm_generator_inst.un3_threshold_cry_4 ));
    InMux I__8052 (
            .O(N__37934),
            .I(N__37931));
    LocalMux I__8051 (
            .O(N__37931),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ));
    InMux I__8050 (
            .O(N__37928),
            .I(N__37924));
    InMux I__8049 (
            .O(N__37927),
            .I(N__37921));
    LocalMux I__8048 (
            .O(N__37924),
            .I(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ));
    LocalMux I__8047 (
            .O(N__37921),
            .I(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ));
    InMux I__8046 (
            .O(N__37916),
            .I(\pwm_generator_inst.un3_threshold_cry_5 ));
    InMux I__8045 (
            .O(N__37913),
            .I(N__37910));
    LocalMux I__8044 (
            .O(N__37910),
            .I(N__37895));
    InMux I__8043 (
            .O(N__37909),
            .I(N__37892));
    CascadeMux I__8042 (
            .O(N__37908),
            .I(N__37875));
    CascadeMux I__8041 (
            .O(N__37907),
            .I(N__37871));
    CascadeMux I__8040 (
            .O(N__37906),
            .I(N__37867));
    CascadeMux I__8039 (
            .O(N__37905),
            .I(N__37862));
    CascadeMux I__8038 (
            .O(N__37904),
            .I(N__37858));
    CascadeMux I__8037 (
            .O(N__37903),
            .I(N__37854));
    CascadeMux I__8036 (
            .O(N__37902),
            .I(N__37850));
    CascadeMux I__8035 (
            .O(N__37901),
            .I(N__37847));
    CascadeMux I__8034 (
            .O(N__37900),
            .I(N__37843));
    CascadeMux I__8033 (
            .O(N__37899),
            .I(N__37839));
    CascadeMux I__8032 (
            .O(N__37898),
            .I(N__37835));
    Span4Mux_s2_v I__8031 (
            .O(N__37895),
            .I(N__37826));
    LocalMux I__8030 (
            .O(N__37892),
            .I(N__37826));
    InMux I__8029 (
            .O(N__37891),
            .I(N__37819));
    InMux I__8028 (
            .O(N__37890),
            .I(N__37819));
    InMux I__8027 (
            .O(N__37889),
            .I(N__37819));
    InMux I__8026 (
            .O(N__37888),
            .I(N__37810));
    InMux I__8025 (
            .O(N__37887),
            .I(N__37810));
    InMux I__8024 (
            .O(N__37886),
            .I(N__37810));
    InMux I__8023 (
            .O(N__37885),
            .I(N__37810));
    InMux I__8022 (
            .O(N__37884),
            .I(N__37807));
    InMux I__8021 (
            .O(N__37883),
            .I(N__37802));
    InMux I__8020 (
            .O(N__37882),
            .I(N__37802));
    InMux I__8019 (
            .O(N__37881),
            .I(N__37799));
    InMux I__8018 (
            .O(N__37880),
            .I(N__37779));
    InMux I__8017 (
            .O(N__37879),
            .I(N__37779));
    InMux I__8016 (
            .O(N__37878),
            .I(N__37764));
    InMux I__8015 (
            .O(N__37875),
            .I(N__37764));
    InMux I__8014 (
            .O(N__37874),
            .I(N__37764));
    InMux I__8013 (
            .O(N__37871),
            .I(N__37764));
    InMux I__8012 (
            .O(N__37870),
            .I(N__37764));
    InMux I__8011 (
            .O(N__37867),
            .I(N__37764));
    InMux I__8010 (
            .O(N__37866),
            .I(N__37764));
    InMux I__8009 (
            .O(N__37865),
            .I(N__37747));
    InMux I__8008 (
            .O(N__37862),
            .I(N__37747));
    InMux I__8007 (
            .O(N__37861),
            .I(N__37747));
    InMux I__8006 (
            .O(N__37858),
            .I(N__37747));
    InMux I__8005 (
            .O(N__37857),
            .I(N__37747));
    InMux I__8004 (
            .O(N__37854),
            .I(N__37747));
    InMux I__8003 (
            .O(N__37853),
            .I(N__37747));
    InMux I__8002 (
            .O(N__37850),
            .I(N__37747));
    InMux I__8001 (
            .O(N__37847),
            .I(N__37730));
    InMux I__8000 (
            .O(N__37846),
            .I(N__37730));
    InMux I__7999 (
            .O(N__37843),
            .I(N__37730));
    InMux I__7998 (
            .O(N__37842),
            .I(N__37730));
    InMux I__7997 (
            .O(N__37839),
            .I(N__37730));
    InMux I__7996 (
            .O(N__37838),
            .I(N__37730));
    InMux I__7995 (
            .O(N__37835),
            .I(N__37730));
    InMux I__7994 (
            .O(N__37834),
            .I(N__37730));
    CascadeMux I__7993 (
            .O(N__37833),
            .I(N__37726));
    CascadeMux I__7992 (
            .O(N__37832),
            .I(N__37722));
    CascadeMux I__7991 (
            .O(N__37831),
            .I(N__37718));
    Span4Mux_v I__7990 (
            .O(N__37826),
            .I(N__37709));
    LocalMux I__7989 (
            .O(N__37819),
            .I(N__37709));
    LocalMux I__7988 (
            .O(N__37810),
            .I(N__37709));
    LocalMux I__7987 (
            .O(N__37807),
            .I(N__37702));
    LocalMux I__7986 (
            .O(N__37802),
            .I(N__37702));
    LocalMux I__7985 (
            .O(N__37799),
            .I(N__37702));
    InMux I__7984 (
            .O(N__37798),
            .I(N__37699));
    InMux I__7983 (
            .O(N__37797),
            .I(N__37694));
    InMux I__7982 (
            .O(N__37796),
            .I(N__37694));
    InMux I__7981 (
            .O(N__37795),
            .I(N__37691));
    InMux I__7980 (
            .O(N__37794),
            .I(N__37688));
    InMux I__7979 (
            .O(N__37793),
            .I(N__37685));
    InMux I__7978 (
            .O(N__37792),
            .I(N__37682));
    InMux I__7977 (
            .O(N__37791),
            .I(N__37679));
    InMux I__7976 (
            .O(N__37790),
            .I(N__37672));
    InMux I__7975 (
            .O(N__37789),
            .I(N__37672));
    InMux I__7974 (
            .O(N__37788),
            .I(N__37672));
    InMux I__7973 (
            .O(N__37787),
            .I(N__37663));
    InMux I__7972 (
            .O(N__37786),
            .I(N__37663));
    InMux I__7971 (
            .O(N__37785),
            .I(N__37663));
    InMux I__7970 (
            .O(N__37784),
            .I(N__37663));
    LocalMux I__7969 (
            .O(N__37779),
            .I(N__37660));
    LocalMux I__7968 (
            .O(N__37764),
            .I(N__37655));
    LocalMux I__7967 (
            .O(N__37747),
            .I(N__37655));
    LocalMux I__7966 (
            .O(N__37730),
            .I(N__37652));
    InMux I__7965 (
            .O(N__37729),
            .I(N__37637));
    InMux I__7964 (
            .O(N__37726),
            .I(N__37637));
    InMux I__7963 (
            .O(N__37725),
            .I(N__37637));
    InMux I__7962 (
            .O(N__37722),
            .I(N__37637));
    InMux I__7961 (
            .O(N__37721),
            .I(N__37637));
    InMux I__7960 (
            .O(N__37718),
            .I(N__37637));
    InMux I__7959 (
            .O(N__37717),
            .I(N__37637));
    CascadeMux I__7958 (
            .O(N__37716),
            .I(N__37633));
    Span4Mux_v I__7957 (
            .O(N__37709),
            .I(N__37629));
    Span12Mux_s7_v I__7956 (
            .O(N__37702),
            .I(N__37620));
    LocalMux I__7955 (
            .O(N__37699),
            .I(N__37620));
    LocalMux I__7954 (
            .O(N__37694),
            .I(N__37620));
    LocalMux I__7953 (
            .O(N__37691),
            .I(N__37620));
    LocalMux I__7952 (
            .O(N__37688),
            .I(N__37607));
    LocalMux I__7951 (
            .O(N__37685),
            .I(N__37607));
    LocalMux I__7950 (
            .O(N__37682),
            .I(N__37607));
    LocalMux I__7949 (
            .O(N__37679),
            .I(N__37607));
    LocalMux I__7948 (
            .O(N__37672),
            .I(N__37607));
    LocalMux I__7947 (
            .O(N__37663),
            .I(N__37607));
    Span4Mux_h I__7946 (
            .O(N__37660),
            .I(N__37604));
    Span4Mux_v I__7945 (
            .O(N__37655),
            .I(N__37601));
    Span4Mux_h I__7944 (
            .O(N__37652),
            .I(N__37596));
    LocalMux I__7943 (
            .O(N__37637),
            .I(N__37596));
    InMux I__7942 (
            .O(N__37636),
            .I(N__37589));
    InMux I__7941 (
            .O(N__37633),
            .I(N__37589));
    InMux I__7940 (
            .O(N__37632),
            .I(N__37589));
    Sp12to4 I__7939 (
            .O(N__37629),
            .I(N__37586));
    Span12Mux_v I__7938 (
            .O(N__37620),
            .I(N__37581));
    Span12Mux_s10_v I__7937 (
            .O(N__37607),
            .I(N__37581));
    Span4Mux_v I__7936 (
            .O(N__37604),
            .I(N__37578));
    Span4Mux_v I__7935 (
            .O(N__37601),
            .I(N__37573));
    Span4Mux_v I__7934 (
            .O(N__37596),
            .I(N__37573));
    LocalMux I__7933 (
            .O(N__37589),
            .I(N__37570));
    Span12Mux_h I__7932 (
            .O(N__37586),
            .I(N__37565));
    Span12Mux_h I__7931 (
            .O(N__37581),
            .I(N__37565));
    Span4Mux_v I__7930 (
            .O(N__37578),
            .I(N__37562));
    Span4Mux_v I__7929 (
            .O(N__37573),
            .I(N__37559));
    Span4Mux_v I__7928 (
            .O(N__37570),
            .I(N__37556));
    Odrv12 I__7927 (
            .O(N__37565),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__7926 (
            .O(N__37562),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__7925 (
            .O(N__37559),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__7924 (
            .O(N__37556),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__7923 (
            .O(N__37547),
            .I(N__37544));
    InMux I__7922 (
            .O(N__37544),
            .I(N__37541));
    LocalMux I__7921 (
            .O(N__37541),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ));
    InMux I__7920 (
            .O(N__37538),
            .I(N__37535));
    LocalMux I__7919 (
            .O(N__37535),
            .I(N__37531));
    InMux I__7918 (
            .O(N__37534),
            .I(N__37528));
    Odrv4 I__7917 (
            .O(N__37531),
            .I(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ));
    LocalMux I__7916 (
            .O(N__37528),
            .I(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ));
    InMux I__7915 (
            .O(N__37523),
            .I(\pwm_generator_inst.un3_threshold_cry_6 ));
    InMux I__7914 (
            .O(N__37520),
            .I(N__37517));
    LocalMux I__7913 (
            .O(N__37517),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ));
    InMux I__7912 (
            .O(N__37514),
            .I(N__37511));
    LocalMux I__7911 (
            .O(N__37511),
            .I(N__37508));
    Span4Mux_v I__7910 (
            .O(N__37508),
            .I(N__37505));
    Odrv4 I__7909 (
            .O(N__37505),
            .I(\pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ));
    InMux I__7908 (
            .O(N__37502),
            .I(bfn_14_29_0_));
    InMux I__7907 (
            .O(N__37499),
            .I(N__37496));
    LocalMux I__7906 (
            .O(N__37496),
            .I(\pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ));
    InMux I__7905 (
            .O(N__37493),
            .I(N__37490));
    LocalMux I__7904 (
            .O(N__37490),
            .I(\pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ));
    InMux I__7903 (
            .O(N__37487),
            .I(\pwm_generator_inst.un15_threshold_1_cry_17 ));
    InMux I__7902 (
            .O(N__37484),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18 ));
    InMux I__7901 (
            .O(N__37481),
            .I(N__37478));
    LocalMux I__7900 (
            .O(N__37478),
            .I(N__37475));
    Odrv4 I__7899 (
            .O(N__37475),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ));
    CascadeMux I__7898 (
            .O(N__37472),
            .I(N__37469));
    InMux I__7897 (
            .O(N__37469),
            .I(N__37464));
    InMux I__7896 (
            .O(N__37468),
            .I(N__37459));
    InMux I__7895 (
            .O(N__37467),
            .I(N__37459));
    LocalMux I__7894 (
            .O(N__37464),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    LocalMux I__7893 (
            .O(N__37459),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    InMux I__7892 (
            .O(N__37454),
            .I(N__37449));
    InMux I__7891 (
            .O(N__37453),
            .I(N__37444));
    InMux I__7890 (
            .O(N__37452),
            .I(N__37444));
    LocalMux I__7889 (
            .O(N__37449),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    LocalMux I__7888 (
            .O(N__37444),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    InMux I__7887 (
            .O(N__37439),
            .I(N__37435));
    InMux I__7886 (
            .O(N__37438),
            .I(N__37431));
    LocalMux I__7885 (
            .O(N__37435),
            .I(N__37428));
    InMux I__7884 (
            .O(N__37434),
            .I(N__37425));
    LocalMux I__7883 (
            .O(N__37431),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    Odrv4 I__7882 (
            .O(N__37428),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    LocalMux I__7881 (
            .O(N__37425),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    CascadeMux I__7880 (
            .O(N__37418),
            .I(N__37414));
    InMux I__7879 (
            .O(N__37417),
            .I(N__37410));
    InMux I__7878 (
            .O(N__37414),
            .I(N__37407));
    InMux I__7877 (
            .O(N__37413),
            .I(N__37404));
    LocalMux I__7876 (
            .O(N__37410),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    LocalMux I__7875 (
            .O(N__37407),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    LocalMux I__7874 (
            .O(N__37404),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    InMux I__7873 (
            .O(N__37397),
            .I(N__37394));
    LocalMux I__7872 (
            .O(N__37394),
            .I(N__37390));
    InMux I__7871 (
            .O(N__37393),
            .I(N__37387));
    Span4Mux_v I__7870 (
            .O(N__37390),
            .I(N__37382));
    LocalMux I__7869 (
            .O(N__37387),
            .I(N__37382));
    Span4Mux_h I__7868 (
            .O(N__37382),
            .I(N__37379));
    Span4Mux_h I__7867 (
            .O(N__37379),
            .I(N__37376));
    Span4Mux_v I__7866 (
            .O(N__37376),
            .I(N__37373));
    Odrv4 I__7865 (
            .O(N__37373),
            .I(\pwm_generator_inst.un3_threshold ));
    InMux I__7864 (
            .O(N__37370),
            .I(N__37367));
    LocalMux I__7863 (
            .O(N__37367),
            .I(N__37364));
    Span12Mux_h I__7862 (
            .O(N__37364),
            .I(N__37361));
    Odrv12 I__7861 (
            .O(N__37361),
            .I(\pwm_generator_inst.O_12 ));
    InMux I__7860 (
            .O(N__37358),
            .I(N__37355));
    LocalMux I__7859 (
            .O(N__37355),
            .I(N__37351));
    InMux I__7858 (
            .O(N__37354),
            .I(N__37348));
    Odrv4 I__7857 (
            .O(N__37351),
            .I(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ));
    LocalMux I__7856 (
            .O(N__37348),
            .I(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ));
    InMux I__7855 (
            .O(N__37343),
            .I(\pwm_generator_inst.un3_threshold_cry_0 ));
    InMux I__7854 (
            .O(N__37340),
            .I(N__37337));
    LocalMux I__7853 (
            .O(N__37337),
            .I(N__37334));
    Span4Mux_v I__7852 (
            .O(N__37334),
            .I(N__37331));
    Span4Mux_h I__7851 (
            .O(N__37331),
            .I(N__37328));
    Span4Mux_h I__7850 (
            .O(N__37328),
            .I(N__37325));
    Odrv4 I__7849 (
            .O(N__37325),
            .I(\pwm_generator_inst.O_13 ));
    InMux I__7848 (
            .O(N__37322),
            .I(\pwm_generator_inst.un3_threshold_cry_1 ));
    InMux I__7847 (
            .O(N__37319),
            .I(N__37316));
    LocalMux I__7846 (
            .O(N__37316),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ));
    InMux I__7845 (
            .O(N__37313),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9 ));
    CascadeMux I__7844 (
            .O(N__37310),
            .I(N__37302));
    CascadeMux I__7843 (
            .O(N__37309),
            .I(N__37299));
    CascadeMux I__7842 (
            .O(N__37308),
            .I(N__37292));
    CascadeMux I__7841 (
            .O(N__37307),
            .I(N__37289));
    CascadeMux I__7840 (
            .O(N__37306),
            .I(N__37285));
    InMux I__7839 (
            .O(N__37305),
            .I(N__37281));
    InMux I__7838 (
            .O(N__37302),
            .I(N__37278));
    InMux I__7837 (
            .O(N__37299),
            .I(N__37273));
    InMux I__7836 (
            .O(N__37298),
            .I(N__37273));
    InMux I__7835 (
            .O(N__37297),
            .I(N__37268));
    InMux I__7834 (
            .O(N__37296),
            .I(N__37268));
    InMux I__7833 (
            .O(N__37295),
            .I(N__37265));
    InMux I__7832 (
            .O(N__37292),
            .I(N__37262));
    InMux I__7831 (
            .O(N__37289),
            .I(N__37253));
    InMux I__7830 (
            .O(N__37288),
            .I(N__37253));
    InMux I__7829 (
            .O(N__37285),
            .I(N__37253));
    InMux I__7828 (
            .O(N__37284),
            .I(N__37253));
    LocalMux I__7827 (
            .O(N__37281),
            .I(N__37246));
    LocalMux I__7826 (
            .O(N__37278),
            .I(N__37246));
    LocalMux I__7825 (
            .O(N__37273),
            .I(N__37246));
    LocalMux I__7824 (
            .O(N__37268),
            .I(N__37241));
    LocalMux I__7823 (
            .O(N__37265),
            .I(N__37241));
    LocalMux I__7822 (
            .O(N__37262),
            .I(N__37238));
    LocalMux I__7821 (
            .O(N__37253),
            .I(N__37235));
    Span4Mux_v I__7820 (
            .O(N__37246),
            .I(N__37230));
    Span4Mux_h I__7819 (
            .O(N__37241),
            .I(N__37230));
    Odrv12 I__7818 (
            .O(N__37238),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    Odrv12 I__7817 (
            .O(N__37235),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    Odrv4 I__7816 (
            .O(N__37230),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    InMux I__7815 (
            .O(N__37223),
            .I(N__37220));
    LocalMux I__7814 (
            .O(N__37220),
            .I(N__37217));
    Odrv4 I__7813 (
            .O(N__37217),
            .I(\pwm_generator_inst.un19_threshold_axb_1 ));
    InMux I__7812 (
            .O(N__37214),
            .I(\pwm_generator_inst.un15_threshold_1_cry_10 ));
    InMux I__7811 (
            .O(N__37211),
            .I(N__37208));
    LocalMux I__7810 (
            .O(N__37208),
            .I(\pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ));
    InMux I__7809 (
            .O(N__37205),
            .I(\pwm_generator_inst.un15_threshold_1_cry_11 ));
    InMux I__7808 (
            .O(N__37202),
            .I(N__37199));
    LocalMux I__7807 (
            .O(N__37199),
            .I(\pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ));
    InMux I__7806 (
            .O(N__37196),
            .I(\pwm_generator_inst.un15_threshold_1_cry_12 ));
    InMux I__7805 (
            .O(N__37193),
            .I(N__37190));
    LocalMux I__7804 (
            .O(N__37190),
            .I(\pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ));
    InMux I__7803 (
            .O(N__37187),
            .I(\pwm_generator_inst.un15_threshold_1_cry_13 ));
    InMux I__7802 (
            .O(N__37184),
            .I(N__37181));
    LocalMux I__7801 (
            .O(N__37181),
            .I(\pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ));
    InMux I__7800 (
            .O(N__37178),
            .I(\pwm_generator_inst.un15_threshold_1_cry_14 ));
    InMux I__7799 (
            .O(N__37175),
            .I(N__37171));
    InMux I__7798 (
            .O(N__37174),
            .I(N__37167));
    LocalMux I__7797 (
            .O(N__37171),
            .I(N__37164));
    InMux I__7796 (
            .O(N__37170),
            .I(N__37161));
    LocalMux I__7795 (
            .O(N__37167),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    Odrv4 I__7794 (
            .O(N__37164),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    LocalMux I__7793 (
            .O(N__37161),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    InMux I__7792 (
            .O(N__37154),
            .I(N__37151));
    LocalMux I__7791 (
            .O(N__37151),
            .I(N__37148));
    Odrv4 I__7790 (
            .O(N__37148),
            .I(\pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ));
    InMux I__7789 (
            .O(N__37145),
            .I(bfn_14_27_0_));
    InMux I__7788 (
            .O(N__37142),
            .I(N__37139));
    LocalMux I__7787 (
            .O(N__37139),
            .I(\pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ));
    InMux I__7786 (
            .O(N__37136),
            .I(\pwm_generator_inst.un15_threshold_1_cry_16 ));
    InMux I__7785 (
            .O(N__37133),
            .I(N__37130));
    LocalMux I__7784 (
            .O(N__37130),
            .I(\pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ));
    InMux I__7783 (
            .O(N__37127),
            .I(N__37124));
    LocalMux I__7782 (
            .O(N__37124),
            .I(\pwm_generator_inst.un15_threshold_1_axb_2 ));
    InMux I__7781 (
            .O(N__37121),
            .I(N__37118));
    LocalMux I__7780 (
            .O(N__37118),
            .I(N__37115));
    Span4Mux_v I__7779 (
            .O(N__37115),
            .I(N__37112));
    Span4Mux_h I__7778 (
            .O(N__37112),
            .I(N__37109));
    Span4Mux_h I__7777 (
            .O(N__37109),
            .I(N__37106));
    Odrv4 I__7776 (
            .O(N__37106),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__7775 (
            .O(N__37103),
            .I(N__37100));
    LocalMux I__7774 (
            .O(N__37100),
            .I(\pwm_generator_inst.un15_threshold_1_axb_3 ));
    InMux I__7773 (
            .O(N__37097),
            .I(N__37094));
    LocalMux I__7772 (
            .O(N__37094),
            .I(N__37091));
    Span4Mux_v I__7771 (
            .O(N__37091),
            .I(N__37088));
    Span4Mux_h I__7770 (
            .O(N__37088),
            .I(N__37085));
    Span4Mux_h I__7769 (
            .O(N__37085),
            .I(N__37082));
    Odrv4 I__7768 (
            .O(N__37082),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__7767 (
            .O(N__37079),
            .I(N__37076));
    LocalMux I__7766 (
            .O(N__37076),
            .I(\pwm_generator_inst.un15_threshold_1_axb_4 ));
    InMux I__7765 (
            .O(N__37073),
            .I(N__37070));
    LocalMux I__7764 (
            .O(N__37070),
            .I(N__37067));
    Span4Mux_h I__7763 (
            .O(N__37067),
            .I(N__37064));
    Span4Mux_h I__7762 (
            .O(N__37064),
            .I(N__37061));
    Span4Mux_h I__7761 (
            .O(N__37061),
            .I(N__37058));
    Odrv4 I__7760 (
            .O(N__37058),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__7759 (
            .O(N__37055),
            .I(N__37052));
    LocalMux I__7758 (
            .O(N__37052),
            .I(\pwm_generator_inst.un15_threshold_1_axb_5 ));
    InMux I__7757 (
            .O(N__37049),
            .I(N__37046));
    LocalMux I__7756 (
            .O(N__37046),
            .I(N__37043));
    Span4Mux_h I__7755 (
            .O(N__37043),
            .I(N__37040));
    Span4Mux_h I__7754 (
            .O(N__37040),
            .I(N__37037));
    Span4Mux_h I__7753 (
            .O(N__37037),
            .I(N__37034));
    Odrv4 I__7752 (
            .O(N__37034),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__7751 (
            .O(N__37031),
            .I(N__37028));
    LocalMux I__7750 (
            .O(N__37028),
            .I(\pwm_generator_inst.un15_threshold_1_axb_6 ));
    InMux I__7749 (
            .O(N__37025),
            .I(N__37022));
    LocalMux I__7748 (
            .O(N__37022),
            .I(N__37019));
    Span12Mux_s7_v I__7747 (
            .O(N__37019),
            .I(N__37016));
    Odrv12 I__7746 (
            .O(N__37016),
            .I(\pwm_generator_inst.O_7 ));
    InMux I__7745 (
            .O(N__37013),
            .I(N__37010));
    LocalMux I__7744 (
            .O(N__37010),
            .I(\pwm_generator_inst.un15_threshold_1_axb_7 ));
    InMux I__7743 (
            .O(N__37007),
            .I(N__37004));
    LocalMux I__7742 (
            .O(N__37004),
            .I(N__37001));
    Span4Mux_v I__7741 (
            .O(N__37001),
            .I(N__36998));
    Span4Mux_h I__7740 (
            .O(N__36998),
            .I(N__36995));
    Span4Mux_h I__7739 (
            .O(N__36995),
            .I(N__36992));
    Odrv4 I__7738 (
            .O(N__36992),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__7737 (
            .O(N__36989),
            .I(N__36986));
    LocalMux I__7736 (
            .O(N__36986),
            .I(\pwm_generator_inst.un15_threshold_1_axb_8 ));
    InMux I__7735 (
            .O(N__36983),
            .I(N__36980));
    LocalMux I__7734 (
            .O(N__36980),
            .I(N__36977));
    Span4Mux_h I__7733 (
            .O(N__36977),
            .I(N__36974));
    Span4Mux_h I__7732 (
            .O(N__36974),
            .I(N__36971));
    Span4Mux_h I__7731 (
            .O(N__36971),
            .I(N__36968));
    Odrv4 I__7730 (
            .O(N__36968),
            .I(\pwm_generator_inst.O_9 ));
    InMux I__7729 (
            .O(N__36965),
            .I(N__36962));
    LocalMux I__7728 (
            .O(N__36962),
            .I(\pwm_generator_inst.un15_threshold_1_axb_9 ));
    CascadeMux I__7727 (
            .O(N__36959),
            .I(N__36955));
    InMux I__7726 (
            .O(N__36958),
            .I(N__36951));
    InMux I__7725 (
            .O(N__36955),
            .I(N__36948));
    InMux I__7724 (
            .O(N__36954),
            .I(N__36945));
    LocalMux I__7723 (
            .O(N__36951),
            .I(N__36938));
    LocalMux I__7722 (
            .O(N__36948),
            .I(N__36938));
    LocalMux I__7721 (
            .O(N__36945),
            .I(N__36938));
    Odrv4 I__7720 (
            .O(N__36938),
            .I(il_max_comp1_D2));
    InMux I__7719 (
            .O(N__36935),
            .I(N__36932));
    LocalMux I__7718 (
            .O(N__36932),
            .I(N__36928));
    InMux I__7717 (
            .O(N__36931),
            .I(N__36925));
    Span4Mux_h I__7716 (
            .O(N__36928),
            .I(N__36922));
    LocalMux I__7715 (
            .O(N__36925),
            .I(N__36919));
    Span4Mux_h I__7714 (
            .O(N__36922),
            .I(N__36916));
    Span4Mux_s3_h I__7713 (
            .O(N__36919),
            .I(N__36913));
    Span4Mux_v I__7712 (
            .O(N__36916),
            .I(N__36908));
    Span4Mux_h I__7711 (
            .O(N__36913),
            .I(N__36908));
    Odrv4 I__7710 (
            .O(N__36908),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    InMux I__7709 (
            .O(N__36905),
            .I(N__36902));
    LocalMux I__7708 (
            .O(N__36902),
            .I(N__36898));
    InMux I__7707 (
            .O(N__36901),
            .I(N__36895));
    Span4Mux_h I__7706 (
            .O(N__36898),
            .I(N__36892));
    LocalMux I__7705 (
            .O(N__36895),
            .I(N__36889));
    Span4Mux_v I__7704 (
            .O(N__36892),
            .I(N__36886));
    Span4Mux_s3_h I__7703 (
            .O(N__36889),
            .I(N__36883));
    Span4Mux_v I__7702 (
            .O(N__36886),
            .I(N__36880));
    Span4Mux_h I__7701 (
            .O(N__36883),
            .I(N__36877));
    Odrv4 I__7700 (
            .O(N__36880),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    Odrv4 I__7699 (
            .O(N__36877),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    CascadeMux I__7698 (
            .O(N__36872),
            .I(N__36869));
    InMux I__7697 (
            .O(N__36869),
            .I(N__36861));
    InMux I__7696 (
            .O(N__36868),
            .I(N__36861));
    InMux I__7695 (
            .O(N__36867),
            .I(N__36858));
    InMux I__7694 (
            .O(N__36866),
            .I(N__36855));
    LocalMux I__7693 (
            .O(N__36861),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__7692 (
            .O(N__36858),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__7691 (
            .O(N__36855),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    InMux I__7690 (
            .O(N__36848),
            .I(N__36842));
    InMux I__7689 (
            .O(N__36847),
            .I(N__36835));
    InMux I__7688 (
            .O(N__36846),
            .I(N__36835));
    InMux I__7687 (
            .O(N__36845),
            .I(N__36835));
    LocalMux I__7686 (
            .O(N__36842),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__7685 (
            .O(N__36835),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    InMux I__7684 (
            .O(N__36830),
            .I(N__36826));
    InMux I__7683 (
            .O(N__36829),
            .I(N__36823));
    LocalMux I__7682 (
            .O(N__36826),
            .I(N__36820));
    LocalMux I__7681 (
            .O(N__36823),
            .I(N__36817));
    Span4Mux_h I__7680 (
            .O(N__36820),
            .I(N__36814));
    Span12Mux_v I__7679 (
            .O(N__36817),
            .I(N__36811));
    Span4Mux_h I__7678 (
            .O(N__36814),
            .I(N__36808));
    Odrv12 I__7677 (
            .O(N__36811),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    Odrv4 I__7676 (
            .O(N__36808),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    InMux I__7675 (
            .O(N__36803),
            .I(N__36800));
    LocalMux I__7674 (
            .O(N__36800),
            .I(N__36797));
    Span4Mux_h I__7673 (
            .O(N__36797),
            .I(N__36794));
    Span4Mux_h I__7672 (
            .O(N__36794),
            .I(N__36791));
    Span4Mux_h I__7671 (
            .O(N__36791),
            .I(N__36788));
    Odrv4 I__7670 (
            .O(N__36788),
            .I(\pwm_generator_inst.O_0 ));
    InMux I__7669 (
            .O(N__36785),
            .I(N__36782));
    LocalMux I__7668 (
            .O(N__36782),
            .I(\pwm_generator_inst.un15_threshold_1_axb_0 ));
    InMux I__7667 (
            .O(N__36779),
            .I(N__36776));
    LocalMux I__7666 (
            .O(N__36776),
            .I(N__36773));
    Span4Mux_h I__7665 (
            .O(N__36773),
            .I(N__36770));
    Span4Mux_h I__7664 (
            .O(N__36770),
            .I(N__36767));
    Span4Mux_h I__7663 (
            .O(N__36767),
            .I(N__36764));
    Odrv4 I__7662 (
            .O(N__36764),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__7661 (
            .O(N__36761),
            .I(N__36758));
    LocalMux I__7660 (
            .O(N__36758),
            .I(\pwm_generator_inst.un15_threshold_1_axb_1 ));
    InMux I__7659 (
            .O(N__36755),
            .I(N__36752));
    LocalMux I__7658 (
            .O(N__36752),
            .I(N__36749));
    Span12Mux_h I__7657 (
            .O(N__36749),
            .I(N__36746));
    Odrv12 I__7656 (
            .O(N__36746),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__7655 (
            .O(N__36743),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    InMux I__7654 (
            .O(N__36740),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    InMux I__7653 (
            .O(N__36737),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__7652 (
            .O(N__36734),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__7651 (
            .O(N__36731),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    InMux I__7650 (
            .O(N__36728),
            .I(N__36690));
    InMux I__7649 (
            .O(N__36727),
            .I(N__36690));
    InMux I__7648 (
            .O(N__36726),
            .I(N__36690));
    InMux I__7647 (
            .O(N__36725),
            .I(N__36690));
    InMux I__7646 (
            .O(N__36724),
            .I(N__36681));
    InMux I__7645 (
            .O(N__36723),
            .I(N__36681));
    InMux I__7644 (
            .O(N__36722),
            .I(N__36681));
    InMux I__7643 (
            .O(N__36721),
            .I(N__36681));
    InMux I__7642 (
            .O(N__36720),
            .I(N__36672));
    InMux I__7641 (
            .O(N__36719),
            .I(N__36672));
    InMux I__7640 (
            .O(N__36718),
            .I(N__36672));
    InMux I__7639 (
            .O(N__36717),
            .I(N__36672));
    InMux I__7638 (
            .O(N__36716),
            .I(N__36663));
    InMux I__7637 (
            .O(N__36715),
            .I(N__36663));
    InMux I__7636 (
            .O(N__36714),
            .I(N__36663));
    InMux I__7635 (
            .O(N__36713),
            .I(N__36663));
    InMux I__7634 (
            .O(N__36712),
            .I(N__36654));
    InMux I__7633 (
            .O(N__36711),
            .I(N__36654));
    InMux I__7632 (
            .O(N__36710),
            .I(N__36654));
    InMux I__7631 (
            .O(N__36709),
            .I(N__36654));
    InMux I__7630 (
            .O(N__36708),
            .I(N__36649));
    InMux I__7629 (
            .O(N__36707),
            .I(N__36649));
    InMux I__7628 (
            .O(N__36706),
            .I(N__36640));
    InMux I__7627 (
            .O(N__36705),
            .I(N__36640));
    InMux I__7626 (
            .O(N__36704),
            .I(N__36640));
    InMux I__7625 (
            .O(N__36703),
            .I(N__36640));
    InMux I__7624 (
            .O(N__36702),
            .I(N__36631));
    InMux I__7623 (
            .O(N__36701),
            .I(N__36631));
    InMux I__7622 (
            .O(N__36700),
            .I(N__36631));
    InMux I__7621 (
            .O(N__36699),
            .I(N__36631));
    LocalMux I__7620 (
            .O(N__36690),
            .I(N__36626));
    LocalMux I__7619 (
            .O(N__36681),
            .I(N__36626));
    LocalMux I__7618 (
            .O(N__36672),
            .I(N__36619));
    LocalMux I__7617 (
            .O(N__36663),
            .I(N__36619));
    LocalMux I__7616 (
            .O(N__36654),
            .I(N__36619));
    LocalMux I__7615 (
            .O(N__36649),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    LocalMux I__7614 (
            .O(N__36640),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    LocalMux I__7613 (
            .O(N__36631),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__7612 (
            .O(N__36626),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv12 I__7611 (
            .O(N__36619),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    CEMux I__7610 (
            .O(N__36608),
            .I(N__36602));
    CEMux I__7609 (
            .O(N__36607),
            .I(N__36598));
    CEMux I__7608 (
            .O(N__36606),
            .I(N__36590));
    CEMux I__7607 (
            .O(N__36605),
            .I(N__36587));
    LocalMux I__7606 (
            .O(N__36602),
            .I(N__36584));
    CEMux I__7605 (
            .O(N__36601),
            .I(N__36581));
    LocalMux I__7604 (
            .O(N__36598),
            .I(N__36555));
    CEMux I__7603 (
            .O(N__36597),
            .I(N__36552));
    CEMux I__7602 (
            .O(N__36596),
            .I(N__36549));
    CEMux I__7601 (
            .O(N__36595),
            .I(N__36539));
    CEMux I__7600 (
            .O(N__36594),
            .I(N__36535));
    CEMux I__7599 (
            .O(N__36593),
            .I(N__36532));
    LocalMux I__7598 (
            .O(N__36590),
            .I(N__36522));
    LocalMux I__7597 (
            .O(N__36587),
            .I(N__36522));
    Span4Mux_v I__7596 (
            .O(N__36584),
            .I(N__36522));
    LocalMux I__7595 (
            .O(N__36581),
            .I(N__36522));
    InMux I__7594 (
            .O(N__36580),
            .I(N__36513));
    InMux I__7593 (
            .O(N__36579),
            .I(N__36513));
    InMux I__7592 (
            .O(N__36578),
            .I(N__36513));
    InMux I__7591 (
            .O(N__36577),
            .I(N__36513));
    InMux I__7590 (
            .O(N__36576),
            .I(N__36506));
    InMux I__7589 (
            .O(N__36575),
            .I(N__36506));
    InMux I__7588 (
            .O(N__36574),
            .I(N__36506));
    InMux I__7587 (
            .O(N__36573),
            .I(N__36497));
    InMux I__7586 (
            .O(N__36572),
            .I(N__36497));
    InMux I__7585 (
            .O(N__36571),
            .I(N__36497));
    InMux I__7584 (
            .O(N__36570),
            .I(N__36497));
    InMux I__7583 (
            .O(N__36569),
            .I(N__36488));
    InMux I__7582 (
            .O(N__36568),
            .I(N__36488));
    InMux I__7581 (
            .O(N__36567),
            .I(N__36488));
    InMux I__7580 (
            .O(N__36566),
            .I(N__36488));
    InMux I__7579 (
            .O(N__36565),
            .I(N__36479));
    InMux I__7578 (
            .O(N__36564),
            .I(N__36479));
    InMux I__7577 (
            .O(N__36563),
            .I(N__36479));
    InMux I__7576 (
            .O(N__36562),
            .I(N__36479));
    InMux I__7575 (
            .O(N__36561),
            .I(N__36470));
    InMux I__7574 (
            .O(N__36560),
            .I(N__36470));
    InMux I__7573 (
            .O(N__36559),
            .I(N__36470));
    InMux I__7572 (
            .O(N__36558),
            .I(N__36470));
    Span4Mux_v I__7571 (
            .O(N__36555),
            .I(N__36464));
    LocalMux I__7570 (
            .O(N__36552),
            .I(N__36464));
    LocalMux I__7569 (
            .O(N__36549),
            .I(N__36461));
    InMux I__7568 (
            .O(N__36548),
            .I(N__36454));
    InMux I__7567 (
            .O(N__36547),
            .I(N__36454));
    InMux I__7566 (
            .O(N__36546),
            .I(N__36454));
    InMux I__7565 (
            .O(N__36545),
            .I(N__36445));
    InMux I__7564 (
            .O(N__36544),
            .I(N__36445));
    InMux I__7563 (
            .O(N__36543),
            .I(N__36445));
    InMux I__7562 (
            .O(N__36542),
            .I(N__36445));
    LocalMux I__7561 (
            .O(N__36539),
            .I(N__36441));
    CEMux I__7560 (
            .O(N__36538),
            .I(N__36438));
    LocalMux I__7559 (
            .O(N__36535),
            .I(N__36435));
    LocalMux I__7558 (
            .O(N__36532),
            .I(N__36432));
    CEMux I__7557 (
            .O(N__36531),
            .I(N__36429));
    Span4Mux_v I__7556 (
            .O(N__36522),
            .I(N__36426));
    LocalMux I__7555 (
            .O(N__36513),
            .I(N__36417));
    LocalMux I__7554 (
            .O(N__36506),
            .I(N__36417));
    LocalMux I__7553 (
            .O(N__36497),
            .I(N__36417));
    LocalMux I__7552 (
            .O(N__36488),
            .I(N__36417));
    LocalMux I__7551 (
            .O(N__36479),
            .I(N__36412));
    LocalMux I__7550 (
            .O(N__36470),
            .I(N__36412));
    InMux I__7549 (
            .O(N__36469),
            .I(N__36409));
    Span4Mux_h I__7548 (
            .O(N__36464),
            .I(N__36404));
    Span4Mux_v I__7547 (
            .O(N__36461),
            .I(N__36404));
    LocalMux I__7546 (
            .O(N__36454),
            .I(N__36399));
    LocalMux I__7545 (
            .O(N__36445),
            .I(N__36399));
    CEMux I__7544 (
            .O(N__36444),
            .I(N__36396));
    Span4Mux_h I__7543 (
            .O(N__36441),
            .I(N__36393));
    LocalMux I__7542 (
            .O(N__36438),
            .I(N__36386));
    Span4Mux_v I__7541 (
            .O(N__36435),
            .I(N__36386));
    Span4Mux_h I__7540 (
            .O(N__36432),
            .I(N__36386));
    LocalMux I__7539 (
            .O(N__36429),
            .I(N__36383));
    Span4Mux_v I__7538 (
            .O(N__36426),
            .I(N__36380));
    Span4Mux_v I__7537 (
            .O(N__36417),
            .I(N__36375));
    Span4Mux_v I__7536 (
            .O(N__36412),
            .I(N__36375));
    LocalMux I__7535 (
            .O(N__36409),
            .I(N__36372));
    Span4Mux_h I__7534 (
            .O(N__36404),
            .I(N__36367));
    Span4Mux_h I__7533 (
            .O(N__36399),
            .I(N__36367));
    LocalMux I__7532 (
            .O(N__36396),
            .I(N__36364));
    Span4Mux_h I__7531 (
            .O(N__36393),
            .I(N__36357));
    Span4Mux_v I__7530 (
            .O(N__36386),
            .I(N__36357));
    Span4Mux_v I__7529 (
            .O(N__36383),
            .I(N__36357));
    Span4Mux_h I__7528 (
            .O(N__36380),
            .I(N__36354));
    Span4Mux_v I__7527 (
            .O(N__36375),
            .I(N__36351));
    Span4Mux_h I__7526 (
            .O(N__36372),
            .I(N__36346));
    Span4Mux_v I__7525 (
            .O(N__36367),
            .I(N__36346));
    Span12Mux_h I__7524 (
            .O(N__36364),
            .I(N__36341));
    Sp12to4 I__7523 (
            .O(N__36357),
            .I(N__36341));
    Span4Mux_h I__7522 (
            .O(N__36354),
            .I(N__36338));
    Span4Mux_v I__7521 (
            .O(N__36351),
            .I(N__36335));
    Span4Mux_v I__7520 (
            .O(N__36346),
            .I(N__36332));
    Odrv12 I__7519 (
            .O(N__36341),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__7518 (
            .O(N__36338),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__7517 (
            .O(N__36335),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__7516 (
            .O(N__36332),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    InMux I__7515 (
            .O(N__36323),
            .I(N__36320));
    LocalMux I__7514 (
            .O(N__36320),
            .I(N__36317));
    Span4Mux_v I__7513 (
            .O(N__36317),
            .I(N__36313));
    InMux I__7512 (
            .O(N__36316),
            .I(N__36310));
    Span4Mux_h I__7511 (
            .O(N__36313),
            .I(N__36307));
    LocalMux I__7510 (
            .O(N__36310),
            .I(N__36304));
    Span4Mux_h I__7509 (
            .O(N__36307),
            .I(N__36301));
    Span12Mux_v I__7508 (
            .O(N__36304),
            .I(N__36298));
    Odrv4 I__7507 (
            .O(N__36301),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    Odrv12 I__7506 (
            .O(N__36298),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    InMux I__7505 (
            .O(N__36293),
            .I(N__36290));
    LocalMux I__7504 (
            .O(N__36290),
            .I(N__36287));
    Span4Mux_v I__7503 (
            .O(N__36287),
            .I(N__36284));
    Span4Mux_v I__7502 (
            .O(N__36284),
            .I(N__36280));
    InMux I__7501 (
            .O(N__36283),
            .I(N__36277));
    Span4Mux_v I__7500 (
            .O(N__36280),
            .I(N__36274));
    LocalMux I__7499 (
            .O(N__36277),
            .I(state_ns_i_a3_1));
    Odrv4 I__7498 (
            .O(N__36274),
            .I(state_ns_i_a3_1));
    InMux I__7497 (
            .O(N__36269),
            .I(bfn_14_16_0_));
    InMux I__7496 (
            .O(N__36266),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    InMux I__7495 (
            .O(N__36263),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    InMux I__7494 (
            .O(N__36260),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    InMux I__7493 (
            .O(N__36257),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    InMux I__7492 (
            .O(N__36254),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    InMux I__7491 (
            .O(N__36251),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    InMux I__7490 (
            .O(N__36248),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    InMux I__7489 (
            .O(N__36245),
            .I(bfn_14_17_0_));
    InMux I__7488 (
            .O(N__36242),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    InMux I__7487 (
            .O(N__36239),
            .I(bfn_14_15_0_));
    InMux I__7486 (
            .O(N__36236),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    InMux I__7485 (
            .O(N__36233),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    InMux I__7484 (
            .O(N__36230),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    InMux I__7483 (
            .O(N__36227),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    InMux I__7482 (
            .O(N__36224),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    InMux I__7481 (
            .O(N__36221),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    InMux I__7480 (
            .O(N__36218),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    InMux I__7479 (
            .O(N__36215),
            .I(N__36209));
    InMux I__7478 (
            .O(N__36214),
            .I(N__36202));
    InMux I__7477 (
            .O(N__36213),
            .I(N__36202));
    InMux I__7476 (
            .O(N__36212),
            .I(N__36202));
    LocalMux I__7475 (
            .O(N__36209),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    LocalMux I__7474 (
            .O(N__36202),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    InMux I__7473 (
            .O(N__36197),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ));
    InMux I__7472 (
            .O(N__36194),
            .I(N__36160));
    InMux I__7471 (
            .O(N__36193),
            .I(N__36160));
    InMux I__7470 (
            .O(N__36192),
            .I(N__36160));
    InMux I__7469 (
            .O(N__36191),
            .I(N__36160));
    InMux I__7468 (
            .O(N__36190),
            .I(N__36151));
    InMux I__7467 (
            .O(N__36189),
            .I(N__36151));
    InMux I__7466 (
            .O(N__36188),
            .I(N__36151));
    InMux I__7465 (
            .O(N__36187),
            .I(N__36151));
    InMux I__7464 (
            .O(N__36186),
            .I(N__36142));
    InMux I__7463 (
            .O(N__36185),
            .I(N__36142));
    InMux I__7462 (
            .O(N__36184),
            .I(N__36142));
    InMux I__7461 (
            .O(N__36183),
            .I(N__36142));
    InMux I__7460 (
            .O(N__36182),
            .I(N__36135));
    InMux I__7459 (
            .O(N__36181),
            .I(N__36135));
    InMux I__7458 (
            .O(N__36180),
            .I(N__36135));
    InMux I__7457 (
            .O(N__36179),
            .I(N__36126));
    InMux I__7456 (
            .O(N__36178),
            .I(N__36126));
    InMux I__7455 (
            .O(N__36177),
            .I(N__36126));
    InMux I__7454 (
            .O(N__36176),
            .I(N__36126));
    InMux I__7453 (
            .O(N__36175),
            .I(N__36113));
    InMux I__7452 (
            .O(N__36174),
            .I(N__36113));
    InMux I__7451 (
            .O(N__36173),
            .I(N__36113));
    InMux I__7450 (
            .O(N__36172),
            .I(N__36104));
    InMux I__7449 (
            .O(N__36171),
            .I(N__36104));
    InMux I__7448 (
            .O(N__36170),
            .I(N__36104));
    InMux I__7447 (
            .O(N__36169),
            .I(N__36104));
    LocalMux I__7446 (
            .O(N__36160),
            .I(N__36093));
    LocalMux I__7445 (
            .O(N__36151),
            .I(N__36093));
    LocalMux I__7444 (
            .O(N__36142),
            .I(N__36093));
    LocalMux I__7443 (
            .O(N__36135),
            .I(N__36093));
    LocalMux I__7442 (
            .O(N__36126),
            .I(N__36093));
    IoInMux I__7441 (
            .O(N__36125),
            .I(N__36090));
    InMux I__7440 (
            .O(N__36124),
            .I(N__36081));
    InMux I__7439 (
            .O(N__36123),
            .I(N__36081));
    InMux I__7438 (
            .O(N__36122),
            .I(N__36081));
    InMux I__7437 (
            .O(N__36121),
            .I(N__36081));
    InMux I__7436 (
            .O(N__36120),
            .I(N__36078));
    LocalMux I__7435 (
            .O(N__36113),
            .I(N__36071));
    LocalMux I__7434 (
            .O(N__36104),
            .I(N__36071));
    Span4Mux_v I__7433 (
            .O(N__36093),
            .I(N__36071));
    LocalMux I__7432 (
            .O(N__36090),
            .I(N__36068));
    LocalMux I__7431 (
            .O(N__36081),
            .I(N__36065));
    LocalMux I__7430 (
            .O(N__36078),
            .I(N__36060));
    Span4Mux_v I__7429 (
            .O(N__36071),
            .I(N__36060));
    IoSpan4Mux I__7428 (
            .O(N__36068),
            .I(N__36057));
    Odrv12 I__7427 (
            .O(N__36065),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv4 I__7426 (
            .O(N__36060),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv4 I__7425 (
            .O(N__36057),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    InMux I__7424 (
            .O(N__36050),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ));
    CascadeMux I__7423 (
            .O(N__36047),
            .I(N__36042));
    CascadeMux I__7422 (
            .O(N__36046),
            .I(N__36038));
    InMux I__7421 (
            .O(N__36045),
            .I(N__36035));
    InMux I__7420 (
            .O(N__36042),
            .I(N__36028));
    InMux I__7419 (
            .O(N__36041),
            .I(N__36028));
    InMux I__7418 (
            .O(N__36038),
            .I(N__36028));
    LocalMux I__7417 (
            .O(N__36035),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    LocalMux I__7416 (
            .O(N__36028),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    InMux I__7415 (
            .O(N__36023),
            .I(bfn_14_14_0_));
    InMux I__7414 (
            .O(N__36020),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    InMux I__7413 (
            .O(N__36017),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    InMux I__7412 (
            .O(N__36014),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    InMux I__7411 (
            .O(N__36011),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    InMux I__7410 (
            .O(N__36008),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    InMux I__7409 (
            .O(N__36005),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    InMux I__7408 (
            .O(N__36002),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ));
    InMux I__7407 (
            .O(N__35999),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ));
    InMux I__7406 (
            .O(N__35996),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ));
    InMux I__7405 (
            .O(N__35993),
            .I(bfn_14_13_0_));
    InMux I__7404 (
            .O(N__35990),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ));
    InMux I__7403 (
            .O(N__35987),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ));
    CascadeMux I__7402 (
            .O(N__35984),
            .I(N__35979));
    InMux I__7401 (
            .O(N__35983),
            .I(N__35976));
    InMux I__7400 (
            .O(N__35982),
            .I(N__35971));
    InMux I__7399 (
            .O(N__35979),
            .I(N__35971));
    LocalMux I__7398 (
            .O(N__35976),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    LocalMux I__7397 (
            .O(N__35971),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    InMux I__7396 (
            .O(N__35966),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ));
    CascadeMux I__7395 (
            .O(N__35963),
            .I(N__35959));
    InMux I__7394 (
            .O(N__35962),
            .I(N__35955));
    InMux I__7393 (
            .O(N__35959),
            .I(N__35952));
    InMux I__7392 (
            .O(N__35958),
            .I(N__35949));
    LocalMux I__7391 (
            .O(N__35955),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    LocalMux I__7390 (
            .O(N__35952),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    LocalMux I__7389 (
            .O(N__35949),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    InMux I__7388 (
            .O(N__35942),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ));
    InMux I__7387 (
            .O(N__35939),
            .I(N__35935));
    InMux I__7386 (
            .O(N__35938),
            .I(N__35932));
    LocalMux I__7385 (
            .O(N__35935),
            .I(N__35929));
    LocalMux I__7384 (
            .O(N__35932),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__7383 (
            .O(N__35929),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__7382 (
            .O(N__35924),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__7381 (
            .O(N__35921),
            .I(N__35917));
    InMux I__7380 (
            .O(N__35920),
            .I(N__35914));
    LocalMux I__7379 (
            .O(N__35917),
            .I(N__35911));
    LocalMux I__7378 (
            .O(N__35914),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__7377 (
            .O(N__35911),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__7376 (
            .O(N__35906),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__7375 (
            .O(N__35903),
            .I(N__35899));
    InMux I__7374 (
            .O(N__35902),
            .I(N__35896));
    LocalMux I__7373 (
            .O(N__35899),
            .I(N__35893));
    LocalMux I__7372 (
            .O(N__35896),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv12 I__7371 (
            .O(N__35893),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__7370 (
            .O(N__35888),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ));
    CascadeMux I__7369 (
            .O(N__35885),
            .I(N__35880));
    InMux I__7368 (
            .O(N__35884),
            .I(N__35877));
    InMux I__7367 (
            .O(N__35883),
            .I(N__35872));
    InMux I__7366 (
            .O(N__35880),
            .I(N__35872));
    LocalMux I__7365 (
            .O(N__35877),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    LocalMux I__7364 (
            .O(N__35872),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__7363 (
            .O(N__35867),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__7362 (
            .O(N__35864),
            .I(N__35859));
    InMux I__7361 (
            .O(N__35863),
            .I(N__35856));
    InMux I__7360 (
            .O(N__35862),
            .I(N__35853));
    LocalMux I__7359 (
            .O(N__35859),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__7358 (
            .O(N__35856),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__7357 (
            .O(N__35853),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__7356 (
            .O(N__35846),
            .I(bfn_14_12_0_));
    InMux I__7355 (
            .O(N__35843),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ));
    InMux I__7354 (
            .O(N__35840),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ));
    InMux I__7353 (
            .O(N__35837),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ));
    InMux I__7352 (
            .O(N__35834),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__7351 (
            .O(N__35831),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__7350 (
            .O(N__35828),
            .I(N__35825));
    LocalMux I__7349 (
            .O(N__35825),
            .I(N__35821));
    InMux I__7348 (
            .O(N__35824),
            .I(N__35818));
    Span4Mux_v I__7347 (
            .O(N__35821),
            .I(N__35815));
    LocalMux I__7346 (
            .O(N__35818),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    Odrv4 I__7345 (
            .O(N__35815),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__7344 (
            .O(N__35810),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ));
    InMux I__7343 (
            .O(N__35807),
            .I(N__35803));
    InMux I__7342 (
            .O(N__35806),
            .I(N__35800));
    LocalMux I__7341 (
            .O(N__35803),
            .I(N__35797));
    LocalMux I__7340 (
            .O(N__35800),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    Odrv4 I__7339 (
            .O(N__35797),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__7338 (
            .O(N__35792),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__7337 (
            .O(N__35789),
            .I(N__35785));
    InMux I__7336 (
            .O(N__35788),
            .I(N__35782));
    LocalMux I__7335 (
            .O(N__35785),
            .I(N__35779));
    LocalMux I__7334 (
            .O(N__35782),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv12 I__7333 (
            .O(N__35779),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__7332 (
            .O(N__35774),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__7331 (
            .O(N__35771),
            .I(N__35767));
    InMux I__7330 (
            .O(N__35770),
            .I(N__35764));
    LocalMux I__7329 (
            .O(N__35767),
            .I(N__35761));
    LocalMux I__7328 (
            .O(N__35764),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    Odrv12 I__7327 (
            .O(N__35761),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__7326 (
            .O(N__35756),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__7325 (
            .O(N__35753),
            .I(N__35749));
    InMux I__7324 (
            .O(N__35752),
            .I(N__35746));
    LocalMux I__7323 (
            .O(N__35749),
            .I(N__35743));
    LocalMux I__7322 (
            .O(N__35746),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__7321 (
            .O(N__35743),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__7320 (
            .O(N__35738),
            .I(bfn_14_11_0_));
    InMux I__7319 (
            .O(N__35735),
            .I(N__35731));
    InMux I__7318 (
            .O(N__35734),
            .I(N__35728));
    LocalMux I__7317 (
            .O(N__35731),
            .I(N__35725));
    LocalMux I__7316 (
            .O(N__35728),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv4 I__7315 (
            .O(N__35725),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__7314 (
            .O(N__35720),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__7313 (
            .O(N__35717),
            .I(N__35713));
    InMux I__7312 (
            .O(N__35716),
            .I(N__35710));
    LocalMux I__7311 (
            .O(N__35713),
            .I(N__35707));
    LocalMux I__7310 (
            .O(N__35710),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv4 I__7309 (
            .O(N__35707),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__7308 (
            .O(N__35702),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__7307 (
            .O(N__35699),
            .I(N__35695));
    InMux I__7306 (
            .O(N__35698),
            .I(N__35692));
    LocalMux I__7305 (
            .O(N__35695),
            .I(N__35689));
    LocalMux I__7304 (
            .O(N__35692),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__7303 (
            .O(N__35689),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__7302 (
            .O(N__35684),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__7301 (
            .O(N__35681),
            .I(N__35678));
    LocalMux I__7300 (
            .O(N__35678),
            .I(N__35675));
    Span4Mux_h I__7299 (
            .O(N__35675),
            .I(N__35672));
    Odrv4 I__7298 (
            .O(N__35672),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt28 ));
    CascadeMux I__7297 (
            .O(N__35669),
            .I(N__35666));
    InMux I__7296 (
            .O(N__35666),
            .I(N__35663));
    LocalMux I__7295 (
            .O(N__35663),
            .I(N__35660));
    Span4Mux_h I__7294 (
            .O(N__35660),
            .I(N__35657));
    Odrv4 I__7293 (
            .O(N__35657),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ));
    InMux I__7292 (
            .O(N__35654),
            .I(N__35651));
    LocalMux I__7291 (
            .O(N__35651),
            .I(N__35648));
    Span4Mux_v I__7290 (
            .O(N__35648),
            .I(N__35645));
    Odrv4 I__7289 (
            .O(N__35645),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ));
    CascadeMux I__7288 (
            .O(N__35642),
            .I(N__35639));
    InMux I__7287 (
            .O(N__35639),
            .I(N__35635));
    CascadeMux I__7286 (
            .O(N__35638),
            .I(N__35632));
    LocalMux I__7285 (
            .O(N__35635),
            .I(N__35629));
    InMux I__7284 (
            .O(N__35632),
            .I(N__35626));
    Span4Mux_v I__7283 (
            .O(N__35629),
            .I(N__35623));
    LocalMux I__7282 (
            .O(N__35626),
            .I(N__35620));
    Odrv4 I__7281 (
            .O(N__35623),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt30 ));
    Odrv12 I__7280 (
            .O(N__35620),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt30 ));
    InMux I__7279 (
            .O(N__35615),
            .I(N__35612));
    LocalMux I__7278 (
            .O(N__35612),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO ));
    InMux I__7277 (
            .O(N__35609),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ));
    InMux I__7276 (
            .O(N__35606),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30 ));
    InMux I__7275 (
            .O(N__35603),
            .I(N__35600));
    LocalMux I__7274 (
            .O(N__35600),
            .I(N__35596));
    InMux I__7273 (
            .O(N__35599),
            .I(N__35593));
    Span4Mux_v I__7272 (
            .O(N__35596),
            .I(N__35590));
    LocalMux I__7271 (
            .O(N__35593),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ));
    Odrv4 I__7270 (
            .O(N__35590),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ));
    InMux I__7269 (
            .O(N__35585),
            .I(N__35582));
    LocalMux I__7268 (
            .O(N__35582),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ));
    CascadeMux I__7267 (
            .O(N__35579),
            .I(N__35575));
    CascadeMux I__7266 (
            .O(N__35578),
            .I(N__35572));
    InMux I__7265 (
            .O(N__35575),
            .I(N__35569));
    InMux I__7264 (
            .O(N__35572),
            .I(N__35565));
    LocalMux I__7263 (
            .O(N__35569),
            .I(N__35562));
    InMux I__7262 (
            .O(N__35568),
            .I(N__35559));
    LocalMux I__7261 (
            .O(N__35565),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv12 I__7260 (
            .O(N__35562),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__7259 (
            .O(N__35559),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__7258 (
            .O(N__35552),
            .I(N__35548));
    InMux I__7257 (
            .O(N__35551),
            .I(N__35545));
    LocalMux I__7256 (
            .O(N__35548),
            .I(N__35542));
    LocalMux I__7255 (
            .O(N__35545),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    Odrv4 I__7254 (
            .O(N__35542),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__7253 (
            .O(N__35537),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ));
    CascadeMux I__7252 (
            .O(N__35534),
            .I(N__35531));
    InMux I__7251 (
            .O(N__35531),
            .I(N__35528));
    LocalMux I__7250 (
            .O(N__35528),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28 ));
    InMux I__7249 (
            .O(N__35525),
            .I(N__35521));
    InMux I__7248 (
            .O(N__35524),
            .I(N__35518));
    LocalMux I__7247 (
            .O(N__35521),
            .I(N__35515));
    LocalMux I__7246 (
            .O(N__35518),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    Odrv4 I__7245 (
            .O(N__35515),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__7244 (
            .O(N__35510),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__7243 (
            .O(N__35507),
            .I(N__35503));
    InMux I__7242 (
            .O(N__35506),
            .I(N__35500));
    LocalMux I__7241 (
            .O(N__35503),
            .I(N__35497));
    LocalMux I__7240 (
            .O(N__35500),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    Odrv4 I__7239 (
            .O(N__35497),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    CascadeMux I__7238 (
            .O(N__35492),
            .I(N__35489));
    InMux I__7237 (
            .O(N__35489),
            .I(N__35486));
    LocalMux I__7236 (
            .O(N__35486),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ));
    InMux I__7235 (
            .O(N__35483),
            .I(N__35480));
    LocalMux I__7234 (
            .O(N__35480),
            .I(N__35477));
    Span4Mux_h I__7233 (
            .O(N__35477),
            .I(N__35474));
    Span4Mux_v I__7232 (
            .O(N__35474),
            .I(N__35471));
    Odrv4 I__7231 (
            .O(N__35471),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ));
    CascadeMux I__7230 (
            .O(N__35468),
            .I(N__35465));
    InMux I__7229 (
            .O(N__35465),
            .I(N__35462));
    LocalMux I__7228 (
            .O(N__35462),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ));
    InMux I__7227 (
            .O(N__35459),
            .I(N__35456));
    LocalMux I__7226 (
            .O(N__35456),
            .I(N__35453));
    Span4Mux_v I__7225 (
            .O(N__35453),
            .I(N__35450));
    Odrv4 I__7224 (
            .O(N__35450),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ));
    CascadeMux I__7223 (
            .O(N__35447),
            .I(N__35444));
    InMux I__7222 (
            .O(N__35444),
            .I(N__35441));
    LocalMux I__7221 (
            .O(N__35441),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ));
    InMux I__7220 (
            .O(N__35438),
            .I(N__35435));
    LocalMux I__7219 (
            .O(N__35435),
            .I(N__35432));
    Span4Mux_h I__7218 (
            .O(N__35432),
            .I(N__35429));
    Odrv4 I__7217 (
            .O(N__35429),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ));
    CascadeMux I__7216 (
            .O(N__35426),
            .I(N__35423));
    InMux I__7215 (
            .O(N__35423),
            .I(N__35420));
    LocalMux I__7214 (
            .O(N__35420),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ));
    InMux I__7213 (
            .O(N__35417),
            .I(N__35414));
    LocalMux I__7212 (
            .O(N__35414),
            .I(N__35411));
    Odrv4 I__7211 (
            .O(N__35411),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt16 ));
    CascadeMux I__7210 (
            .O(N__35408),
            .I(N__35405));
    InMux I__7209 (
            .O(N__35405),
            .I(N__35402));
    LocalMux I__7208 (
            .O(N__35402),
            .I(N__35399));
    Span4Mux_h I__7207 (
            .O(N__35399),
            .I(N__35396));
    Odrv4 I__7206 (
            .O(N__35396),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ));
    CascadeMux I__7205 (
            .O(N__35393),
            .I(N__35390));
    InMux I__7204 (
            .O(N__35390),
            .I(N__35387));
    LocalMux I__7203 (
            .O(N__35387),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ));
    CascadeMux I__7202 (
            .O(N__35384),
            .I(N__35381));
    InMux I__7201 (
            .O(N__35381),
            .I(N__35378));
    LocalMux I__7200 (
            .O(N__35378),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ));
    InMux I__7199 (
            .O(N__35375),
            .I(N__35372));
    LocalMux I__7198 (
            .O(N__35372),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ));
    InMux I__7197 (
            .O(N__35369),
            .I(N__35366));
    LocalMux I__7196 (
            .O(N__35366),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ));
    CascadeMux I__7195 (
            .O(N__35363),
            .I(N__35360));
    InMux I__7194 (
            .O(N__35360),
            .I(N__35357));
    LocalMux I__7193 (
            .O(N__35357),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ));
    CascadeMux I__7192 (
            .O(N__35354),
            .I(N__35351));
    InMux I__7191 (
            .O(N__35351),
            .I(N__35348));
    LocalMux I__7190 (
            .O(N__35348),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ));
    CascadeMux I__7189 (
            .O(N__35345),
            .I(N__35342));
    InMux I__7188 (
            .O(N__35342),
            .I(N__35339));
    LocalMux I__7187 (
            .O(N__35339),
            .I(N__35336));
    Odrv4 I__7186 (
            .O(N__35336),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ));
    CascadeMux I__7185 (
            .O(N__35333),
            .I(N__35330));
    InMux I__7184 (
            .O(N__35330),
            .I(N__35327));
    LocalMux I__7183 (
            .O(N__35327),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ));
    CascadeMux I__7182 (
            .O(N__35324),
            .I(N__35316));
    CascadeMux I__7181 (
            .O(N__35323),
            .I(N__35312));
    CascadeMux I__7180 (
            .O(N__35322),
            .I(N__35308));
    InMux I__7179 (
            .O(N__35321),
            .I(N__35303));
    InMux I__7178 (
            .O(N__35320),
            .I(N__35303));
    InMux I__7177 (
            .O(N__35319),
            .I(N__35290));
    InMux I__7176 (
            .O(N__35316),
            .I(N__35290));
    InMux I__7175 (
            .O(N__35315),
            .I(N__35290));
    InMux I__7174 (
            .O(N__35312),
            .I(N__35290));
    InMux I__7173 (
            .O(N__35311),
            .I(N__35290));
    InMux I__7172 (
            .O(N__35308),
            .I(N__35290));
    LocalMux I__7171 (
            .O(N__35303),
            .I(N__35287));
    LocalMux I__7170 (
            .O(N__35290),
            .I(N__35284));
    Span12Mux_h I__7169 (
            .O(N__35287),
            .I(N__35279));
    Span12Mux_s7_v I__7168 (
            .O(N__35284),
            .I(N__35279));
    Span12Mux_h I__7167 (
            .O(N__35279),
            .I(N__35276));
    Odrv12 I__7166 (
            .O(N__35276),
            .I(\pwm_generator_inst.un2_threshold_1_25 ));
    CascadeMux I__7165 (
            .O(N__35273),
            .I(N__35270));
    InMux I__7164 (
            .O(N__35270),
            .I(N__35267));
    LocalMux I__7163 (
            .O(N__35267),
            .I(N__35264));
    Span4Mux_s2_v I__7162 (
            .O(N__35264),
            .I(N__35261));
    Span4Mux_v I__7161 (
            .O(N__35261),
            .I(N__35258));
    Odrv4 I__7160 (
            .O(N__35258),
            .I(\pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ));
    InMux I__7159 (
            .O(N__35255),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_14 ));
    InMux I__7158 (
            .O(N__35252),
            .I(N__35249));
    LocalMux I__7157 (
            .O(N__35249),
            .I(N__35246));
    Span4Mux_v I__7156 (
            .O(N__35246),
            .I(N__35243));
    Odrv4 I__7155 (
            .O(N__35243),
            .I(\pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ));
    InMux I__7154 (
            .O(N__35240),
            .I(bfn_13_30_0_));
    CascadeMux I__7153 (
            .O(N__35237),
            .I(N__35233));
    InMux I__7152 (
            .O(N__35236),
            .I(N__35230));
    InMux I__7151 (
            .O(N__35233),
            .I(N__35227));
    LocalMux I__7150 (
            .O(N__35230),
            .I(N__35224));
    LocalMux I__7149 (
            .O(N__35227),
            .I(N__35219));
    Span4Mux_h I__7148 (
            .O(N__35224),
            .I(N__35219));
    Span4Mux_v I__7147 (
            .O(N__35219),
            .I(N__35213));
    InMux I__7146 (
            .O(N__35218),
            .I(N__35206));
    InMux I__7145 (
            .O(N__35217),
            .I(N__35206));
    InMux I__7144 (
            .O(N__35216),
            .I(N__35206));
    Odrv4 I__7143 (
            .O(N__35213),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    LocalMux I__7142 (
            .O(N__35206),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    InMux I__7141 (
            .O(N__35201),
            .I(N__35198));
    LocalMux I__7140 (
            .O(N__35198),
            .I(N__35195));
    Span4Mux_h I__7139 (
            .O(N__35195),
            .I(N__35192));
    Span4Mux_v I__7138 (
            .O(N__35192),
            .I(N__35186));
    InMux I__7137 (
            .O(N__35191),
            .I(N__35179));
    InMux I__7136 (
            .O(N__35190),
            .I(N__35179));
    InMux I__7135 (
            .O(N__35189),
            .I(N__35179));
    Odrv4 I__7134 (
            .O(N__35186),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    LocalMux I__7133 (
            .O(N__35179),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    InMux I__7132 (
            .O(N__35174),
            .I(N__35169));
    InMux I__7131 (
            .O(N__35173),
            .I(N__35166));
    CascadeMux I__7130 (
            .O(N__35172),
            .I(N__35163));
    LocalMux I__7129 (
            .O(N__35169),
            .I(N__35158));
    LocalMux I__7128 (
            .O(N__35166),
            .I(N__35158));
    InMux I__7127 (
            .O(N__35163),
            .I(N__35153));
    Span4Mux_h I__7126 (
            .O(N__35158),
            .I(N__35150));
    InMux I__7125 (
            .O(N__35157),
            .I(N__35145));
    InMux I__7124 (
            .O(N__35156),
            .I(N__35145));
    LocalMux I__7123 (
            .O(N__35153),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    Odrv4 I__7122 (
            .O(N__35150),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    LocalMux I__7121 (
            .O(N__35145),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    InMux I__7120 (
            .O(N__35138),
            .I(N__35135));
    LocalMux I__7119 (
            .O(N__35135),
            .I(N__35132));
    Span4Mux_h I__7118 (
            .O(N__35132),
            .I(N__35128));
    InMux I__7117 (
            .O(N__35131),
            .I(N__35125));
    Odrv4 I__7116 (
            .O(N__35128),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    LocalMux I__7115 (
            .O(N__35125),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    InMux I__7114 (
            .O(N__35120),
            .I(N__35117));
    LocalMux I__7113 (
            .O(N__35117),
            .I(N__35113));
    InMux I__7112 (
            .O(N__35116),
            .I(N__35110));
    Span4Mux_v I__7111 (
            .O(N__35113),
            .I(N__35107));
    LocalMux I__7110 (
            .O(N__35110),
            .I(N__35104));
    Span4Mux_v I__7109 (
            .O(N__35107),
            .I(N__35101));
    Span4Mux_h I__7108 (
            .O(N__35104),
            .I(N__35098));
    Odrv4 I__7107 (
            .O(N__35101),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ));
    Odrv4 I__7106 (
            .O(N__35098),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ));
    CascadeMux I__7105 (
            .O(N__35093),
            .I(N__35089));
    InMux I__7104 (
            .O(N__35092),
            .I(N__35086));
    InMux I__7103 (
            .O(N__35089),
            .I(N__35083));
    LocalMux I__7102 (
            .O(N__35086),
            .I(N__35080));
    LocalMux I__7101 (
            .O(N__35083),
            .I(N__35077));
    Span12Mux_h I__7100 (
            .O(N__35080),
            .I(N__35071));
    Span4Mux_v I__7099 (
            .O(N__35077),
            .I(N__35068));
    InMux I__7098 (
            .O(N__35076),
            .I(N__35063));
    InMux I__7097 (
            .O(N__35075),
            .I(N__35063));
    InMux I__7096 (
            .O(N__35074),
            .I(N__35060));
    Span12Mux_v I__7095 (
            .O(N__35071),
            .I(N__35057));
    Span4Mux_v I__7094 (
            .O(N__35068),
            .I(N__35052));
    LocalMux I__7093 (
            .O(N__35063),
            .I(N__35052));
    LocalMux I__7092 (
            .O(N__35060),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    Odrv12 I__7091 (
            .O(N__35057),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    Odrv4 I__7090 (
            .O(N__35052),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    CascadeMux I__7089 (
            .O(N__35045),
            .I(N__35042));
    InMux I__7088 (
            .O(N__35042),
            .I(N__35038));
    InMux I__7087 (
            .O(N__35041),
            .I(N__35035));
    LocalMux I__7086 (
            .O(N__35038),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    LocalMux I__7085 (
            .O(N__35035),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    CascadeMux I__7084 (
            .O(N__35030),
            .I(N__35027));
    InMux I__7083 (
            .O(N__35027),
            .I(N__35024));
    LocalMux I__7082 (
            .O(N__35024),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ));
    InMux I__7081 (
            .O(N__35021),
            .I(N__35018));
    LocalMux I__7080 (
            .O(N__35018),
            .I(N__35015));
    Span4Mux_v I__7079 (
            .O(N__35015),
            .I(N__35012));
    Odrv4 I__7078 (
            .O(N__35012),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ));
    CascadeMux I__7077 (
            .O(N__35009),
            .I(N__35006));
    InMux I__7076 (
            .O(N__35006),
            .I(N__35003));
    LocalMux I__7075 (
            .O(N__35003),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ));
    InMux I__7074 (
            .O(N__35000),
            .I(N__34997));
    LocalMux I__7073 (
            .O(N__34997),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ));
    InMux I__7072 (
            .O(N__34994),
            .I(N__34991));
    LocalMux I__7071 (
            .O(N__34991),
            .I(N__34988));
    Span4Mux_v I__7070 (
            .O(N__34988),
            .I(N__34985));
    Sp12to4 I__7069 (
            .O(N__34985),
            .I(N__34982));
    Span12Mux_h I__7068 (
            .O(N__34982),
            .I(N__34979));
    Odrv12 I__7067 (
            .O(N__34979),
            .I(\pwm_generator_inst.un2_threshold_2_7 ));
    CascadeMux I__7066 (
            .O(N__34976),
            .I(N__34973));
    InMux I__7065 (
            .O(N__34973),
            .I(N__34970));
    LocalMux I__7064 (
            .O(N__34970),
            .I(N__34967));
    Span4Mux_v I__7063 (
            .O(N__34967),
            .I(N__34964));
    Sp12to4 I__7062 (
            .O(N__34964),
            .I(N__34961));
    Odrv12 I__7061 (
            .O(N__34961),
            .I(\pwm_generator_inst.un2_threshold_1_22 ));
    InMux I__7060 (
            .O(N__34958),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_6 ));
    InMux I__7059 (
            .O(N__34955),
            .I(N__34952));
    LocalMux I__7058 (
            .O(N__34952),
            .I(N__34949));
    Span4Mux_v I__7057 (
            .O(N__34949),
            .I(N__34946));
    Span4Mux_h I__7056 (
            .O(N__34946),
            .I(N__34943));
    Span4Mux_h I__7055 (
            .O(N__34943),
            .I(N__34940));
    Span4Mux_h I__7054 (
            .O(N__34940),
            .I(N__34937));
    Odrv4 I__7053 (
            .O(N__34937),
            .I(\pwm_generator_inst.un2_threshold_2_8 ));
    CascadeMux I__7052 (
            .O(N__34934),
            .I(N__34931));
    InMux I__7051 (
            .O(N__34931),
            .I(N__34928));
    LocalMux I__7050 (
            .O(N__34928),
            .I(N__34925));
    Span12Mux_s10_v I__7049 (
            .O(N__34925),
            .I(N__34922));
    Span12Mux_h I__7048 (
            .O(N__34922),
            .I(N__34919));
    Odrv12 I__7047 (
            .O(N__34919),
            .I(\pwm_generator_inst.un2_threshold_1_23 ));
    InMux I__7046 (
            .O(N__34916),
            .I(bfn_13_29_0_));
    InMux I__7045 (
            .O(N__34913),
            .I(N__34910));
    LocalMux I__7044 (
            .O(N__34910),
            .I(N__34907));
    Span4Mux_v I__7043 (
            .O(N__34907),
            .I(N__34904));
    Span4Mux_h I__7042 (
            .O(N__34904),
            .I(N__34901));
    Span4Mux_h I__7041 (
            .O(N__34901),
            .I(N__34898));
    Span4Mux_h I__7040 (
            .O(N__34898),
            .I(N__34895));
    Odrv4 I__7039 (
            .O(N__34895),
            .I(\pwm_generator_inst.un2_threshold_2_9 ));
    CascadeMux I__7038 (
            .O(N__34892),
            .I(N__34889));
    InMux I__7037 (
            .O(N__34889),
            .I(N__34886));
    LocalMux I__7036 (
            .O(N__34886),
            .I(N__34883));
    Span12Mux_s8_v I__7035 (
            .O(N__34883),
            .I(N__34880));
    Span12Mux_h I__7034 (
            .O(N__34880),
            .I(N__34877));
    Odrv12 I__7033 (
            .O(N__34877),
            .I(\pwm_generator_inst.un2_threshold_1_24 ));
    InMux I__7032 (
            .O(N__34874),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_8 ));
    InMux I__7031 (
            .O(N__34871),
            .I(N__34868));
    LocalMux I__7030 (
            .O(N__34868),
            .I(N__34865));
    Span4Mux_v I__7029 (
            .O(N__34865),
            .I(N__34862));
    Sp12to4 I__7028 (
            .O(N__34862),
            .I(N__34859));
    Span12Mux_h I__7027 (
            .O(N__34859),
            .I(N__34856));
    Odrv12 I__7026 (
            .O(N__34856),
            .I(\pwm_generator_inst.un2_threshold_2_10 ));
    InMux I__7025 (
            .O(N__34853),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_9 ));
    CascadeMux I__7024 (
            .O(N__34850),
            .I(N__34847));
    InMux I__7023 (
            .O(N__34847),
            .I(N__34844));
    LocalMux I__7022 (
            .O(N__34844),
            .I(N__34841));
    Span4Mux_s3_v I__7021 (
            .O(N__34841),
            .I(N__34838));
    Sp12to4 I__7020 (
            .O(N__34838),
            .I(N__34835));
    Span12Mux_h I__7019 (
            .O(N__34835),
            .I(N__34832));
    Odrv12 I__7018 (
            .O(N__34832),
            .I(\pwm_generator_inst.un2_threshold_2_11 ));
    InMux I__7017 (
            .O(N__34829),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_10 ));
    InMux I__7016 (
            .O(N__34826),
            .I(N__34823));
    LocalMux I__7015 (
            .O(N__34823),
            .I(N__34820));
    Span4Mux_s2_v I__7014 (
            .O(N__34820),
            .I(N__34817));
    Span4Mux_v I__7013 (
            .O(N__34817),
            .I(N__34814));
    Sp12to4 I__7012 (
            .O(N__34814),
            .I(N__34811));
    Odrv12 I__7011 (
            .O(N__34811),
            .I(\pwm_generator_inst.un2_threshold_2_12 ));
    InMux I__7010 (
            .O(N__34808),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11 ));
    CascadeMux I__7009 (
            .O(N__34805),
            .I(N__34802));
    InMux I__7008 (
            .O(N__34802),
            .I(N__34799));
    LocalMux I__7007 (
            .O(N__34799),
            .I(N__34796));
    Sp12to4 I__7006 (
            .O(N__34796),
            .I(N__34793));
    Span12Mux_h I__7005 (
            .O(N__34793),
            .I(N__34790));
    Odrv12 I__7004 (
            .O(N__34790),
            .I(\pwm_generator_inst.un2_threshold_2_13 ));
    InMux I__7003 (
            .O(N__34787),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_12 ));
    InMux I__7002 (
            .O(N__34784),
            .I(N__34781));
    LocalMux I__7001 (
            .O(N__34781),
            .I(N__34778));
    Span4Mux_v I__7000 (
            .O(N__34778),
            .I(N__34775));
    Sp12to4 I__6999 (
            .O(N__34775),
            .I(N__34772));
    Span12Mux_h I__6998 (
            .O(N__34772),
            .I(N__34769));
    Odrv12 I__6997 (
            .O(N__34769),
            .I(\pwm_generator_inst.un2_threshold_2_14 ));
    InMux I__6996 (
            .O(N__34766),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_13 ));
    InMux I__6995 (
            .O(N__34763),
            .I(N__34760));
    LocalMux I__6994 (
            .O(N__34760),
            .I(N__34757));
    Odrv12 I__6993 (
            .O(N__34757),
            .I(\pwm_generator_inst.un19_threshold_axb_7 ));
    InMux I__6992 (
            .O(N__34754),
            .I(N__34751));
    LocalMux I__6991 (
            .O(N__34751),
            .I(N__34748));
    Span4Mux_v I__6990 (
            .O(N__34748),
            .I(N__34745));
    Span4Mux_h I__6989 (
            .O(N__34745),
            .I(N__34742));
    Span4Mux_h I__6988 (
            .O(N__34742),
            .I(N__34739));
    Span4Mux_h I__6987 (
            .O(N__34739),
            .I(N__34736));
    Odrv4 I__6986 (
            .O(N__34736),
            .I(\pwm_generator_inst.un2_threshold_2_0 ));
    CascadeMux I__6985 (
            .O(N__34733),
            .I(N__34730));
    InMux I__6984 (
            .O(N__34730),
            .I(N__34727));
    LocalMux I__6983 (
            .O(N__34727),
            .I(N__34724));
    Span12Mux_s11_v I__6982 (
            .O(N__34724),
            .I(N__34721));
    Span12Mux_h I__6981 (
            .O(N__34721),
            .I(N__34718));
    Odrv12 I__6980 (
            .O(N__34718),
            .I(\pwm_generator_inst.un2_threshold_1_15 ));
    InMux I__6979 (
            .O(N__34715),
            .I(N__34712));
    LocalMux I__6978 (
            .O(N__34712),
            .I(N__34709));
    Span4Mux_v I__6977 (
            .O(N__34709),
            .I(N__34706));
    Sp12to4 I__6976 (
            .O(N__34706),
            .I(N__34703));
    Span12Mux_h I__6975 (
            .O(N__34703),
            .I(N__34700));
    Odrv12 I__6974 (
            .O(N__34700),
            .I(\pwm_generator_inst.un2_threshold_2_1 ));
    CascadeMux I__6973 (
            .O(N__34697),
            .I(N__34694));
    InMux I__6972 (
            .O(N__34694),
            .I(N__34691));
    LocalMux I__6971 (
            .O(N__34691),
            .I(N__34688));
    Span12Mux_s9_v I__6970 (
            .O(N__34688),
            .I(N__34685));
    Span12Mux_h I__6969 (
            .O(N__34685),
            .I(N__34682));
    Odrv12 I__6968 (
            .O(N__34682),
            .I(\pwm_generator_inst.un2_threshold_1_16 ));
    InMux I__6967 (
            .O(N__34679),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_0 ));
    InMux I__6966 (
            .O(N__34676),
            .I(N__34673));
    LocalMux I__6965 (
            .O(N__34673),
            .I(N__34670));
    Span4Mux_v I__6964 (
            .O(N__34670),
            .I(N__34667));
    Span4Mux_h I__6963 (
            .O(N__34667),
            .I(N__34664));
    Span4Mux_h I__6962 (
            .O(N__34664),
            .I(N__34661));
    Span4Mux_h I__6961 (
            .O(N__34661),
            .I(N__34658));
    Odrv4 I__6960 (
            .O(N__34658),
            .I(\pwm_generator_inst.un2_threshold_2_2 ));
    CascadeMux I__6959 (
            .O(N__34655),
            .I(N__34652));
    InMux I__6958 (
            .O(N__34652),
            .I(N__34649));
    LocalMux I__6957 (
            .O(N__34649),
            .I(N__34646));
    Span12Mux_s4_v I__6956 (
            .O(N__34646),
            .I(N__34643));
    Span12Mux_h I__6955 (
            .O(N__34643),
            .I(N__34640));
    Odrv12 I__6954 (
            .O(N__34640),
            .I(\pwm_generator_inst.un2_threshold_1_17 ));
    InMux I__6953 (
            .O(N__34637),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1 ));
    InMux I__6952 (
            .O(N__34634),
            .I(N__34631));
    LocalMux I__6951 (
            .O(N__34631),
            .I(N__34628));
    Span4Mux_v I__6950 (
            .O(N__34628),
            .I(N__34625));
    Sp12to4 I__6949 (
            .O(N__34625),
            .I(N__34622));
    Span12Mux_h I__6948 (
            .O(N__34622),
            .I(N__34619));
    Odrv12 I__6947 (
            .O(N__34619),
            .I(\pwm_generator_inst.un2_threshold_2_3 ));
    CascadeMux I__6946 (
            .O(N__34616),
            .I(N__34613));
    InMux I__6945 (
            .O(N__34613),
            .I(N__34610));
    LocalMux I__6944 (
            .O(N__34610),
            .I(N__34607));
    Span4Mux_h I__6943 (
            .O(N__34607),
            .I(N__34604));
    Span4Mux_h I__6942 (
            .O(N__34604),
            .I(N__34601));
    Span4Mux_h I__6941 (
            .O(N__34601),
            .I(N__34598));
    Odrv4 I__6940 (
            .O(N__34598),
            .I(\pwm_generator_inst.un2_threshold_1_18 ));
    InMux I__6939 (
            .O(N__34595),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2 ));
    InMux I__6938 (
            .O(N__34592),
            .I(N__34589));
    LocalMux I__6937 (
            .O(N__34589),
            .I(N__34586));
    Span4Mux_s3_v I__6936 (
            .O(N__34586),
            .I(N__34583));
    Span4Mux_v I__6935 (
            .O(N__34583),
            .I(N__34580));
    Sp12to4 I__6934 (
            .O(N__34580),
            .I(N__34577));
    Odrv12 I__6933 (
            .O(N__34577),
            .I(\pwm_generator_inst.un2_threshold_2_4 ));
    CascadeMux I__6932 (
            .O(N__34574),
            .I(N__34571));
    InMux I__6931 (
            .O(N__34571),
            .I(N__34568));
    LocalMux I__6930 (
            .O(N__34568),
            .I(N__34565));
    Span12Mux_h I__6929 (
            .O(N__34565),
            .I(N__34562));
    Odrv12 I__6928 (
            .O(N__34562),
            .I(\pwm_generator_inst.un2_threshold_1_19 ));
    InMux I__6927 (
            .O(N__34559),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3 ));
    InMux I__6926 (
            .O(N__34556),
            .I(N__34553));
    LocalMux I__6925 (
            .O(N__34553),
            .I(N__34550));
    Span12Mux_h I__6924 (
            .O(N__34550),
            .I(N__34547));
    Span12Mux_h I__6923 (
            .O(N__34547),
            .I(N__34544));
    Odrv12 I__6922 (
            .O(N__34544),
            .I(\pwm_generator_inst.un2_threshold_2_5 ));
    CascadeMux I__6921 (
            .O(N__34541),
            .I(N__34538));
    InMux I__6920 (
            .O(N__34538),
            .I(N__34535));
    LocalMux I__6919 (
            .O(N__34535),
            .I(N__34532));
    Span4Mux_h I__6918 (
            .O(N__34532),
            .I(N__34529));
    Span4Mux_h I__6917 (
            .O(N__34529),
            .I(N__34526));
    Span4Mux_h I__6916 (
            .O(N__34526),
            .I(N__34523));
    Odrv4 I__6915 (
            .O(N__34523),
            .I(\pwm_generator_inst.un2_threshold_1_20 ));
    InMux I__6914 (
            .O(N__34520),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_4 ));
    InMux I__6913 (
            .O(N__34517),
            .I(N__34514));
    LocalMux I__6912 (
            .O(N__34514),
            .I(N__34511));
    Span4Mux_v I__6911 (
            .O(N__34511),
            .I(N__34508));
    Sp12to4 I__6910 (
            .O(N__34508),
            .I(N__34505));
    Span12Mux_h I__6909 (
            .O(N__34505),
            .I(N__34502));
    Odrv12 I__6908 (
            .O(N__34502),
            .I(\pwm_generator_inst.un2_threshold_2_6 ));
    CascadeMux I__6907 (
            .O(N__34499),
            .I(N__34496));
    InMux I__6906 (
            .O(N__34496),
            .I(N__34493));
    LocalMux I__6905 (
            .O(N__34493),
            .I(N__34490));
    Span4Mux_h I__6904 (
            .O(N__34490),
            .I(N__34487));
    Span4Mux_h I__6903 (
            .O(N__34487),
            .I(N__34484));
    Span4Mux_h I__6902 (
            .O(N__34484),
            .I(N__34481));
    Odrv4 I__6901 (
            .O(N__34481),
            .I(\pwm_generator_inst.un2_threshold_1_21 ));
    InMux I__6900 (
            .O(N__34478),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_5 ));
    InMux I__6899 (
            .O(N__34475),
            .I(\pwm_generator_inst.un19_threshold_cry_8 ));
    InMux I__6898 (
            .O(N__34472),
            .I(N__34469));
    LocalMux I__6897 (
            .O(N__34469),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433 ));
    InMux I__6896 (
            .O(N__34466),
            .I(N__34463));
    LocalMux I__6895 (
            .O(N__34463),
            .I(\pwm_generator_inst.un19_threshold_axb_5 ));
    InMux I__6894 (
            .O(N__34460),
            .I(N__34457));
    LocalMux I__6893 (
            .O(N__34457),
            .I(\pwm_generator_inst.un19_threshold_axb_3 ));
    InMux I__6892 (
            .O(N__34454),
            .I(N__34451));
    LocalMux I__6891 (
            .O(N__34451),
            .I(\pwm_generator_inst.un19_threshold_axb_6 ));
    InMux I__6890 (
            .O(N__34448),
            .I(N__34445));
    LocalMux I__6889 (
            .O(N__34445),
            .I(\pwm_generator_inst.un19_threshold_axb_4 ));
    InMux I__6888 (
            .O(N__34442),
            .I(N__34439));
    LocalMux I__6887 (
            .O(N__34439),
            .I(\pwm_generator_inst.un19_threshold_axb_0 ));
    InMux I__6886 (
            .O(N__34436),
            .I(N__34433));
    LocalMux I__6885 (
            .O(N__34433),
            .I(\pwm_generator_inst.un19_threshold_axb_8 ));
    InMux I__6884 (
            .O(N__34430),
            .I(N__34427));
    LocalMux I__6883 (
            .O(N__34427),
            .I(N__34424));
    Odrv4 I__6882 (
            .O(N__34424),
            .I(\pwm_generator_inst.un19_threshold_axb_2 ));
    CascadeMux I__6881 (
            .O(N__34421),
            .I(N__34418));
    InMux I__6880 (
            .O(N__34418),
            .I(N__34415));
    LocalMux I__6879 (
            .O(N__34415),
            .I(\pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ));
    InMux I__6878 (
            .O(N__34412),
            .I(\pwm_generator_inst.un19_threshold_cry_0 ));
    CascadeMux I__6877 (
            .O(N__34409),
            .I(N__34406));
    InMux I__6876 (
            .O(N__34406),
            .I(N__34403));
    LocalMux I__6875 (
            .O(N__34403),
            .I(\pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ));
    InMux I__6874 (
            .O(N__34400),
            .I(\pwm_generator_inst.un19_threshold_cry_1 ));
    InMux I__6873 (
            .O(N__34397),
            .I(N__34394));
    LocalMux I__6872 (
            .O(N__34394),
            .I(\pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ));
    InMux I__6871 (
            .O(N__34391),
            .I(\pwm_generator_inst.un19_threshold_cry_2 ));
    InMux I__6870 (
            .O(N__34388),
            .I(N__34385));
    LocalMux I__6869 (
            .O(N__34385),
            .I(\pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ));
    InMux I__6868 (
            .O(N__34382),
            .I(\pwm_generator_inst.un19_threshold_cry_3 ));
    CascadeMux I__6867 (
            .O(N__34379),
            .I(N__34376));
    InMux I__6866 (
            .O(N__34376),
            .I(N__34373));
    LocalMux I__6865 (
            .O(N__34373),
            .I(\pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ));
    InMux I__6864 (
            .O(N__34370),
            .I(\pwm_generator_inst.un19_threshold_cry_4 ));
    InMux I__6863 (
            .O(N__34367),
            .I(N__34364));
    LocalMux I__6862 (
            .O(N__34364),
            .I(\pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ));
    InMux I__6861 (
            .O(N__34361),
            .I(\pwm_generator_inst.un19_threshold_cry_5 ));
    InMux I__6860 (
            .O(N__34358),
            .I(N__34355));
    LocalMux I__6859 (
            .O(N__34355),
            .I(\pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ));
    InMux I__6858 (
            .O(N__34352),
            .I(\pwm_generator_inst.un19_threshold_cry_6 ));
    CascadeMux I__6857 (
            .O(N__34349),
            .I(N__34346));
    InMux I__6856 (
            .O(N__34346),
            .I(N__34343));
    LocalMux I__6855 (
            .O(N__34343),
            .I(\pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ));
    InMux I__6854 (
            .O(N__34340),
            .I(bfn_13_25_0_));
    InMux I__6853 (
            .O(N__34337),
            .I(N__34334));
    LocalMux I__6852 (
            .O(N__34334),
            .I(N__34329));
    InMux I__6851 (
            .O(N__34333),
            .I(N__34326));
    InMux I__6850 (
            .O(N__34332),
            .I(N__34323));
    Span4Mux_v I__6849 (
            .O(N__34329),
            .I(N__34320));
    LocalMux I__6848 (
            .O(N__34326),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__6847 (
            .O(N__34323),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    Odrv4 I__6846 (
            .O(N__34320),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__6845 (
            .O(N__34313),
            .I(N__34309));
    InMux I__6844 (
            .O(N__34312),
            .I(N__34305));
    LocalMux I__6843 (
            .O(N__34309),
            .I(N__34302));
    InMux I__6842 (
            .O(N__34308),
            .I(N__34299));
    LocalMux I__6841 (
            .O(N__34305),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    Odrv4 I__6840 (
            .O(N__34302),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__6839 (
            .O(N__34299),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    InMux I__6838 (
            .O(N__34292),
            .I(N__34287));
    InMux I__6837 (
            .O(N__34291),
            .I(N__34284));
    InMux I__6836 (
            .O(N__34290),
            .I(N__34281));
    LocalMux I__6835 (
            .O(N__34287),
            .I(N__34278));
    LocalMux I__6834 (
            .O(N__34284),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__6833 (
            .O(N__34281),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    Odrv4 I__6832 (
            .O(N__34278),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    InMux I__6831 (
            .O(N__34271),
            .I(N__34266));
    InMux I__6830 (
            .O(N__34270),
            .I(N__34263));
    InMux I__6829 (
            .O(N__34269),
            .I(N__34260));
    LocalMux I__6828 (
            .O(N__34266),
            .I(N__34257));
    LocalMux I__6827 (
            .O(N__34263),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__6826 (
            .O(N__34260),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    Odrv4 I__6825 (
            .O(N__34257),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    CascadeMux I__6824 (
            .O(N__34250),
            .I(\pwm_generator_inst.un1_counterlto2_0_cascade_ ));
    InMux I__6823 (
            .O(N__34247),
            .I(N__34242));
    InMux I__6822 (
            .O(N__34246),
            .I(N__34239));
    InMux I__6821 (
            .O(N__34245),
            .I(N__34236));
    LocalMux I__6820 (
            .O(N__34242),
            .I(N__34233));
    LocalMux I__6819 (
            .O(N__34239),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__6818 (
            .O(N__34236),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    Odrv4 I__6817 (
            .O(N__34233),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    InMux I__6816 (
            .O(N__34226),
            .I(N__34210));
    InMux I__6815 (
            .O(N__34225),
            .I(N__34210));
    InMux I__6814 (
            .O(N__34224),
            .I(N__34210));
    InMux I__6813 (
            .O(N__34223),
            .I(N__34210));
    InMux I__6812 (
            .O(N__34222),
            .I(N__34195));
    InMux I__6811 (
            .O(N__34221),
            .I(N__34195));
    InMux I__6810 (
            .O(N__34220),
            .I(N__34195));
    InMux I__6809 (
            .O(N__34219),
            .I(N__34195));
    LocalMux I__6808 (
            .O(N__34210),
            .I(N__34188));
    InMux I__6807 (
            .O(N__34209),
            .I(N__34183));
    InMux I__6806 (
            .O(N__34208),
            .I(N__34183));
    InMux I__6805 (
            .O(N__34207),
            .I(N__34174));
    InMux I__6804 (
            .O(N__34206),
            .I(N__34174));
    InMux I__6803 (
            .O(N__34205),
            .I(N__34174));
    InMux I__6802 (
            .O(N__34204),
            .I(N__34174));
    LocalMux I__6801 (
            .O(N__34195),
            .I(N__34171));
    InMux I__6800 (
            .O(N__34194),
            .I(N__34162));
    InMux I__6799 (
            .O(N__34193),
            .I(N__34162));
    InMux I__6798 (
            .O(N__34192),
            .I(N__34162));
    InMux I__6797 (
            .O(N__34191),
            .I(N__34162));
    Span4Mux_v I__6796 (
            .O(N__34188),
            .I(N__34143));
    LocalMux I__6795 (
            .O(N__34183),
            .I(N__34143));
    LocalMux I__6794 (
            .O(N__34174),
            .I(N__34143));
    Span4Mux_v I__6793 (
            .O(N__34171),
            .I(N__34143));
    LocalMux I__6792 (
            .O(N__34162),
            .I(N__34143));
    InMux I__6791 (
            .O(N__34161),
            .I(N__34134));
    InMux I__6790 (
            .O(N__34160),
            .I(N__34134));
    InMux I__6789 (
            .O(N__34159),
            .I(N__34134));
    InMux I__6788 (
            .O(N__34158),
            .I(N__34134));
    InMux I__6787 (
            .O(N__34157),
            .I(N__34125));
    InMux I__6786 (
            .O(N__34156),
            .I(N__34125));
    InMux I__6785 (
            .O(N__34155),
            .I(N__34125));
    InMux I__6784 (
            .O(N__34154),
            .I(N__34125));
    Span4Mux_v I__6783 (
            .O(N__34143),
            .I(N__34116));
    LocalMux I__6782 (
            .O(N__34134),
            .I(N__34116));
    LocalMux I__6781 (
            .O(N__34125),
            .I(N__34113));
    InMux I__6780 (
            .O(N__34124),
            .I(N__34104));
    InMux I__6779 (
            .O(N__34123),
            .I(N__34104));
    InMux I__6778 (
            .O(N__34122),
            .I(N__34104));
    InMux I__6777 (
            .O(N__34121),
            .I(N__34104));
    Span4Mux_h I__6776 (
            .O(N__34116),
            .I(N__34099));
    Span4Mux_h I__6775 (
            .O(N__34113),
            .I(N__34099));
    LocalMux I__6774 (
            .O(N__34104),
            .I(N__34096));
    Span4Mux_h I__6773 (
            .O(N__34099),
            .I(N__34093));
    Odrv12 I__6772 (
            .O(N__34096),
            .I(\current_shift_inst.timer_s1.running_i ));
    Odrv4 I__6771 (
            .O(N__34093),
            .I(\current_shift_inst.timer_s1.running_i ));
    InMux I__6770 (
            .O(N__34088),
            .I(N__34083));
    InMux I__6769 (
            .O(N__34087),
            .I(N__34080));
    InMux I__6768 (
            .O(N__34086),
            .I(N__34077));
    LocalMux I__6767 (
            .O(N__34083),
            .I(N__34074));
    LocalMux I__6766 (
            .O(N__34080),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__6765 (
            .O(N__34077),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    Odrv4 I__6764 (
            .O(N__34074),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    InMux I__6763 (
            .O(N__34067),
            .I(N__34063));
    InMux I__6762 (
            .O(N__34066),
            .I(N__34059));
    LocalMux I__6761 (
            .O(N__34063),
            .I(N__34056));
    InMux I__6760 (
            .O(N__34062),
            .I(N__34053));
    LocalMux I__6759 (
            .O(N__34059),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    Odrv4 I__6758 (
            .O(N__34056),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__6757 (
            .O(N__34053),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    InMux I__6756 (
            .O(N__34046),
            .I(N__34041));
    InMux I__6755 (
            .O(N__34045),
            .I(N__34038));
    InMux I__6754 (
            .O(N__34044),
            .I(N__34035));
    LocalMux I__6753 (
            .O(N__34041),
            .I(N__34032));
    LocalMux I__6752 (
            .O(N__34038),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__6751 (
            .O(N__34035),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    Odrv4 I__6750 (
            .O(N__34032),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    InMux I__6749 (
            .O(N__34025),
            .I(N__34020));
    InMux I__6748 (
            .O(N__34024),
            .I(N__34017));
    InMux I__6747 (
            .O(N__34023),
            .I(N__34014));
    LocalMux I__6746 (
            .O(N__34020),
            .I(N__34011));
    LocalMux I__6745 (
            .O(N__34017),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__6744 (
            .O(N__34014),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    Odrv4 I__6743 (
            .O(N__34011),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    InMux I__6742 (
            .O(N__34004),
            .I(N__33999));
    InMux I__6741 (
            .O(N__34003),
            .I(N__33996));
    InMux I__6740 (
            .O(N__34002),
            .I(N__33993));
    LocalMux I__6739 (
            .O(N__33999),
            .I(N__33990));
    LocalMux I__6738 (
            .O(N__33996),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__6737 (
            .O(N__33993),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    Odrv4 I__6736 (
            .O(N__33990),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    CascadeMux I__6735 (
            .O(N__33983),
            .I(\pwm_generator_inst.un1_counterlto9_2_cascade_ ));
    InMux I__6734 (
            .O(N__33980),
            .I(N__33977));
    LocalMux I__6733 (
            .O(N__33977),
            .I(\pwm_generator_inst.un1_counterlt9 ));
    InMux I__6732 (
            .O(N__33974),
            .I(N__33956));
    InMux I__6731 (
            .O(N__33973),
            .I(N__33956));
    InMux I__6730 (
            .O(N__33972),
            .I(N__33956));
    InMux I__6729 (
            .O(N__33971),
            .I(N__33956));
    InMux I__6728 (
            .O(N__33970),
            .I(N__33951));
    InMux I__6727 (
            .O(N__33969),
            .I(N__33951));
    InMux I__6726 (
            .O(N__33968),
            .I(N__33942));
    InMux I__6725 (
            .O(N__33967),
            .I(N__33942));
    InMux I__6724 (
            .O(N__33966),
            .I(N__33942));
    InMux I__6723 (
            .O(N__33965),
            .I(N__33942));
    LocalMux I__6722 (
            .O(N__33956),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__6721 (
            .O(N__33951),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__6720 (
            .O(N__33942),
            .I(\pwm_generator_inst.un1_counter_0 ));
    InMux I__6719 (
            .O(N__33935),
            .I(N__33932));
    LocalMux I__6718 (
            .O(N__33932),
            .I(N__33928));
    InMux I__6717 (
            .O(N__33931),
            .I(N__33925));
    Span4Mux_h I__6716 (
            .O(N__33928),
            .I(N__33922));
    LocalMux I__6715 (
            .O(N__33925),
            .I(N__33919));
    Sp12to4 I__6714 (
            .O(N__33922),
            .I(N__33916));
    Span4Mux_s3_h I__6713 (
            .O(N__33919),
            .I(N__33913));
    Span12Mux_v I__6712 (
            .O(N__33916),
            .I(N__33910));
    Span4Mux_h I__6711 (
            .O(N__33913),
            .I(N__33907));
    Odrv12 I__6710 (
            .O(N__33910),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    Odrv4 I__6709 (
            .O(N__33907),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    InMux I__6708 (
            .O(N__33902),
            .I(N__33899));
    LocalMux I__6707 (
            .O(N__33899),
            .I(N__33895));
    InMux I__6706 (
            .O(N__33898),
            .I(N__33892));
    Span4Mux_v I__6705 (
            .O(N__33895),
            .I(N__33889));
    LocalMux I__6704 (
            .O(N__33892),
            .I(N__33886));
    Sp12to4 I__6703 (
            .O(N__33889),
            .I(N__33883));
    Span4Mux_s3_h I__6702 (
            .O(N__33886),
            .I(N__33880));
    Span12Mux_h I__6701 (
            .O(N__33883),
            .I(N__33877));
    Span4Mux_h I__6700 (
            .O(N__33880),
            .I(N__33874));
    Odrv12 I__6699 (
            .O(N__33877),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    Odrv4 I__6698 (
            .O(N__33874),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    InMux I__6697 (
            .O(N__33869),
            .I(N__33866));
    LocalMux I__6696 (
            .O(N__33866),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ));
    CascadeMux I__6695 (
            .O(N__33863),
            .I(N__33860));
    InMux I__6694 (
            .O(N__33860),
            .I(N__33856));
    CascadeMux I__6693 (
            .O(N__33859),
            .I(N__33853));
    LocalMux I__6692 (
            .O(N__33856),
            .I(N__33850));
    InMux I__6691 (
            .O(N__33853),
            .I(N__33845));
    Span4Mux_v I__6690 (
            .O(N__33850),
            .I(N__33842));
    InMux I__6689 (
            .O(N__33849),
            .I(N__33839));
    InMux I__6688 (
            .O(N__33848),
            .I(N__33836));
    LocalMux I__6687 (
            .O(N__33845),
            .I(N__33833));
    Span4Mux_h I__6686 (
            .O(N__33842),
            .I(N__33826));
    LocalMux I__6685 (
            .O(N__33839),
            .I(N__33826));
    LocalMux I__6684 (
            .O(N__33836),
            .I(N__33826));
    Span4Mux_v I__6683 (
            .O(N__33833),
            .I(N__33823));
    Span4Mux_v I__6682 (
            .O(N__33826),
            .I(N__33820));
    Odrv4 I__6681 (
            .O(N__33823),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    Odrv4 I__6680 (
            .O(N__33820),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    InMux I__6679 (
            .O(N__33815),
            .I(N__33812));
    LocalMux I__6678 (
            .O(N__33812),
            .I(N__33807));
    CascadeMux I__6677 (
            .O(N__33811),
            .I(N__33804));
    InMux I__6676 (
            .O(N__33810),
            .I(N__33801));
    Span4Mux_h I__6675 (
            .O(N__33807),
            .I(N__33798));
    InMux I__6674 (
            .O(N__33804),
            .I(N__33795));
    LocalMux I__6673 (
            .O(N__33801),
            .I(\current_shift_inst.un4_control_input1_28 ));
    Odrv4 I__6672 (
            .O(N__33798),
            .I(\current_shift_inst.un4_control_input1_28 ));
    LocalMux I__6671 (
            .O(N__33795),
            .I(\current_shift_inst.un4_control_input1_28 ));
    InMux I__6670 (
            .O(N__33788),
            .I(N__33785));
    LocalMux I__6669 (
            .O(N__33785),
            .I(N__33782));
    Odrv4 I__6668 (
            .O(N__33782),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ));
    InMux I__6667 (
            .O(N__33779),
            .I(N__33776));
    LocalMux I__6666 (
            .O(N__33776),
            .I(N__33773));
    Span4Mux_h I__6665 (
            .O(N__33773),
            .I(N__33768));
    InMux I__6664 (
            .O(N__33772),
            .I(N__33765));
    InMux I__6663 (
            .O(N__33771),
            .I(N__33762));
    Span4Mux_v I__6662 (
            .O(N__33768),
            .I(N__33759));
    LocalMux I__6661 (
            .O(N__33765),
            .I(N__33754));
    LocalMux I__6660 (
            .O(N__33762),
            .I(N__33754));
    Span4Mux_h I__6659 (
            .O(N__33759),
            .I(N__33751));
    Span4Mux_v I__6658 (
            .O(N__33754),
            .I(N__33748));
    Odrv4 I__6657 (
            .O(N__33751),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    Odrv4 I__6656 (
            .O(N__33748),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    CEMux I__6655 (
            .O(N__33743),
            .I(N__33719));
    CEMux I__6654 (
            .O(N__33742),
            .I(N__33719));
    CEMux I__6653 (
            .O(N__33741),
            .I(N__33719));
    CEMux I__6652 (
            .O(N__33740),
            .I(N__33719));
    CEMux I__6651 (
            .O(N__33739),
            .I(N__33719));
    CEMux I__6650 (
            .O(N__33738),
            .I(N__33719));
    CEMux I__6649 (
            .O(N__33737),
            .I(N__33719));
    CEMux I__6648 (
            .O(N__33736),
            .I(N__33719));
    GlobalMux I__6647 (
            .O(N__33719),
            .I(N__33716));
    gio2CtrlBuf I__6646 (
            .O(N__33716),
            .I(\current_shift_inst.timer_s1.N_162_i_g ));
    InMux I__6645 (
            .O(N__33713),
            .I(N__33709));
    CascadeMux I__6644 (
            .O(N__33712),
            .I(N__33705));
    LocalMux I__6643 (
            .O(N__33709),
            .I(N__33702));
    InMux I__6642 (
            .O(N__33708),
            .I(N__33699));
    InMux I__6641 (
            .O(N__33705),
            .I(N__33696));
    Span4Mux_h I__6640 (
            .O(N__33702),
            .I(N__33688));
    LocalMux I__6639 (
            .O(N__33699),
            .I(N__33688));
    LocalMux I__6638 (
            .O(N__33696),
            .I(N__33688));
    InMux I__6637 (
            .O(N__33695),
            .I(N__33685));
    Span4Mux_h I__6636 (
            .O(N__33688),
            .I(N__33682));
    LocalMux I__6635 (
            .O(N__33685),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    Odrv4 I__6634 (
            .O(N__33682),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    InMux I__6633 (
            .O(N__33677),
            .I(N__33674));
    LocalMux I__6632 (
            .O(N__33674),
            .I(\current_shift_inst.un4_control_input1_1 ));
    CascadeMux I__6631 (
            .O(N__33671),
            .I(\current_shift_inst.un4_control_input1_1_cascade_ ));
    InMux I__6630 (
            .O(N__33668),
            .I(N__33664));
    InMux I__6629 (
            .O(N__33667),
            .I(N__33661));
    LocalMux I__6628 (
            .O(N__33664),
            .I(N__33658));
    LocalMux I__6627 (
            .O(N__33661),
            .I(N__33655));
    Span4Mux_v I__6626 (
            .O(N__33658),
            .I(N__33650));
    Span4Mux_v I__6625 (
            .O(N__33655),
            .I(N__33650));
    Span4Mux_h I__6624 (
            .O(N__33650),
            .I(N__33645));
    InMux I__6623 (
            .O(N__33649),
            .I(N__33642));
    InMux I__6622 (
            .O(N__33648),
            .I(N__33639));
    Odrv4 I__6621 (
            .O(N__33645),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__6620 (
            .O(N__33642),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__6619 (
            .O(N__33639),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    CascadeMux I__6618 (
            .O(N__33632),
            .I(N__33629));
    InMux I__6617 (
            .O(N__33629),
            .I(N__33626));
    LocalMux I__6616 (
            .O(N__33626),
            .I(N__33623));
    Span4Mux_v I__6615 (
            .O(N__33623),
            .I(N__33620));
    Odrv4 I__6614 (
            .O(N__33620),
            .I(\current_shift_inst.un38_control_input_cry_0_s0_sf ));
    CascadeMux I__6613 (
            .O(N__33617),
            .I(N__33612));
    CascadeMux I__6612 (
            .O(N__33616),
            .I(N__33597));
    InMux I__6611 (
            .O(N__33615),
            .I(N__33582));
    InMux I__6610 (
            .O(N__33612),
            .I(N__33582));
    InMux I__6609 (
            .O(N__33611),
            .I(N__33582));
    InMux I__6608 (
            .O(N__33610),
            .I(N__33573));
    InMux I__6607 (
            .O(N__33609),
            .I(N__33573));
    InMux I__6606 (
            .O(N__33608),
            .I(N__33573));
    InMux I__6605 (
            .O(N__33607),
            .I(N__33573));
    InMux I__6604 (
            .O(N__33606),
            .I(N__33562));
    InMux I__6603 (
            .O(N__33605),
            .I(N__33562));
    InMux I__6602 (
            .O(N__33604),
            .I(N__33542));
    InMux I__6601 (
            .O(N__33603),
            .I(N__33542));
    InMux I__6600 (
            .O(N__33602),
            .I(N__33529));
    InMux I__6599 (
            .O(N__33601),
            .I(N__33529));
    InMux I__6598 (
            .O(N__33600),
            .I(N__33529));
    InMux I__6597 (
            .O(N__33597),
            .I(N__33529));
    InMux I__6596 (
            .O(N__33596),
            .I(N__33529));
    InMux I__6595 (
            .O(N__33595),
            .I(N__33529));
    InMux I__6594 (
            .O(N__33594),
            .I(N__33518));
    InMux I__6593 (
            .O(N__33593),
            .I(N__33518));
    InMux I__6592 (
            .O(N__33592),
            .I(N__33518));
    InMux I__6591 (
            .O(N__33591),
            .I(N__33518));
    InMux I__6590 (
            .O(N__33590),
            .I(N__33518));
    InMux I__6589 (
            .O(N__33589),
            .I(N__33512));
    LocalMux I__6588 (
            .O(N__33582),
            .I(N__33509));
    LocalMux I__6587 (
            .O(N__33573),
            .I(N__33506));
    InMux I__6586 (
            .O(N__33572),
            .I(N__33493));
    InMux I__6585 (
            .O(N__33571),
            .I(N__33493));
    InMux I__6584 (
            .O(N__33570),
            .I(N__33493));
    InMux I__6583 (
            .O(N__33569),
            .I(N__33493));
    InMux I__6582 (
            .O(N__33568),
            .I(N__33493));
    InMux I__6581 (
            .O(N__33567),
            .I(N__33493));
    LocalMux I__6580 (
            .O(N__33562),
            .I(N__33489));
    InMux I__6579 (
            .O(N__33561),
            .I(N__33486));
    InMux I__6578 (
            .O(N__33560),
            .I(N__33471));
    InMux I__6577 (
            .O(N__33559),
            .I(N__33471));
    InMux I__6576 (
            .O(N__33558),
            .I(N__33471));
    InMux I__6575 (
            .O(N__33557),
            .I(N__33471));
    InMux I__6574 (
            .O(N__33556),
            .I(N__33471));
    InMux I__6573 (
            .O(N__33555),
            .I(N__33471));
    InMux I__6572 (
            .O(N__33554),
            .I(N__33471));
    InMux I__6571 (
            .O(N__33553),
            .I(N__33455));
    InMux I__6570 (
            .O(N__33552),
            .I(N__33455));
    InMux I__6569 (
            .O(N__33551),
            .I(N__33455));
    InMux I__6568 (
            .O(N__33550),
            .I(N__33455));
    InMux I__6567 (
            .O(N__33549),
            .I(N__33455));
    InMux I__6566 (
            .O(N__33548),
            .I(N__33447));
    InMux I__6565 (
            .O(N__33547),
            .I(N__33444));
    LocalMux I__6564 (
            .O(N__33542),
            .I(N__33441));
    LocalMux I__6563 (
            .O(N__33529),
            .I(N__33436));
    LocalMux I__6562 (
            .O(N__33518),
            .I(N__33436));
    InMux I__6561 (
            .O(N__33517),
            .I(N__33426));
    InMux I__6560 (
            .O(N__33516),
            .I(N__33426));
    InMux I__6559 (
            .O(N__33515),
            .I(N__33426));
    LocalMux I__6558 (
            .O(N__33512),
            .I(N__33417));
    Span4Mux_v I__6557 (
            .O(N__33509),
            .I(N__33417));
    Span4Mux_v I__6556 (
            .O(N__33506),
            .I(N__33417));
    LocalMux I__6555 (
            .O(N__33493),
            .I(N__33417));
    InMux I__6554 (
            .O(N__33492),
            .I(N__33414));
    Span4Mux_v I__6553 (
            .O(N__33489),
            .I(N__33407));
    LocalMux I__6552 (
            .O(N__33486),
            .I(N__33407));
    LocalMux I__6551 (
            .O(N__33471),
            .I(N__33407));
    InMux I__6550 (
            .O(N__33470),
            .I(N__33389));
    InMux I__6549 (
            .O(N__33469),
            .I(N__33389));
    InMux I__6548 (
            .O(N__33468),
            .I(N__33389));
    InMux I__6547 (
            .O(N__33467),
            .I(N__33389));
    InMux I__6546 (
            .O(N__33466),
            .I(N__33389));
    LocalMux I__6545 (
            .O(N__33455),
            .I(N__33386));
    InMux I__6544 (
            .O(N__33454),
            .I(N__33372));
    InMux I__6543 (
            .O(N__33453),
            .I(N__33372));
    InMux I__6542 (
            .O(N__33452),
            .I(N__33372));
    InMux I__6541 (
            .O(N__33451),
            .I(N__33372));
    InMux I__6540 (
            .O(N__33450),
            .I(N__33372));
    LocalMux I__6539 (
            .O(N__33447),
            .I(N__33367));
    LocalMux I__6538 (
            .O(N__33444),
            .I(N__33367));
    Span4Mux_h I__6537 (
            .O(N__33441),
            .I(N__33364));
    Span4Mux_v I__6536 (
            .O(N__33436),
            .I(N__33361));
    InMux I__6535 (
            .O(N__33435),
            .I(N__33354));
    InMux I__6534 (
            .O(N__33434),
            .I(N__33354));
    InMux I__6533 (
            .O(N__33433),
            .I(N__33354));
    LocalMux I__6532 (
            .O(N__33426),
            .I(N__33349));
    Span4Mux_h I__6531 (
            .O(N__33417),
            .I(N__33349));
    LocalMux I__6530 (
            .O(N__33414),
            .I(N__33344));
    Span4Mux_v I__6529 (
            .O(N__33407),
            .I(N__33344));
    InMux I__6528 (
            .O(N__33406),
            .I(N__33329));
    InMux I__6527 (
            .O(N__33405),
            .I(N__33329));
    InMux I__6526 (
            .O(N__33404),
            .I(N__33329));
    InMux I__6525 (
            .O(N__33403),
            .I(N__33329));
    InMux I__6524 (
            .O(N__33402),
            .I(N__33329));
    InMux I__6523 (
            .O(N__33401),
            .I(N__33329));
    InMux I__6522 (
            .O(N__33400),
            .I(N__33329));
    LocalMux I__6521 (
            .O(N__33389),
            .I(N__33324));
    Span4Mux_h I__6520 (
            .O(N__33386),
            .I(N__33324));
    InMux I__6519 (
            .O(N__33385),
            .I(N__33317));
    InMux I__6518 (
            .O(N__33384),
            .I(N__33317));
    InMux I__6517 (
            .O(N__33383),
            .I(N__33317));
    LocalMux I__6516 (
            .O(N__33372),
            .I(N__33310));
    Span4Mux_h I__6515 (
            .O(N__33367),
            .I(N__33310));
    Span4Mux_v I__6514 (
            .O(N__33364),
            .I(N__33310));
    Odrv4 I__6513 (
            .O(N__33361),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__6512 (
            .O(N__33354),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__6511 (
            .O(N__33349),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__6510 (
            .O(N__33344),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__6509 (
            .O(N__33329),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__6508 (
            .O(N__33324),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__6507 (
            .O(N__33317),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__6506 (
            .O(N__33310),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    CascadeMux I__6505 (
            .O(N__33293),
            .I(N__33282));
    InMux I__6504 (
            .O(N__33292),
            .I(N__33255));
    InMux I__6503 (
            .O(N__33291),
            .I(N__33242));
    InMux I__6502 (
            .O(N__33290),
            .I(N__33242));
    InMux I__6501 (
            .O(N__33289),
            .I(N__33242));
    InMux I__6500 (
            .O(N__33288),
            .I(N__33242));
    InMux I__6499 (
            .O(N__33287),
            .I(N__33242));
    InMux I__6498 (
            .O(N__33286),
            .I(N__33242));
    InMux I__6497 (
            .O(N__33285),
            .I(N__33235));
    InMux I__6496 (
            .O(N__33282),
            .I(N__33235));
    InMux I__6495 (
            .O(N__33281),
            .I(N__33235));
    CascadeMux I__6494 (
            .O(N__33280),
            .I(N__33231));
    CascadeMux I__6493 (
            .O(N__33279),
            .I(N__33225));
    CascadeMux I__6492 (
            .O(N__33278),
            .I(N__33215));
    CascadeMux I__6491 (
            .O(N__33277),
            .I(N__33212));
    CascadeMux I__6490 (
            .O(N__33276),
            .I(N__33205));
    CascadeMux I__6489 (
            .O(N__33275),
            .I(N__33202));
    CascadeMux I__6488 (
            .O(N__33274),
            .I(N__33199));
    InMux I__6487 (
            .O(N__33273),
            .I(N__33194));
    InMux I__6486 (
            .O(N__33272),
            .I(N__33194));
    CascadeMux I__6485 (
            .O(N__33271),
            .I(N__33188));
    CascadeMux I__6484 (
            .O(N__33270),
            .I(N__33181));
    CascadeMux I__6483 (
            .O(N__33269),
            .I(N__33176));
    CascadeMux I__6482 (
            .O(N__33268),
            .I(N__33173));
    CascadeMux I__6481 (
            .O(N__33267),
            .I(N__33170));
    CascadeMux I__6480 (
            .O(N__33266),
            .I(N__33162));
    CascadeMux I__6479 (
            .O(N__33265),
            .I(N__33157));
    CascadeMux I__6478 (
            .O(N__33264),
            .I(N__33153));
    CascadeMux I__6477 (
            .O(N__33263),
            .I(N__33149));
    CascadeMux I__6476 (
            .O(N__33262),
            .I(N__33144));
    CascadeMux I__6475 (
            .O(N__33261),
            .I(N__33140));
    CascadeMux I__6474 (
            .O(N__33260),
            .I(N__33136));
    CascadeMux I__6473 (
            .O(N__33259),
            .I(N__33132));
    CascadeMux I__6472 (
            .O(N__33258),
            .I(N__33115));
    LocalMux I__6471 (
            .O(N__33255),
            .I(N__33111));
    LocalMux I__6470 (
            .O(N__33242),
            .I(N__33106));
    LocalMux I__6469 (
            .O(N__33235),
            .I(N__33106));
    InMux I__6468 (
            .O(N__33234),
            .I(N__33103));
    InMux I__6467 (
            .O(N__33231),
            .I(N__33092));
    InMux I__6466 (
            .O(N__33230),
            .I(N__33092));
    InMux I__6465 (
            .O(N__33229),
            .I(N__33092));
    InMux I__6464 (
            .O(N__33228),
            .I(N__33092));
    InMux I__6463 (
            .O(N__33225),
            .I(N__33092));
    InMux I__6462 (
            .O(N__33224),
            .I(N__33087));
    InMux I__6461 (
            .O(N__33223),
            .I(N__33087));
    CascadeMux I__6460 (
            .O(N__33222),
            .I(N__33083));
    CascadeMux I__6459 (
            .O(N__33221),
            .I(N__33080));
    CascadeMux I__6458 (
            .O(N__33220),
            .I(N__33076));
    CascadeMux I__6457 (
            .O(N__33219),
            .I(N__33072));
    CascadeMux I__6456 (
            .O(N__33218),
            .I(N__33069));
    InMux I__6455 (
            .O(N__33215),
            .I(N__33060));
    InMux I__6454 (
            .O(N__33212),
            .I(N__33060));
    InMux I__6453 (
            .O(N__33211),
            .I(N__33045));
    InMux I__6452 (
            .O(N__33210),
            .I(N__33045));
    InMux I__6451 (
            .O(N__33209),
            .I(N__33045));
    InMux I__6450 (
            .O(N__33208),
            .I(N__33045));
    InMux I__6449 (
            .O(N__33205),
            .I(N__33045));
    InMux I__6448 (
            .O(N__33202),
            .I(N__33045));
    InMux I__6447 (
            .O(N__33199),
            .I(N__33045));
    LocalMux I__6446 (
            .O(N__33194),
            .I(N__33042));
    CascadeMux I__6445 (
            .O(N__33193),
            .I(N__33038));
    CascadeMux I__6444 (
            .O(N__33192),
            .I(N__33034));
    CascadeMux I__6443 (
            .O(N__33191),
            .I(N__33030));
    InMux I__6442 (
            .O(N__33188),
            .I(N__33024));
    InMux I__6441 (
            .O(N__33187),
            .I(N__33024));
    InMux I__6440 (
            .O(N__33186),
            .I(N__33011));
    InMux I__6439 (
            .O(N__33185),
            .I(N__33011));
    InMux I__6438 (
            .O(N__33184),
            .I(N__33011));
    InMux I__6437 (
            .O(N__33181),
            .I(N__33011));
    InMux I__6436 (
            .O(N__33180),
            .I(N__33011));
    InMux I__6435 (
            .O(N__33179),
            .I(N__33011));
    InMux I__6434 (
            .O(N__33176),
            .I(N__33004));
    InMux I__6433 (
            .O(N__33173),
            .I(N__33004));
    InMux I__6432 (
            .O(N__33170),
            .I(N__33004));
    InMux I__6431 (
            .O(N__33169),
            .I(N__32991));
    InMux I__6430 (
            .O(N__33168),
            .I(N__32991));
    InMux I__6429 (
            .O(N__33167),
            .I(N__32991));
    InMux I__6428 (
            .O(N__33166),
            .I(N__32991));
    InMux I__6427 (
            .O(N__33165),
            .I(N__32991));
    InMux I__6426 (
            .O(N__33162),
            .I(N__32991));
    InMux I__6425 (
            .O(N__33161),
            .I(N__32974));
    InMux I__6424 (
            .O(N__33160),
            .I(N__32974));
    InMux I__6423 (
            .O(N__33157),
            .I(N__32974));
    InMux I__6422 (
            .O(N__33156),
            .I(N__32974));
    InMux I__6421 (
            .O(N__33153),
            .I(N__32974));
    InMux I__6420 (
            .O(N__33152),
            .I(N__32974));
    InMux I__6419 (
            .O(N__33149),
            .I(N__32974));
    InMux I__6418 (
            .O(N__33148),
            .I(N__32974));
    InMux I__6417 (
            .O(N__33147),
            .I(N__32957));
    InMux I__6416 (
            .O(N__33144),
            .I(N__32957));
    InMux I__6415 (
            .O(N__33143),
            .I(N__32957));
    InMux I__6414 (
            .O(N__33140),
            .I(N__32957));
    InMux I__6413 (
            .O(N__33139),
            .I(N__32957));
    InMux I__6412 (
            .O(N__33136),
            .I(N__32957));
    InMux I__6411 (
            .O(N__33135),
            .I(N__32957));
    InMux I__6410 (
            .O(N__33132),
            .I(N__32957));
    CascadeMux I__6409 (
            .O(N__33131),
            .I(N__32954));
    CascadeMux I__6408 (
            .O(N__33130),
            .I(N__32950));
    CascadeMux I__6407 (
            .O(N__33129),
            .I(N__32946));
    CascadeMux I__6406 (
            .O(N__33128),
            .I(N__32942));
    CascadeMux I__6405 (
            .O(N__33127),
            .I(N__32937));
    CascadeMux I__6404 (
            .O(N__33126),
            .I(N__32933));
    CascadeMux I__6403 (
            .O(N__33125),
            .I(N__32929));
    CascadeMux I__6402 (
            .O(N__33124),
            .I(N__32925));
    CascadeMux I__6401 (
            .O(N__33123),
            .I(N__32921));
    CascadeMux I__6400 (
            .O(N__33122),
            .I(N__32917));
    CascadeMux I__6399 (
            .O(N__33121),
            .I(N__32913));
    InMux I__6398 (
            .O(N__33120),
            .I(N__32899));
    InMux I__6397 (
            .O(N__33119),
            .I(N__32899));
    InMux I__6396 (
            .O(N__33118),
            .I(N__32899));
    InMux I__6395 (
            .O(N__33115),
            .I(N__32899));
    InMux I__6394 (
            .O(N__33114),
            .I(N__32899));
    Span4Mux_v I__6393 (
            .O(N__33111),
            .I(N__32892));
    Span4Mux_v I__6392 (
            .O(N__33106),
            .I(N__32892));
    LocalMux I__6391 (
            .O(N__33103),
            .I(N__32892));
    LocalMux I__6390 (
            .O(N__33092),
            .I(N__32889));
    LocalMux I__6389 (
            .O(N__33087),
            .I(N__32886));
    InMux I__6388 (
            .O(N__33086),
            .I(N__32883));
    InMux I__6387 (
            .O(N__33083),
            .I(N__32878));
    InMux I__6386 (
            .O(N__33080),
            .I(N__32878));
    InMux I__6385 (
            .O(N__33079),
            .I(N__32867));
    InMux I__6384 (
            .O(N__33076),
            .I(N__32867));
    InMux I__6383 (
            .O(N__33075),
            .I(N__32867));
    InMux I__6382 (
            .O(N__33072),
            .I(N__32867));
    InMux I__6381 (
            .O(N__33069),
            .I(N__32867));
    CascadeMux I__6380 (
            .O(N__33068),
            .I(N__32864));
    CascadeMux I__6379 (
            .O(N__33067),
            .I(N__32860));
    CascadeMux I__6378 (
            .O(N__33066),
            .I(N__32856));
    CascadeMux I__6377 (
            .O(N__33065),
            .I(N__32852));
    LocalMux I__6376 (
            .O(N__33060),
            .I(N__32848));
    LocalMux I__6375 (
            .O(N__33045),
            .I(N__32843));
    Span4Mux_v I__6374 (
            .O(N__33042),
            .I(N__32843));
    InMux I__6373 (
            .O(N__33041),
            .I(N__32828));
    InMux I__6372 (
            .O(N__33038),
            .I(N__32828));
    InMux I__6371 (
            .O(N__33037),
            .I(N__32828));
    InMux I__6370 (
            .O(N__33034),
            .I(N__32828));
    InMux I__6369 (
            .O(N__33033),
            .I(N__32828));
    InMux I__6368 (
            .O(N__33030),
            .I(N__32828));
    InMux I__6367 (
            .O(N__33029),
            .I(N__32828));
    LocalMux I__6366 (
            .O(N__33024),
            .I(N__32815));
    LocalMux I__6365 (
            .O(N__33011),
            .I(N__32815));
    LocalMux I__6364 (
            .O(N__33004),
            .I(N__32815));
    LocalMux I__6363 (
            .O(N__32991),
            .I(N__32815));
    LocalMux I__6362 (
            .O(N__32974),
            .I(N__32815));
    LocalMux I__6361 (
            .O(N__32957),
            .I(N__32815));
    InMux I__6360 (
            .O(N__32954),
            .I(N__32798));
    InMux I__6359 (
            .O(N__32953),
            .I(N__32798));
    InMux I__6358 (
            .O(N__32950),
            .I(N__32798));
    InMux I__6357 (
            .O(N__32949),
            .I(N__32798));
    InMux I__6356 (
            .O(N__32946),
            .I(N__32798));
    InMux I__6355 (
            .O(N__32945),
            .I(N__32798));
    InMux I__6354 (
            .O(N__32942),
            .I(N__32798));
    InMux I__6353 (
            .O(N__32941),
            .I(N__32798));
    InMux I__6352 (
            .O(N__32940),
            .I(N__32781));
    InMux I__6351 (
            .O(N__32937),
            .I(N__32781));
    InMux I__6350 (
            .O(N__32936),
            .I(N__32781));
    InMux I__6349 (
            .O(N__32933),
            .I(N__32781));
    InMux I__6348 (
            .O(N__32932),
            .I(N__32781));
    InMux I__6347 (
            .O(N__32929),
            .I(N__32781));
    InMux I__6346 (
            .O(N__32928),
            .I(N__32781));
    InMux I__6345 (
            .O(N__32925),
            .I(N__32781));
    InMux I__6344 (
            .O(N__32924),
            .I(N__32768));
    InMux I__6343 (
            .O(N__32921),
            .I(N__32768));
    InMux I__6342 (
            .O(N__32920),
            .I(N__32768));
    InMux I__6341 (
            .O(N__32917),
            .I(N__32768));
    InMux I__6340 (
            .O(N__32916),
            .I(N__32768));
    InMux I__6339 (
            .O(N__32913),
            .I(N__32768));
    CascadeMux I__6338 (
            .O(N__32912),
            .I(N__32765));
    CascadeMux I__6337 (
            .O(N__32911),
            .I(N__32761));
    CascadeMux I__6336 (
            .O(N__32910),
            .I(N__32757));
    LocalMux I__6335 (
            .O(N__32899),
            .I(N__32753));
    Span4Mux_v I__6334 (
            .O(N__32892),
            .I(N__32750));
    Span4Mux_h I__6333 (
            .O(N__32889),
            .I(N__32747));
    Span4Mux_v I__6332 (
            .O(N__32886),
            .I(N__32738));
    LocalMux I__6331 (
            .O(N__32883),
            .I(N__32738));
    LocalMux I__6330 (
            .O(N__32878),
            .I(N__32738));
    LocalMux I__6329 (
            .O(N__32867),
            .I(N__32738));
    InMux I__6328 (
            .O(N__32864),
            .I(N__32721));
    InMux I__6327 (
            .O(N__32863),
            .I(N__32721));
    InMux I__6326 (
            .O(N__32860),
            .I(N__32721));
    InMux I__6325 (
            .O(N__32859),
            .I(N__32721));
    InMux I__6324 (
            .O(N__32856),
            .I(N__32721));
    InMux I__6323 (
            .O(N__32855),
            .I(N__32721));
    InMux I__6322 (
            .O(N__32852),
            .I(N__32721));
    InMux I__6321 (
            .O(N__32851),
            .I(N__32721));
    Span4Mux_h I__6320 (
            .O(N__32848),
            .I(N__32706));
    Span4Mux_h I__6319 (
            .O(N__32843),
            .I(N__32706));
    LocalMux I__6318 (
            .O(N__32828),
            .I(N__32706));
    Span4Mux_v I__6317 (
            .O(N__32815),
            .I(N__32706));
    LocalMux I__6316 (
            .O(N__32798),
            .I(N__32706));
    LocalMux I__6315 (
            .O(N__32781),
            .I(N__32706));
    LocalMux I__6314 (
            .O(N__32768),
            .I(N__32706));
    InMux I__6313 (
            .O(N__32765),
            .I(N__32693));
    InMux I__6312 (
            .O(N__32764),
            .I(N__32693));
    InMux I__6311 (
            .O(N__32761),
            .I(N__32693));
    InMux I__6310 (
            .O(N__32760),
            .I(N__32693));
    InMux I__6309 (
            .O(N__32757),
            .I(N__32693));
    InMux I__6308 (
            .O(N__32756),
            .I(N__32693));
    Odrv12 I__6307 (
            .O(N__32753),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__6306 (
            .O(N__32750),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__6305 (
            .O(N__32747),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__6304 (
            .O(N__32738),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__6303 (
            .O(N__32721),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__6302 (
            .O(N__32706),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__6301 (
            .O(N__32693),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    CascadeMux I__6300 (
            .O(N__32678),
            .I(N__32675));
    InMux I__6299 (
            .O(N__32675),
            .I(N__32671));
    InMux I__6298 (
            .O(N__32674),
            .I(N__32668));
    LocalMux I__6297 (
            .O(N__32671),
            .I(N__32662));
    LocalMux I__6296 (
            .O(N__32668),
            .I(N__32662));
    InMux I__6295 (
            .O(N__32667),
            .I(N__32659));
    Span4Mux_h I__6294 (
            .O(N__32662),
            .I(N__32656));
    LocalMux I__6293 (
            .O(N__32659),
            .I(N__32653));
    Span4Mux_h I__6292 (
            .O(N__32656),
            .I(N__32649));
    Span4Mux_h I__6291 (
            .O(N__32653),
            .I(N__32646));
    InMux I__6290 (
            .O(N__32652),
            .I(N__32643));
    Odrv4 I__6289 (
            .O(N__32649),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    Odrv4 I__6288 (
            .O(N__32646),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    LocalMux I__6287 (
            .O(N__32643),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    InMux I__6286 (
            .O(N__32636),
            .I(N__32633));
    LocalMux I__6285 (
            .O(N__32633),
            .I(N__32629));
    InMux I__6284 (
            .O(N__32632),
            .I(N__32626));
    Span4Mux_h I__6283 (
            .O(N__32629),
            .I(N__32620));
    LocalMux I__6282 (
            .O(N__32626),
            .I(N__32620));
    InMux I__6281 (
            .O(N__32625),
            .I(N__32617));
    Odrv4 I__6280 (
            .O(N__32620),
            .I(\current_shift_inst.un4_control_input1_3 ));
    LocalMux I__6279 (
            .O(N__32617),
            .I(\current_shift_inst.un4_control_input1_3 ));
    InMux I__6278 (
            .O(N__32612),
            .I(N__32609));
    LocalMux I__6277 (
            .O(N__32609),
            .I(N__32606));
    Span4Mux_h I__6276 (
            .O(N__32606),
            .I(N__32603));
    Odrv4 I__6275 (
            .O(N__32603),
            .I(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ));
    IoInMux I__6274 (
            .O(N__32600),
            .I(N__32597));
    LocalMux I__6273 (
            .O(N__32597),
            .I(N__32594));
    Span12Mux_s0_v I__6272 (
            .O(N__32594),
            .I(N__32591));
    Odrv12 I__6271 (
            .O(N__32591),
            .I(\current_shift_inst.timer_s1.N_162_i ));
    CEMux I__6270 (
            .O(N__32588),
            .I(N__32585));
    LocalMux I__6269 (
            .O(N__32585),
            .I(N__32579));
    CEMux I__6268 (
            .O(N__32584),
            .I(N__32576));
    CEMux I__6267 (
            .O(N__32583),
            .I(N__32573));
    CEMux I__6266 (
            .O(N__32582),
            .I(N__32570));
    Span4Mux_v I__6265 (
            .O(N__32579),
            .I(N__32565));
    LocalMux I__6264 (
            .O(N__32576),
            .I(N__32565));
    LocalMux I__6263 (
            .O(N__32573),
            .I(N__32562));
    LocalMux I__6262 (
            .O(N__32570),
            .I(N__32559));
    Span4Mux_v I__6261 (
            .O(N__32565),
            .I(N__32556));
    Span4Mux_h I__6260 (
            .O(N__32562),
            .I(N__32551));
    Span4Mux_v I__6259 (
            .O(N__32559),
            .I(N__32551));
    Sp12to4 I__6258 (
            .O(N__32556),
            .I(N__32548));
    Span4Mux_h I__6257 (
            .O(N__32551),
            .I(N__32545));
    Odrv12 I__6256 (
            .O(N__32548),
            .I(\current_shift_inst.timer_s1.N_163_i ));
    Odrv4 I__6255 (
            .O(N__32545),
            .I(\current_shift_inst.timer_s1.N_163_i ));
    CascadeMux I__6254 (
            .O(N__32540),
            .I(N__32537));
    InMux I__6253 (
            .O(N__32537),
            .I(N__32534));
    LocalMux I__6252 (
            .O(N__32534),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ));
    CascadeMux I__6251 (
            .O(N__32531),
            .I(N__32528));
    InMux I__6250 (
            .O(N__32528),
            .I(N__32525));
    LocalMux I__6249 (
            .O(N__32525),
            .I(\current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ));
    InMux I__6248 (
            .O(N__32522),
            .I(N__32519));
    LocalMux I__6247 (
            .O(N__32519),
            .I(\current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ));
    InMux I__6246 (
            .O(N__32516),
            .I(N__32512));
    InMux I__6245 (
            .O(N__32515),
            .I(N__32509));
    LocalMux I__6244 (
            .O(N__32512),
            .I(N__32506));
    LocalMux I__6243 (
            .O(N__32509),
            .I(N__32503));
    Span4Mux_v I__6242 (
            .O(N__32506),
            .I(N__32500));
    Span4Mux_h I__6241 (
            .O(N__32503),
            .I(N__32496));
    Span4Mux_h I__6240 (
            .O(N__32500),
            .I(N__32493));
    InMux I__6239 (
            .O(N__32499),
            .I(N__32490));
    Odrv4 I__6238 (
            .O(N__32496),
            .I(\current_shift_inst.un4_control_input1_18 ));
    Odrv4 I__6237 (
            .O(N__32493),
            .I(\current_shift_inst.un4_control_input1_18 ));
    LocalMux I__6236 (
            .O(N__32490),
            .I(\current_shift_inst.un4_control_input1_18 ));
    CascadeMux I__6235 (
            .O(N__32483),
            .I(N__32479));
    CascadeMux I__6234 (
            .O(N__32482),
            .I(N__32476));
    InMux I__6233 (
            .O(N__32479),
            .I(N__32473));
    InMux I__6232 (
            .O(N__32476),
            .I(N__32470));
    LocalMux I__6231 (
            .O(N__32473),
            .I(N__32467));
    LocalMux I__6230 (
            .O(N__32470),
            .I(N__32464));
    Span4Mux_v I__6229 (
            .O(N__32467),
            .I(N__32461));
    Span4Mux_h I__6228 (
            .O(N__32464),
            .I(N__32456));
    Span4Mux_v I__6227 (
            .O(N__32461),
            .I(N__32453));
    InMux I__6226 (
            .O(N__32460),
            .I(N__32450));
    InMux I__6225 (
            .O(N__32459),
            .I(N__32447));
    Span4Mux_h I__6224 (
            .O(N__32456),
            .I(N__32444));
    Sp12to4 I__6223 (
            .O(N__32453),
            .I(N__32437));
    LocalMux I__6222 (
            .O(N__32450),
            .I(N__32437));
    LocalMux I__6221 (
            .O(N__32447),
            .I(N__32437));
    Odrv4 I__6220 (
            .O(N__32444),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    Odrv12 I__6219 (
            .O(N__32437),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    InMux I__6218 (
            .O(N__32432),
            .I(N__32429));
    LocalMux I__6217 (
            .O(N__32429),
            .I(\current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ));
    InMux I__6216 (
            .O(N__32426),
            .I(N__32423));
    LocalMux I__6215 (
            .O(N__32423),
            .I(N__32419));
    InMux I__6214 (
            .O(N__32422),
            .I(N__32415));
    Span4Mux_v I__6213 (
            .O(N__32419),
            .I(N__32412));
    InMux I__6212 (
            .O(N__32418),
            .I(N__32409));
    LocalMux I__6211 (
            .O(N__32415),
            .I(N__32406));
    Span4Mux_h I__6210 (
            .O(N__32412),
            .I(N__32401));
    LocalMux I__6209 (
            .O(N__32409),
            .I(N__32401));
    Span12Mux_v I__6208 (
            .O(N__32406),
            .I(N__32397));
    Span4Mux_v I__6207 (
            .O(N__32401),
            .I(N__32394));
    InMux I__6206 (
            .O(N__32400),
            .I(N__32391));
    Odrv12 I__6205 (
            .O(N__32397),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    Odrv4 I__6204 (
            .O(N__32394),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    LocalMux I__6203 (
            .O(N__32391),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    CascadeMux I__6202 (
            .O(N__32384),
            .I(N__32381));
    InMux I__6201 (
            .O(N__32381),
            .I(N__32378));
    LocalMux I__6200 (
            .O(N__32378),
            .I(N__32375));
    Span4Mux_v I__6199 (
            .O(N__32375),
            .I(N__32371));
    InMux I__6198 (
            .O(N__32374),
            .I(N__32368));
    Span4Mux_h I__6197 (
            .O(N__32371),
            .I(N__32363));
    LocalMux I__6196 (
            .O(N__32368),
            .I(N__32363));
    Span4Mux_h I__6195 (
            .O(N__32363),
            .I(N__32359));
    InMux I__6194 (
            .O(N__32362),
            .I(N__32356));
    Odrv4 I__6193 (
            .O(N__32359),
            .I(\current_shift_inst.un4_control_input1_5 ));
    LocalMux I__6192 (
            .O(N__32356),
            .I(\current_shift_inst.un4_control_input1_5 ));
    CascadeMux I__6191 (
            .O(N__32351),
            .I(N__32348));
    InMux I__6190 (
            .O(N__32348),
            .I(N__32345));
    LocalMux I__6189 (
            .O(N__32345),
            .I(N__32342));
    Odrv4 I__6188 (
            .O(N__32342),
            .I(\current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ));
    InMux I__6187 (
            .O(N__32339),
            .I(N__32335));
    InMux I__6186 (
            .O(N__32338),
            .I(N__32332));
    LocalMux I__6185 (
            .O(N__32335),
            .I(N__32329));
    LocalMux I__6184 (
            .O(N__32332),
            .I(N__32325));
    Span4Mux_h I__6183 (
            .O(N__32329),
            .I(N__32322));
    InMux I__6182 (
            .O(N__32328),
            .I(N__32319));
    Span4Mux_h I__6181 (
            .O(N__32325),
            .I(N__32315));
    Span4Mux_v I__6180 (
            .O(N__32322),
            .I(N__32310));
    LocalMux I__6179 (
            .O(N__32319),
            .I(N__32310));
    InMux I__6178 (
            .O(N__32318),
            .I(N__32307));
    Span4Mux_v I__6177 (
            .O(N__32315),
            .I(N__32302));
    Span4Mux_h I__6176 (
            .O(N__32310),
            .I(N__32302));
    LocalMux I__6175 (
            .O(N__32307),
            .I(N__32299));
    Odrv4 I__6174 (
            .O(N__32302),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    Odrv4 I__6173 (
            .O(N__32299),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    InMux I__6172 (
            .O(N__32294),
            .I(N__32291));
    LocalMux I__6171 (
            .O(N__32291),
            .I(N__32287));
    InMux I__6170 (
            .O(N__32290),
            .I(N__32284));
    Span4Mux_h I__6169 (
            .O(N__32287),
            .I(N__32280));
    LocalMux I__6168 (
            .O(N__32284),
            .I(N__32277));
    InMux I__6167 (
            .O(N__32283),
            .I(N__32274));
    Odrv4 I__6166 (
            .O(N__32280),
            .I(\current_shift_inst.un4_control_input1_13 ));
    Odrv4 I__6165 (
            .O(N__32277),
            .I(\current_shift_inst.un4_control_input1_13 ));
    LocalMux I__6164 (
            .O(N__32274),
            .I(\current_shift_inst.un4_control_input1_13 ));
    CascadeMux I__6163 (
            .O(N__32267),
            .I(N__32264));
    InMux I__6162 (
            .O(N__32264),
            .I(N__32261));
    LocalMux I__6161 (
            .O(N__32261),
            .I(N__32258));
    Span4Mux_h I__6160 (
            .O(N__32258),
            .I(N__32255));
    Odrv4 I__6159 (
            .O(N__32255),
            .I(\current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ));
    CascadeMux I__6158 (
            .O(N__32252),
            .I(N__32249));
    InMux I__6157 (
            .O(N__32249),
            .I(N__32245));
    InMux I__6156 (
            .O(N__32248),
            .I(N__32242));
    LocalMux I__6155 (
            .O(N__32245),
            .I(N__32239));
    LocalMux I__6154 (
            .O(N__32242),
            .I(N__32235));
    Span4Mux_h I__6153 (
            .O(N__32239),
            .I(N__32231));
    InMux I__6152 (
            .O(N__32238),
            .I(N__32228));
    Span4Mux_h I__6151 (
            .O(N__32235),
            .I(N__32225));
    InMux I__6150 (
            .O(N__32234),
            .I(N__32222));
    Span4Mux_v I__6149 (
            .O(N__32231),
            .I(N__32219));
    LocalMux I__6148 (
            .O(N__32228),
            .I(N__32216));
    Span4Mux_v I__6147 (
            .O(N__32225),
            .I(N__32211));
    LocalMux I__6146 (
            .O(N__32222),
            .I(N__32211));
    Span4Mux_h I__6145 (
            .O(N__32219),
            .I(N__32208));
    Span4Mux_h I__6144 (
            .O(N__32216),
            .I(N__32205));
    Span4Mux_h I__6143 (
            .O(N__32211),
            .I(N__32202));
    Odrv4 I__6142 (
            .O(N__32208),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    Odrv4 I__6141 (
            .O(N__32205),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    Odrv4 I__6140 (
            .O(N__32202),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    InMux I__6139 (
            .O(N__32195),
            .I(N__32191));
    InMux I__6138 (
            .O(N__32194),
            .I(N__32188));
    LocalMux I__6137 (
            .O(N__32191),
            .I(N__32184));
    LocalMux I__6136 (
            .O(N__32188),
            .I(N__32181));
    InMux I__6135 (
            .O(N__32187),
            .I(N__32178));
    Span4Mux_v I__6134 (
            .O(N__32184),
            .I(N__32175));
    Span4Mux_h I__6133 (
            .O(N__32181),
            .I(N__32170));
    LocalMux I__6132 (
            .O(N__32178),
            .I(N__32170));
    Odrv4 I__6131 (
            .O(N__32175),
            .I(\current_shift_inst.un4_control_input1_15 ));
    Odrv4 I__6130 (
            .O(N__32170),
            .I(\current_shift_inst.un4_control_input1_15 ));
    InMux I__6129 (
            .O(N__32165),
            .I(N__32162));
    LocalMux I__6128 (
            .O(N__32162),
            .I(N__32159));
    Odrv4 I__6127 (
            .O(N__32159),
            .I(\current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ));
    InMux I__6126 (
            .O(N__32156),
            .I(N__32152));
    InMux I__6125 (
            .O(N__32155),
            .I(N__32149));
    LocalMux I__6124 (
            .O(N__32152),
            .I(N__32144));
    LocalMux I__6123 (
            .O(N__32149),
            .I(N__32144));
    Span4Mux_v I__6122 (
            .O(N__32144),
            .I(N__32140));
    InMux I__6121 (
            .O(N__32143),
            .I(N__32136));
    Span4Mux_v I__6120 (
            .O(N__32140),
            .I(N__32133));
    InMux I__6119 (
            .O(N__32139),
            .I(N__32130));
    LocalMux I__6118 (
            .O(N__32136),
            .I(N__32127));
    Span4Mux_h I__6117 (
            .O(N__32133),
            .I(N__32122));
    LocalMux I__6116 (
            .O(N__32130),
            .I(N__32122));
    Odrv12 I__6115 (
            .O(N__32127),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    Odrv4 I__6114 (
            .O(N__32122),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    InMux I__6113 (
            .O(N__32117),
            .I(N__32114));
    LocalMux I__6112 (
            .O(N__32114),
            .I(N__32109));
    InMux I__6111 (
            .O(N__32113),
            .I(N__32106));
    InMux I__6110 (
            .O(N__32112),
            .I(N__32103));
    Span4Mux_h I__6109 (
            .O(N__32109),
            .I(N__32098));
    LocalMux I__6108 (
            .O(N__32106),
            .I(N__32098));
    LocalMux I__6107 (
            .O(N__32103),
            .I(N__32095));
    Span4Mux_v I__6106 (
            .O(N__32098),
            .I(N__32092));
    Span4Mux_h I__6105 (
            .O(N__32095),
            .I(N__32089));
    Odrv4 I__6104 (
            .O(N__32092),
            .I(\current_shift_inst.un4_control_input1_14 ));
    Odrv4 I__6103 (
            .O(N__32089),
            .I(\current_shift_inst.un4_control_input1_14 ));
    CascadeMux I__6102 (
            .O(N__32084),
            .I(N__32081));
    InMux I__6101 (
            .O(N__32081),
            .I(N__32078));
    LocalMux I__6100 (
            .O(N__32078),
            .I(N__32075));
    Odrv4 I__6099 (
            .O(N__32075),
            .I(\current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ));
    InMux I__6098 (
            .O(N__32072),
            .I(N__32069));
    LocalMux I__6097 (
            .O(N__32069),
            .I(N__32066));
    Span4Mux_h I__6096 (
            .O(N__32066),
            .I(N__32063));
    Sp12to4 I__6095 (
            .O(N__32063),
            .I(N__32060));
    Span12Mux_v I__6094 (
            .O(N__32060),
            .I(N__32057));
    Odrv12 I__6093 (
            .O(N__32057),
            .I(il_max_comp1_D1));
    InMux I__6092 (
            .O(N__32054),
            .I(N__32050));
    InMux I__6091 (
            .O(N__32053),
            .I(N__32047));
    LocalMux I__6090 (
            .O(N__32050),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ));
    LocalMux I__6089 (
            .O(N__32047),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ));
    InMux I__6088 (
            .O(N__32042),
            .I(N__32036));
    InMux I__6087 (
            .O(N__32041),
            .I(N__32036));
    LocalMux I__6086 (
            .O(N__32036),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ));
    InMux I__6085 (
            .O(N__32033),
            .I(N__32030));
    LocalMux I__6084 (
            .O(N__32030),
            .I(N__32027));
    Odrv12 I__6083 (
            .O(N__32027),
            .I(\phase_controller_inst2.stoper_tr.un4_running_df30 ));
    InMux I__6082 (
            .O(N__32024),
            .I(N__32015));
    InMux I__6081 (
            .O(N__32023),
            .I(N__32015));
    InMux I__6080 (
            .O(N__32022),
            .I(N__32015));
    LocalMux I__6079 (
            .O(N__32015),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ));
    CascadeMux I__6078 (
            .O(N__32012),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13_cascade_));
    InMux I__6077 (
            .O(N__32009),
            .I(N__32006));
    LocalMux I__6076 (
            .O(N__32006),
            .I(N__32003));
    Span4Mux_h I__6075 (
            .O(N__32003),
            .I(N__32000));
    Span4Mux_v I__6074 (
            .O(N__32000),
            .I(N__31996));
    InMux I__6073 (
            .O(N__31999),
            .I(N__31993));
    Odrv4 I__6072 (
            .O(N__31996),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    LocalMux I__6071 (
            .O(N__31993),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    CascadeMux I__6070 (
            .O(N__31988),
            .I(N__31985));
    InMux I__6069 (
            .O(N__31985),
            .I(N__31979));
    InMux I__6068 (
            .O(N__31984),
            .I(N__31974));
    InMux I__6067 (
            .O(N__31983),
            .I(N__31974));
    InMux I__6066 (
            .O(N__31982),
            .I(N__31971));
    LocalMux I__6065 (
            .O(N__31979),
            .I(N__31968));
    LocalMux I__6064 (
            .O(N__31974),
            .I(N__31965));
    LocalMux I__6063 (
            .O(N__31971),
            .I(N__31962));
    Span4Mux_v I__6062 (
            .O(N__31968),
            .I(N__31959));
    Span4Mux_h I__6061 (
            .O(N__31965),
            .I(N__31955));
    Span12Mux_v I__6060 (
            .O(N__31962),
            .I(N__31952));
    Span4Mux_h I__6059 (
            .O(N__31959),
            .I(N__31949));
    InMux I__6058 (
            .O(N__31958),
            .I(N__31946));
    Span4Mux_h I__6057 (
            .O(N__31955),
            .I(N__31943));
    Odrv12 I__6056 (
            .O(N__31952),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    Odrv4 I__6055 (
            .O(N__31949),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    LocalMux I__6054 (
            .O(N__31946),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    Odrv4 I__6053 (
            .O(N__31943),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    InMux I__6052 (
            .O(N__31934),
            .I(N__31928));
    InMux I__6051 (
            .O(N__31933),
            .I(N__31928));
    LocalMux I__6050 (
            .O(N__31928),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ));
    CascadeMux I__6049 (
            .O(N__31925),
            .I(N__31922));
    InMux I__6048 (
            .O(N__31922),
            .I(N__31918));
    InMux I__6047 (
            .O(N__31921),
            .I(N__31915));
    LocalMux I__6046 (
            .O(N__31918),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ));
    LocalMux I__6045 (
            .O(N__31915),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ));
    InMux I__6044 (
            .O(N__31910),
            .I(N__31907));
    LocalMux I__6043 (
            .O(N__31907),
            .I(N__31903));
    InMux I__6042 (
            .O(N__31906),
            .I(N__31900));
    Odrv4 I__6041 (
            .O(N__31903),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    LocalMux I__6040 (
            .O(N__31900),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    CascadeMux I__6039 (
            .O(N__31895),
            .I(elapsed_time_ns_1_RNI69DN9_0_28_cascade_));
    InMux I__6038 (
            .O(N__31892),
            .I(N__31885));
    InMux I__6037 (
            .O(N__31891),
            .I(N__31885));
    InMux I__6036 (
            .O(N__31890),
            .I(N__31882));
    LocalMux I__6035 (
            .O(N__31885),
            .I(N__31879));
    LocalMux I__6034 (
            .O(N__31882),
            .I(N__31873));
    Span4Mux_v I__6033 (
            .O(N__31879),
            .I(N__31873));
    InMux I__6032 (
            .O(N__31878),
            .I(N__31870));
    Span4Mux_h I__6031 (
            .O(N__31873),
            .I(N__31865));
    LocalMux I__6030 (
            .O(N__31870),
            .I(N__31865));
    Span4Mux_v I__6029 (
            .O(N__31865),
            .I(N__31862));
    Odrv4 I__6028 (
            .O(N__31862),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    InMux I__6027 (
            .O(N__31859),
            .I(N__31856));
    LocalMux I__6026 (
            .O(N__31856),
            .I(N__31853));
    Span4Mux_h I__6025 (
            .O(N__31853),
            .I(N__31849));
    InMux I__6024 (
            .O(N__31852),
            .I(N__31846));
    Odrv4 I__6023 (
            .O(N__31849),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ));
    LocalMux I__6022 (
            .O(N__31846),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ));
    InMux I__6021 (
            .O(N__31841),
            .I(N__31838));
    LocalMux I__6020 (
            .O(N__31838),
            .I(N__31834));
    InMux I__6019 (
            .O(N__31837),
            .I(N__31831));
    Span4Mux_v I__6018 (
            .O(N__31834),
            .I(N__31825));
    LocalMux I__6017 (
            .O(N__31831),
            .I(N__31825));
    InMux I__6016 (
            .O(N__31830),
            .I(N__31822));
    Span4Mux_v I__6015 (
            .O(N__31825),
            .I(N__31819));
    LocalMux I__6014 (
            .O(N__31822),
            .I(N__31816));
    Sp12to4 I__6013 (
            .O(N__31819),
            .I(N__31813));
    Span12Mux_v I__6012 (
            .O(N__31816),
            .I(N__31808));
    Span12Mux_h I__6011 (
            .O(N__31813),
            .I(N__31808));
    Odrv12 I__6010 (
            .O(N__31808),
            .I(il_min_comp2_c));
    InMux I__6009 (
            .O(N__31805),
            .I(N__31802));
    LocalMux I__6008 (
            .O(N__31802),
            .I(N__31796));
    InMux I__6007 (
            .O(N__31801),
            .I(N__31793));
    InMux I__6006 (
            .O(N__31800),
            .I(N__31790));
    InMux I__6005 (
            .O(N__31799),
            .I(N__31787));
    Span4Mux_v I__6004 (
            .O(N__31796),
            .I(N__31784));
    LocalMux I__6003 (
            .O(N__31793),
            .I(N__31781));
    LocalMux I__6002 (
            .O(N__31790),
            .I(\phase_controller_inst2.hc_time_passed ));
    LocalMux I__6001 (
            .O(N__31787),
            .I(\phase_controller_inst2.hc_time_passed ));
    Odrv4 I__6000 (
            .O(N__31784),
            .I(\phase_controller_inst2.hc_time_passed ));
    Odrv12 I__5999 (
            .O(N__31781),
            .I(\phase_controller_inst2.hc_time_passed ));
    CascadeMux I__5998 (
            .O(N__31772),
            .I(N__31769));
    InMux I__5997 (
            .O(N__31769),
            .I(N__31765));
    InMux I__5996 (
            .O(N__31768),
            .I(N__31762));
    LocalMux I__5995 (
            .O(N__31765),
            .I(N__31758));
    LocalMux I__5994 (
            .O(N__31762),
            .I(N__31755));
    CascadeMux I__5993 (
            .O(N__31761),
            .I(N__31752));
    Span4Mux_h I__5992 (
            .O(N__31758),
            .I(N__31749));
    Span4Mux_v I__5991 (
            .O(N__31755),
            .I(N__31746));
    InMux I__5990 (
            .O(N__31752),
            .I(N__31743));
    Span4Mux_v I__5989 (
            .O(N__31749),
            .I(N__31738));
    Span4Mux_h I__5988 (
            .O(N__31746),
            .I(N__31738));
    LocalMux I__5987 (
            .O(N__31743),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    Odrv4 I__5986 (
            .O(N__31738),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    InMux I__5985 (
            .O(N__31733),
            .I(N__31728));
    InMux I__5984 (
            .O(N__31732),
            .I(N__31725));
    InMux I__5983 (
            .O(N__31731),
            .I(N__31722));
    LocalMux I__5982 (
            .O(N__31728),
            .I(N__31719));
    LocalMux I__5981 (
            .O(N__31725),
            .I(N__31716));
    LocalMux I__5980 (
            .O(N__31722),
            .I(N__31712));
    Span4Mux_h I__5979 (
            .O(N__31719),
            .I(N__31709));
    Span12Mux_s4_v I__5978 (
            .O(N__31716),
            .I(N__31706));
    InMux I__5977 (
            .O(N__31715),
            .I(N__31703));
    Span4Mux_h I__5976 (
            .O(N__31712),
            .I(N__31698));
    Span4Mux_v I__5975 (
            .O(N__31709),
            .I(N__31698));
    Span12Mux_v I__5974 (
            .O(N__31706),
            .I(N__31695));
    LocalMux I__5973 (
            .O(N__31703),
            .I(N__31690));
    Span4Mux_v I__5972 (
            .O(N__31698),
            .I(N__31690));
    Odrv12 I__5971 (
            .O(N__31695),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    Odrv4 I__5970 (
            .O(N__31690),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    InMux I__5969 (
            .O(N__31685),
            .I(N__31682));
    LocalMux I__5968 (
            .O(N__31682),
            .I(N__31679));
    Odrv12 I__5967 (
            .O(N__31679),
            .I(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ));
    CascadeMux I__5966 (
            .O(N__31676),
            .I(\phase_controller_inst2.start_timer_tr_RNO_0_0_cascade_ ));
    InMux I__5965 (
            .O(N__31673),
            .I(N__31667));
    InMux I__5964 (
            .O(N__31672),
            .I(N__31667));
    LocalMux I__5963 (
            .O(N__31667),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    CascadeMux I__5962 (
            .O(N__31664),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ));
    CascadeMux I__5961 (
            .O(N__31661),
            .I(N__31656));
    InMux I__5960 (
            .O(N__31660),
            .I(N__31653));
    InMux I__5959 (
            .O(N__31659),
            .I(N__31648));
    InMux I__5958 (
            .O(N__31656),
            .I(N__31648));
    LocalMux I__5957 (
            .O(N__31653),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ));
    LocalMux I__5956 (
            .O(N__31648),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ));
    CascadeMux I__5955 (
            .O(N__31643),
            .I(N__31638));
    InMux I__5954 (
            .O(N__31642),
            .I(N__31635));
    InMux I__5953 (
            .O(N__31641),
            .I(N__31630));
    InMux I__5952 (
            .O(N__31638),
            .I(N__31630));
    LocalMux I__5951 (
            .O(N__31635),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ));
    LocalMux I__5950 (
            .O(N__31630),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ));
    InMux I__5949 (
            .O(N__31625),
            .I(N__31622));
    LocalMux I__5948 (
            .O(N__31622),
            .I(N__31619));
    Span4Mux_h I__5947 (
            .O(N__31619),
            .I(N__31616));
    Odrv4 I__5946 (
            .O(N__31616),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ));
    InMux I__5945 (
            .O(N__31613),
            .I(N__31609));
    InMux I__5944 (
            .O(N__31612),
            .I(N__31605));
    LocalMux I__5943 (
            .O(N__31609),
            .I(N__31602));
    InMux I__5942 (
            .O(N__31608),
            .I(N__31599));
    LocalMux I__5941 (
            .O(N__31605),
            .I(N__31592));
    Span12Mux_h I__5940 (
            .O(N__31602),
            .I(N__31592));
    LocalMux I__5939 (
            .O(N__31599),
            .I(N__31592));
    Odrv12 I__5938 (
            .O(N__31592),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    InMux I__5937 (
            .O(N__31589),
            .I(N__31586));
    LocalMux I__5936 (
            .O(N__31586),
            .I(N__31581));
    InMux I__5935 (
            .O(N__31585),
            .I(N__31578));
    InMux I__5934 (
            .O(N__31584),
            .I(N__31575));
    Span4Mux_v I__5933 (
            .O(N__31581),
            .I(N__31571));
    LocalMux I__5932 (
            .O(N__31578),
            .I(N__31568));
    LocalMux I__5931 (
            .O(N__31575),
            .I(N__31565));
    InMux I__5930 (
            .O(N__31574),
            .I(N__31562));
    Span4Mux_h I__5929 (
            .O(N__31571),
            .I(N__31555));
    Span4Mux_h I__5928 (
            .O(N__31568),
            .I(N__31555));
    Span4Mux_v I__5927 (
            .O(N__31565),
            .I(N__31555));
    LocalMux I__5926 (
            .O(N__31562),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    Odrv4 I__5925 (
            .O(N__31555),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__5924 (
            .O(N__31550),
            .I(N__31544));
    InMux I__5923 (
            .O(N__31549),
            .I(N__31544));
    LocalMux I__5922 (
            .O(N__31544),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ));
    InMux I__5921 (
            .O(N__31541),
            .I(N__31538));
    LocalMux I__5920 (
            .O(N__31538),
            .I(N__31535));
    Span4Mux_h I__5919 (
            .O(N__31535),
            .I(N__31530));
    InMux I__5918 (
            .O(N__31534),
            .I(N__31527));
    InMux I__5917 (
            .O(N__31533),
            .I(N__31524));
    Span4Mux_h I__5916 (
            .O(N__31530),
            .I(N__31521));
    LocalMux I__5915 (
            .O(N__31527),
            .I(N__31518));
    LocalMux I__5914 (
            .O(N__31524),
            .I(elapsed_time_ns_1_RNI03DN9_0_22));
    Odrv4 I__5913 (
            .O(N__31521),
            .I(elapsed_time_ns_1_RNI03DN9_0_22));
    Odrv4 I__5912 (
            .O(N__31518),
            .I(elapsed_time_ns_1_RNI03DN9_0_22));
    InMux I__5911 (
            .O(N__31511),
            .I(N__31507));
    InMux I__5910 (
            .O(N__31510),
            .I(N__31504));
    LocalMux I__5909 (
            .O(N__31507),
            .I(N__31499));
    LocalMux I__5908 (
            .O(N__31504),
            .I(N__31496));
    InMux I__5907 (
            .O(N__31503),
            .I(N__31493));
    InMux I__5906 (
            .O(N__31502),
            .I(N__31490));
    Span4Mux_v I__5905 (
            .O(N__31499),
            .I(N__31487));
    Span4Mux_v I__5904 (
            .O(N__31496),
            .I(N__31482));
    LocalMux I__5903 (
            .O(N__31493),
            .I(N__31482));
    LocalMux I__5902 (
            .O(N__31490),
            .I(N__31479));
    Span4Mux_h I__5901 (
            .O(N__31487),
            .I(N__31476));
    Span4Mux_h I__5900 (
            .O(N__31482),
            .I(N__31471));
    Span4Mux_v I__5899 (
            .O(N__31479),
            .I(N__31471));
    Odrv4 I__5898 (
            .O(N__31476),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    Odrv4 I__5897 (
            .O(N__31471),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    InMux I__5896 (
            .O(N__31466),
            .I(N__31460));
    InMux I__5895 (
            .O(N__31465),
            .I(N__31460));
    LocalMux I__5894 (
            .O(N__31460),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ));
    InMux I__5893 (
            .O(N__31457),
            .I(N__31454));
    LocalMux I__5892 (
            .O(N__31454),
            .I(N__31451));
    Span4Mux_h I__5891 (
            .O(N__31451),
            .I(N__31448));
    Odrv4 I__5890 (
            .O(N__31448),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt20 ));
    InMux I__5889 (
            .O(N__31445),
            .I(N__31440));
    InMux I__5888 (
            .O(N__31444),
            .I(N__31435));
    InMux I__5887 (
            .O(N__31443),
            .I(N__31435));
    LocalMux I__5886 (
            .O(N__31440),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    LocalMux I__5885 (
            .O(N__31435),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    CascadeMux I__5884 (
            .O(N__31430),
            .I(N__31427));
    InMux I__5883 (
            .O(N__31427),
            .I(N__31420));
    InMux I__5882 (
            .O(N__31426),
            .I(N__31420));
    InMux I__5881 (
            .O(N__31425),
            .I(N__31417));
    LocalMux I__5880 (
            .O(N__31420),
            .I(N__31414));
    LocalMux I__5879 (
            .O(N__31417),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ));
    Odrv4 I__5878 (
            .O(N__31414),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ));
    CascadeMux I__5877 (
            .O(N__31409),
            .I(N__31406));
    InMux I__5876 (
            .O(N__31406),
            .I(N__31403));
    LocalMux I__5875 (
            .O(N__31403),
            .I(N__31400));
    Span4Mux_h I__5874 (
            .O(N__31400),
            .I(N__31397));
    Odrv4 I__5873 (
            .O(N__31397),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ));
    CascadeMux I__5872 (
            .O(N__31394),
            .I(N__31391));
    InMux I__5871 (
            .O(N__31391),
            .I(N__31385));
    InMux I__5870 (
            .O(N__31390),
            .I(N__31385));
    LocalMux I__5869 (
            .O(N__31385),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ));
    InMux I__5868 (
            .O(N__31382),
            .I(N__31379));
    LocalMux I__5867 (
            .O(N__31379),
            .I(N__31375));
    InMux I__5866 (
            .O(N__31378),
            .I(N__31371));
    Span12Mux_h I__5865 (
            .O(N__31375),
            .I(N__31368));
    InMux I__5864 (
            .O(N__31374),
            .I(N__31365));
    LocalMux I__5863 (
            .O(N__31371),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    Odrv12 I__5862 (
            .O(N__31368),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    LocalMux I__5861 (
            .O(N__31365),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    InMux I__5860 (
            .O(N__31358),
            .I(N__31353));
    InMux I__5859 (
            .O(N__31357),
            .I(N__31350));
    InMux I__5858 (
            .O(N__31356),
            .I(N__31347));
    LocalMux I__5857 (
            .O(N__31353),
            .I(N__31343));
    LocalMux I__5856 (
            .O(N__31350),
            .I(N__31338));
    LocalMux I__5855 (
            .O(N__31347),
            .I(N__31338));
    CascadeMux I__5854 (
            .O(N__31346),
            .I(N__31335));
    Span4Mux_v I__5853 (
            .O(N__31343),
            .I(N__31332));
    Span4Mux_v I__5852 (
            .O(N__31338),
            .I(N__31329));
    InMux I__5851 (
            .O(N__31335),
            .I(N__31326));
    Span4Mux_h I__5850 (
            .O(N__31332),
            .I(N__31319));
    Span4Mux_v I__5849 (
            .O(N__31329),
            .I(N__31319));
    LocalMux I__5848 (
            .O(N__31326),
            .I(N__31319));
    Span4Mux_v I__5847 (
            .O(N__31319),
            .I(N__31316));
    Odrv4 I__5846 (
            .O(N__31316),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    InMux I__5845 (
            .O(N__31313),
            .I(N__31307));
    InMux I__5844 (
            .O(N__31312),
            .I(N__31307));
    LocalMux I__5843 (
            .O(N__31307),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ));
    InMux I__5842 (
            .O(N__31304),
            .I(N__31299));
    InMux I__5841 (
            .O(N__31303),
            .I(N__31296));
    InMux I__5840 (
            .O(N__31302),
            .I(N__31293));
    LocalMux I__5839 (
            .O(N__31299),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ));
    LocalMux I__5838 (
            .O(N__31296),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ));
    LocalMux I__5837 (
            .O(N__31293),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ));
    CascadeMux I__5836 (
            .O(N__31286),
            .I(N__31282));
    CascadeMux I__5835 (
            .O(N__31285),
            .I(N__31279));
    InMux I__5834 (
            .O(N__31282),
            .I(N__31276));
    InMux I__5833 (
            .O(N__31279),
            .I(N__31273));
    LocalMux I__5832 (
            .O(N__31276),
            .I(N__31270));
    LocalMux I__5831 (
            .O(N__31273),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ));
    Odrv12 I__5830 (
            .O(N__31270),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ));
    InMux I__5829 (
            .O(N__31265),
            .I(N__31260));
    InMux I__5828 (
            .O(N__31264),
            .I(N__31257));
    InMux I__5827 (
            .O(N__31263),
            .I(N__31254));
    LocalMux I__5826 (
            .O(N__31260),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ));
    LocalMux I__5825 (
            .O(N__31257),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ));
    LocalMux I__5824 (
            .O(N__31254),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ));
    CascadeMux I__5823 (
            .O(N__31247),
            .I(N__31244));
    InMux I__5822 (
            .O(N__31244),
            .I(N__31241));
    LocalMux I__5821 (
            .O(N__31241),
            .I(N__31238));
    Odrv12 I__5820 (
            .O(N__31238),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ));
    InMux I__5819 (
            .O(N__31235),
            .I(N__31231));
    InMux I__5818 (
            .O(N__31234),
            .I(N__31228));
    LocalMux I__5817 (
            .O(N__31231),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    LocalMux I__5816 (
            .O(N__31228),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    InMux I__5815 (
            .O(N__31223),
            .I(N__31219));
    InMux I__5814 (
            .O(N__31222),
            .I(N__31215));
    LocalMux I__5813 (
            .O(N__31219),
            .I(N__31212));
    InMux I__5812 (
            .O(N__31218),
            .I(N__31209));
    LocalMux I__5811 (
            .O(N__31215),
            .I(N__31206));
    Span4Mux_h I__5810 (
            .O(N__31212),
            .I(N__31203));
    LocalMux I__5809 (
            .O(N__31209),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__5808 (
            .O(N__31206),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__5807 (
            .O(N__31203),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    CascadeMux I__5806 (
            .O(N__31196),
            .I(N__31192));
    CascadeMux I__5805 (
            .O(N__31195),
            .I(N__31189));
    InMux I__5804 (
            .O(N__31192),
            .I(N__31186));
    InMux I__5803 (
            .O(N__31189),
            .I(N__31183));
    LocalMux I__5802 (
            .O(N__31186),
            .I(N__31180));
    LocalMux I__5801 (
            .O(N__31183),
            .I(N__31177));
    Span4Mux_h I__5800 (
            .O(N__31180),
            .I(N__31174));
    Odrv4 I__5799 (
            .O(N__31177),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    Odrv4 I__5798 (
            .O(N__31174),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    InMux I__5797 (
            .O(N__31169),
            .I(N__31165));
    InMux I__5796 (
            .O(N__31168),
            .I(N__31161));
    LocalMux I__5795 (
            .O(N__31165),
            .I(N__31158));
    InMux I__5794 (
            .O(N__31164),
            .I(N__31155));
    LocalMux I__5793 (
            .O(N__31161),
            .I(N__31152));
    Span4Mux_h I__5792 (
            .O(N__31158),
            .I(N__31149));
    LocalMux I__5791 (
            .O(N__31155),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__5790 (
            .O(N__31152),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__5789 (
            .O(N__31149),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    CascadeMux I__5788 (
            .O(N__31142),
            .I(N__31139));
    InMux I__5787 (
            .O(N__31139),
            .I(N__31136));
    LocalMux I__5786 (
            .O(N__31136),
            .I(N__31133));
    Span4Mux_v I__5785 (
            .O(N__31133),
            .I(N__31130));
    Odrv4 I__5784 (
            .O(N__31130),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt16 ));
    InMux I__5783 (
            .O(N__31127),
            .I(N__31118));
    InMux I__5782 (
            .O(N__31126),
            .I(N__31118));
    InMux I__5781 (
            .O(N__31125),
            .I(N__31118));
    LocalMux I__5780 (
            .O(N__31118),
            .I(\phase_controller_inst2.tr_time_passed ));
    CascadeMux I__5779 (
            .O(N__31115),
            .I(N__31112));
    InMux I__5778 (
            .O(N__31112),
            .I(N__31108));
    InMux I__5777 (
            .O(N__31111),
            .I(N__31105));
    LocalMux I__5776 (
            .O(N__31108),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    LocalMux I__5775 (
            .O(N__31105),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    CascadeMux I__5774 (
            .O(N__31100),
            .I(\phase_controller_inst2.state_RNI9M3OZ0Z_0_cascade_ ));
    InMux I__5773 (
            .O(N__31097),
            .I(N__31094));
    LocalMux I__5772 (
            .O(N__31094),
            .I(N__31091));
    Span4Mux_v I__5771 (
            .O(N__31091),
            .I(N__31088));
    Odrv4 I__5770 (
            .O(N__31088),
            .I(\phase_controller_inst2.start_timer_hc_0_sqmuxa ));
    InMux I__5769 (
            .O(N__31085),
            .I(N__31082));
    LocalMux I__5768 (
            .O(N__31082),
            .I(N__31079));
    Span4Mux_v I__5767 (
            .O(N__31079),
            .I(N__31076));
    Sp12to4 I__5766 (
            .O(N__31076),
            .I(N__31073));
    Span12Mux_h I__5765 (
            .O(N__31073),
            .I(N__31070));
    Span12Mux_v I__5764 (
            .O(N__31070),
            .I(N__31064));
    InMux I__5763 (
            .O(N__31069),
            .I(N__31057));
    InMux I__5762 (
            .O(N__31068),
            .I(N__31057));
    InMux I__5761 (
            .O(N__31067),
            .I(N__31057));
    Odrv12 I__5760 (
            .O(N__31064),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    LocalMux I__5759 (
            .O(N__31057),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    InMux I__5758 (
            .O(N__31052),
            .I(N__31043));
    InMux I__5757 (
            .O(N__31051),
            .I(N__31043));
    InMux I__5756 (
            .O(N__31050),
            .I(N__31043));
    LocalMux I__5755 (
            .O(N__31043),
            .I(N__31040));
    Span4Mux_v I__5754 (
            .O(N__31040),
            .I(N__31037));
    Span4Mux_h I__5753 (
            .O(N__31037),
            .I(N__31034));
    Span4Mux_h I__5752 (
            .O(N__31034),
            .I(N__31031));
    Odrv4 I__5751 (
            .O(N__31031),
            .I(il_max_comp2_c));
    CascadeMux I__5750 (
            .O(N__31028),
            .I(N__31025));
    InMux I__5749 (
            .O(N__31025),
            .I(N__31022));
    LocalMux I__5748 (
            .O(N__31022),
            .I(N__31019));
    Span4Mux_h I__5747 (
            .O(N__31019),
            .I(N__31016));
    Odrv4 I__5746 (
            .O(N__31016),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt22 ));
    CascadeMux I__5745 (
            .O(N__31013),
            .I(N__31010));
    InMux I__5744 (
            .O(N__31010),
            .I(N__31007));
    LocalMux I__5743 (
            .O(N__31007),
            .I(\pwm_generator_inst.un14_counter_1 ));
    CascadeMux I__5742 (
            .O(N__31004),
            .I(N__31001));
    InMux I__5741 (
            .O(N__31001),
            .I(N__30998));
    LocalMux I__5740 (
            .O(N__30998),
            .I(N__30995));
    Odrv4 I__5739 (
            .O(N__30995),
            .I(\pwm_generator_inst.threshold_0 ));
    CascadeMux I__5738 (
            .O(N__30992),
            .I(N__30989));
    InMux I__5737 (
            .O(N__30989),
            .I(N__30986));
    LocalMux I__5736 (
            .O(N__30986),
            .I(\pwm_generator_inst.threshold_2 ));
    CascadeMux I__5735 (
            .O(N__30983),
            .I(N__30980));
    InMux I__5734 (
            .O(N__30980),
            .I(N__30977));
    LocalMux I__5733 (
            .O(N__30977),
            .I(N__30974));
    Odrv4 I__5732 (
            .O(N__30974),
            .I(\pwm_generator_inst.un14_counter_8 ));
    InMux I__5731 (
            .O(N__30971),
            .I(N__30947));
    InMux I__5730 (
            .O(N__30970),
            .I(N__30947));
    InMux I__5729 (
            .O(N__30969),
            .I(N__30940));
    InMux I__5728 (
            .O(N__30968),
            .I(N__30940));
    InMux I__5727 (
            .O(N__30967),
            .I(N__30940));
    InMux I__5726 (
            .O(N__30966),
            .I(N__30922));
    InMux I__5725 (
            .O(N__30965),
            .I(N__30922));
    InMux I__5724 (
            .O(N__30964),
            .I(N__30922));
    InMux I__5723 (
            .O(N__30963),
            .I(N__30922));
    InMux I__5722 (
            .O(N__30962),
            .I(N__30922));
    InMux I__5721 (
            .O(N__30961),
            .I(N__30922));
    InMux I__5720 (
            .O(N__30960),
            .I(N__30922));
    InMux I__5719 (
            .O(N__30959),
            .I(N__30922));
    InMux I__5718 (
            .O(N__30958),
            .I(N__30907));
    InMux I__5717 (
            .O(N__30957),
            .I(N__30907));
    InMux I__5716 (
            .O(N__30956),
            .I(N__30907));
    InMux I__5715 (
            .O(N__30955),
            .I(N__30907));
    InMux I__5714 (
            .O(N__30954),
            .I(N__30907));
    InMux I__5713 (
            .O(N__30953),
            .I(N__30907));
    InMux I__5712 (
            .O(N__30952),
            .I(N__30907));
    LocalMux I__5711 (
            .O(N__30947),
            .I(N__30904));
    LocalMux I__5710 (
            .O(N__30940),
            .I(N__30901));
    CascadeMux I__5709 (
            .O(N__30939),
            .I(N__30892));
    LocalMux I__5708 (
            .O(N__30922),
            .I(N__30886));
    LocalMux I__5707 (
            .O(N__30907),
            .I(N__30886));
    Span4Mux_v I__5706 (
            .O(N__30904),
            .I(N__30881));
    Span4Mux_v I__5705 (
            .O(N__30901),
            .I(N__30881));
    CascadeMux I__5704 (
            .O(N__30900),
            .I(N__30878));
    CascadeMux I__5703 (
            .O(N__30899),
            .I(N__30874));
    CascadeMux I__5702 (
            .O(N__30898),
            .I(N__30871));
    CascadeMux I__5701 (
            .O(N__30897),
            .I(N__30866));
    CascadeMux I__5700 (
            .O(N__30896),
            .I(N__30863));
    CascadeMux I__5699 (
            .O(N__30895),
            .I(N__30860));
    InMux I__5698 (
            .O(N__30892),
            .I(N__30854));
    InMux I__5697 (
            .O(N__30891),
            .I(N__30854));
    Span12Mux_s10_v I__5696 (
            .O(N__30886),
            .I(N__30851));
    Span4Mux_h I__5695 (
            .O(N__30881),
            .I(N__30848));
    InMux I__5694 (
            .O(N__30878),
            .I(N__30845));
    InMux I__5693 (
            .O(N__30877),
            .I(N__30832));
    InMux I__5692 (
            .O(N__30874),
            .I(N__30832));
    InMux I__5691 (
            .O(N__30871),
            .I(N__30832));
    InMux I__5690 (
            .O(N__30870),
            .I(N__30832));
    InMux I__5689 (
            .O(N__30869),
            .I(N__30832));
    InMux I__5688 (
            .O(N__30866),
            .I(N__30832));
    InMux I__5687 (
            .O(N__30863),
            .I(N__30825));
    InMux I__5686 (
            .O(N__30860),
            .I(N__30825));
    InMux I__5685 (
            .O(N__30859),
            .I(N__30825));
    LocalMux I__5684 (
            .O(N__30854),
            .I(N__30820));
    Span12Mux_h I__5683 (
            .O(N__30851),
            .I(N__30820));
    Sp12to4 I__5682 (
            .O(N__30848),
            .I(N__30817));
    LocalMux I__5681 (
            .O(N__30845),
            .I(N_19_1));
    LocalMux I__5680 (
            .O(N__30832),
            .I(N_19_1));
    LocalMux I__5679 (
            .O(N__30825),
            .I(N_19_1));
    Odrv12 I__5678 (
            .O(N__30820),
            .I(N_19_1));
    Odrv12 I__5677 (
            .O(N__30817),
            .I(N_19_1));
    CascadeMux I__5676 (
            .O(N__30806),
            .I(N__30803));
    InMux I__5675 (
            .O(N__30803),
            .I(N__30800));
    LocalMux I__5674 (
            .O(N__30800),
            .I(\pwm_generator_inst.threshold_9 ));
    IoInMux I__5673 (
            .O(N__30797),
            .I(N__30794));
    LocalMux I__5672 (
            .O(N__30794),
            .I(N__30791));
    IoSpan4Mux I__5671 (
            .O(N__30791),
            .I(N__30788));
    Span4Mux_s0_v I__5670 (
            .O(N__30788),
            .I(N__30785));
    Odrv4 I__5669 (
            .O(N__30785),
            .I(\pll_inst.red_c_i ));
    InMux I__5668 (
            .O(N__30782),
            .I(N__30779));
    LocalMux I__5667 (
            .O(N__30779),
            .I(N__30776));
    Span4Mux_v I__5666 (
            .O(N__30776),
            .I(N__30773));
    Odrv4 I__5665 (
            .O(N__30773),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ));
    InMux I__5664 (
            .O(N__30770),
            .I(N__30764));
    CascadeMux I__5663 (
            .O(N__30769),
            .I(N__30761));
    InMux I__5662 (
            .O(N__30768),
            .I(N__30758));
    InMux I__5661 (
            .O(N__30767),
            .I(N__30755));
    LocalMux I__5660 (
            .O(N__30764),
            .I(N__30752));
    InMux I__5659 (
            .O(N__30761),
            .I(N__30749));
    LocalMux I__5658 (
            .O(N__30758),
            .I(N__30746));
    LocalMux I__5657 (
            .O(N__30755),
            .I(N__30741));
    Span4Mux_h I__5656 (
            .O(N__30752),
            .I(N__30741));
    LocalMux I__5655 (
            .O(N__30749),
            .I(N__30738));
    Span12Mux_s11_v I__5654 (
            .O(N__30746),
            .I(N__30735));
    Span4Mux_v I__5653 (
            .O(N__30741),
            .I(N__30730));
    Span4Mux_h I__5652 (
            .O(N__30738),
            .I(N__30730));
    Odrv12 I__5651 (
            .O(N__30735),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    Odrv4 I__5650 (
            .O(N__30730),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    InMux I__5649 (
            .O(N__30725),
            .I(N__30722));
    LocalMux I__5648 (
            .O(N__30722),
            .I(N__30719));
    Span4Mux_h I__5647 (
            .O(N__30719),
            .I(N__30715));
    InMux I__5646 (
            .O(N__30718),
            .I(N__30711));
    Span4Mux_h I__5645 (
            .O(N__30715),
            .I(N__30708));
    InMux I__5644 (
            .O(N__30714),
            .I(N__30705));
    LocalMux I__5643 (
            .O(N__30711),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    Odrv4 I__5642 (
            .O(N__30708),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    LocalMux I__5641 (
            .O(N__30705),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    InMux I__5640 (
            .O(N__30698),
            .I(\pwm_generator_inst.counter_cry_8 ));
    InMux I__5639 (
            .O(N__30695),
            .I(N__30692));
    LocalMux I__5638 (
            .O(N__30692),
            .I(N__30689));
    Span12Mux_s9_v I__5637 (
            .O(N__30689),
            .I(N__30686));
    Span12Mux_h I__5636 (
            .O(N__30686),
            .I(N__30683));
    Odrv12 I__5635 (
            .O(N__30683),
            .I(\pwm_generator_inst.un2_threshold_2_1_16 ));
    InMux I__5634 (
            .O(N__30680),
            .I(N__30676));
    InMux I__5633 (
            .O(N__30679),
            .I(N__30673));
    LocalMux I__5632 (
            .O(N__30676),
            .I(N__30668));
    LocalMux I__5631 (
            .O(N__30673),
            .I(N__30668));
    Span4Mux_h I__5630 (
            .O(N__30668),
            .I(N__30665));
    Span4Mux_h I__5629 (
            .O(N__30665),
            .I(N__30662));
    Span4Mux_h I__5628 (
            .O(N__30662),
            .I(N__30659));
    Odrv4 I__5627 (
            .O(N__30659),
            .I(\pwm_generator_inst.un2_threshold_2_1_15 ));
    CascadeMux I__5626 (
            .O(N__30656),
            .I(N__30653));
    InMux I__5625 (
            .O(N__30653),
            .I(N__30650));
    LocalMux I__5624 (
            .O(N__30650),
            .I(\pwm_generator_inst.threshold_3 ));
    CascadeMux I__5623 (
            .O(N__30647),
            .I(N__30644));
    InMux I__5622 (
            .O(N__30644),
            .I(N__30641));
    LocalMux I__5621 (
            .O(N__30641),
            .I(\pwm_generator_inst.threshold_4 ));
    CascadeMux I__5620 (
            .O(N__30638),
            .I(N__30635));
    InMux I__5619 (
            .O(N__30635),
            .I(N__30632));
    LocalMux I__5618 (
            .O(N__30632),
            .I(\pwm_generator_inst.threshold_5 ));
    CascadeMux I__5617 (
            .O(N__30629),
            .I(N__30626));
    InMux I__5616 (
            .O(N__30626),
            .I(N__30623));
    LocalMux I__5615 (
            .O(N__30623),
            .I(N__30620));
    Odrv4 I__5614 (
            .O(N__30620),
            .I(\pwm_generator_inst.un14_counter_6 ));
    CascadeMux I__5613 (
            .O(N__30617),
            .I(N__30614));
    InMux I__5612 (
            .O(N__30614),
            .I(N__30611));
    LocalMux I__5611 (
            .O(N__30611),
            .I(\pwm_generator_inst.un14_counter_7 ));
    InMux I__5610 (
            .O(N__30608),
            .I(bfn_12_21_0_));
    InMux I__5609 (
            .O(N__30605),
            .I(\pwm_generator_inst.counter_cry_0 ));
    InMux I__5608 (
            .O(N__30602),
            .I(\pwm_generator_inst.counter_cry_1 ));
    InMux I__5607 (
            .O(N__30599),
            .I(\pwm_generator_inst.counter_cry_2 ));
    InMux I__5606 (
            .O(N__30596),
            .I(\pwm_generator_inst.counter_cry_3 ));
    InMux I__5605 (
            .O(N__30593),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__5604 (
            .O(N__30590),
            .I(\pwm_generator_inst.counter_cry_5 ));
    InMux I__5603 (
            .O(N__30587),
            .I(\pwm_generator_inst.counter_cry_6 ));
    InMux I__5602 (
            .O(N__30584),
            .I(bfn_12_22_0_));
    InMux I__5601 (
            .O(N__30581),
            .I(N__30577));
    InMux I__5600 (
            .O(N__30580),
            .I(N__30574));
    LocalMux I__5599 (
            .O(N__30577),
            .I(N__30570));
    LocalMux I__5598 (
            .O(N__30574),
            .I(N__30567));
    InMux I__5597 (
            .O(N__30573),
            .I(N__30564));
    Span4Mux_h I__5596 (
            .O(N__30570),
            .I(N__30561));
    Span4Mux_v I__5595 (
            .O(N__30567),
            .I(N__30556));
    LocalMux I__5594 (
            .O(N__30564),
            .I(N__30556));
    Span4Mux_h I__5593 (
            .O(N__30561),
            .I(N__30552));
    Span4Mux_h I__5592 (
            .O(N__30556),
            .I(N__30549));
    InMux I__5591 (
            .O(N__30555),
            .I(N__30546));
    Odrv4 I__5590 (
            .O(N__30552),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    Odrv4 I__5589 (
            .O(N__30549),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    LocalMux I__5588 (
            .O(N__30546),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    CascadeMux I__5587 (
            .O(N__30539),
            .I(N__30535));
    InMux I__5586 (
            .O(N__30538),
            .I(N__30532));
    InMux I__5585 (
            .O(N__30535),
            .I(N__30529));
    LocalMux I__5584 (
            .O(N__30532),
            .I(N__30526));
    LocalMux I__5583 (
            .O(N__30529),
            .I(N__30522));
    Span4Mux_h I__5582 (
            .O(N__30526),
            .I(N__30519));
    InMux I__5581 (
            .O(N__30525),
            .I(N__30516));
    Odrv4 I__5580 (
            .O(N__30522),
            .I(\current_shift_inst.un4_control_input1_30 ));
    Odrv4 I__5579 (
            .O(N__30519),
            .I(\current_shift_inst.un4_control_input1_30 ));
    LocalMux I__5578 (
            .O(N__30516),
            .I(\current_shift_inst.un4_control_input1_30 ));
    InMux I__5577 (
            .O(N__30509),
            .I(N__30506));
    LocalMux I__5576 (
            .O(N__30506),
            .I(N__30503));
    Odrv4 I__5575 (
            .O(N__30503),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ));
    InMux I__5574 (
            .O(N__30500),
            .I(N__30496));
    InMux I__5573 (
            .O(N__30499),
            .I(N__30492));
    LocalMux I__5572 (
            .O(N__30496),
            .I(N__30488));
    InMux I__5571 (
            .O(N__30495),
            .I(N__30485));
    LocalMux I__5570 (
            .O(N__30492),
            .I(N__30482));
    InMux I__5569 (
            .O(N__30491),
            .I(N__30479));
    Span4Mux_v I__5568 (
            .O(N__30488),
            .I(N__30476));
    LocalMux I__5567 (
            .O(N__30485),
            .I(N__30473));
    Span4Mux_h I__5566 (
            .O(N__30482),
            .I(N__30468));
    LocalMux I__5565 (
            .O(N__30479),
            .I(N__30468));
    Span4Mux_h I__5564 (
            .O(N__30476),
            .I(N__30465));
    Span4Mux_h I__5563 (
            .O(N__30473),
            .I(N__30462));
    Span4Mux_h I__5562 (
            .O(N__30468),
            .I(N__30459));
    Odrv4 I__5561 (
            .O(N__30465),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    Odrv4 I__5560 (
            .O(N__30462),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    Odrv4 I__5559 (
            .O(N__30459),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    InMux I__5558 (
            .O(N__30452),
            .I(N__30447));
    InMux I__5557 (
            .O(N__30451),
            .I(N__30444));
    InMux I__5556 (
            .O(N__30450),
            .I(N__30441));
    LocalMux I__5555 (
            .O(N__30447),
            .I(N__30438));
    LocalMux I__5554 (
            .O(N__30444),
            .I(N__30435));
    LocalMux I__5553 (
            .O(N__30441),
            .I(N__30432));
    Odrv4 I__5552 (
            .O(N__30438),
            .I(\current_shift_inst.un4_control_input1_12 ));
    Odrv4 I__5551 (
            .O(N__30435),
            .I(\current_shift_inst.un4_control_input1_12 ));
    Odrv4 I__5550 (
            .O(N__30432),
            .I(\current_shift_inst.un4_control_input1_12 ));
    InMux I__5549 (
            .O(N__30425),
            .I(N__30422));
    LocalMux I__5548 (
            .O(N__30422),
            .I(N__30419));
    Odrv12 I__5547 (
            .O(N__30419),
            .I(\current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ));
    CascadeMux I__5546 (
            .O(N__30416),
            .I(N__30413));
    InMux I__5545 (
            .O(N__30413),
            .I(N__30409));
    InMux I__5544 (
            .O(N__30412),
            .I(N__30406));
    LocalMux I__5543 (
            .O(N__30409),
            .I(N__30400));
    LocalMux I__5542 (
            .O(N__30406),
            .I(N__30400));
    InMux I__5541 (
            .O(N__30405),
            .I(N__30397));
    Span4Mux_h I__5540 (
            .O(N__30400),
            .I(N__30393));
    LocalMux I__5539 (
            .O(N__30397),
            .I(N__30390));
    InMux I__5538 (
            .O(N__30396),
            .I(N__30387));
    Span4Mux_h I__5537 (
            .O(N__30393),
            .I(N__30384));
    Span4Mux_v I__5536 (
            .O(N__30390),
            .I(N__30379));
    LocalMux I__5535 (
            .O(N__30387),
            .I(N__30379));
    Odrv4 I__5534 (
            .O(N__30384),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    Odrv4 I__5533 (
            .O(N__30379),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    InMux I__5532 (
            .O(N__30374),
            .I(N__30371));
    LocalMux I__5531 (
            .O(N__30371),
            .I(N__30366));
    InMux I__5530 (
            .O(N__30370),
            .I(N__30363));
    InMux I__5529 (
            .O(N__30369),
            .I(N__30360));
    Odrv4 I__5528 (
            .O(N__30366),
            .I(\current_shift_inst.un4_control_input1_11 ));
    LocalMux I__5527 (
            .O(N__30363),
            .I(\current_shift_inst.un4_control_input1_11 ));
    LocalMux I__5526 (
            .O(N__30360),
            .I(\current_shift_inst.un4_control_input1_11 ));
    CascadeMux I__5525 (
            .O(N__30353),
            .I(N__30350));
    InMux I__5524 (
            .O(N__30350),
            .I(N__30347));
    LocalMux I__5523 (
            .O(N__30347),
            .I(N__30344));
    Span4Mux_v I__5522 (
            .O(N__30344),
            .I(N__30341));
    Odrv4 I__5521 (
            .O(N__30341),
            .I(\current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ));
    CascadeMux I__5520 (
            .O(N__30338),
            .I(N__30334));
    CascadeMux I__5519 (
            .O(N__30337),
            .I(N__30331));
    InMux I__5518 (
            .O(N__30334),
            .I(N__30328));
    InMux I__5517 (
            .O(N__30331),
            .I(N__30324));
    LocalMux I__5516 (
            .O(N__30328),
            .I(N__30321));
    InMux I__5515 (
            .O(N__30327),
            .I(N__30318));
    LocalMux I__5514 (
            .O(N__30324),
            .I(\current_shift_inst.un4_control_input1_23 ));
    Odrv4 I__5513 (
            .O(N__30321),
            .I(\current_shift_inst.un4_control_input1_23 ));
    LocalMux I__5512 (
            .O(N__30318),
            .I(\current_shift_inst.un4_control_input1_23 ));
    InMux I__5511 (
            .O(N__30311),
            .I(N__30307));
    InMux I__5510 (
            .O(N__30310),
            .I(N__30304));
    LocalMux I__5509 (
            .O(N__30307),
            .I(N__30300));
    LocalMux I__5508 (
            .O(N__30304),
            .I(N__30297));
    InMux I__5507 (
            .O(N__30303),
            .I(N__30294));
    Span4Mux_v I__5506 (
            .O(N__30300),
            .I(N__30287));
    Span4Mux_h I__5505 (
            .O(N__30297),
            .I(N__30287));
    LocalMux I__5504 (
            .O(N__30294),
            .I(N__30287));
    Span4Mux_h I__5503 (
            .O(N__30287),
            .I(N__30283));
    InMux I__5502 (
            .O(N__30286),
            .I(N__30280));
    Odrv4 I__5501 (
            .O(N__30283),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    LocalMux I__5500 (
            .O(N__30280),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    CascadeMux I__5499 (
            .O(N__30275),
            .I(N__30272));
    InMux I__5498 (
            .O(N__30272),
            .I(N__30269));
    LocalMux I__5497 (
            .O(N__30269),
            .I(N__30266));
    Span4Mux_v I__5496 (
            .O(N__30266),
            .I(N__30263));
    Odrv4 I__5495 (
            .O(N__30263),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ));
    CascadeMux I__5494 (
            .O(N__30260),
            .I(N__30256));
    InMux I__5493 (
            .O(N__30259),
            .I(N__30253));
    InMux I__5492 (
            .O(N__30256),
            .I(N__30250));
    LocalMux I__5491 (
            .O(N__30253),
            .I(N__30246));
    LocalMux I__5490 (
            .O(N__30250),
            .I(N__30243));
    InMux I__5489 (
            .O(N__30249),
            .I(N__30240));
    Span4Mux_v I__5488 (
            .O(N__30246),
            .I(N__30237));
    Span4Mux_h I__5487 (
            .O(N__30243),
            .I(N__30231));
    LocalMux I__5486 (
            .O(N__30240),
            .I(N__30231));
    Span4Mux_v I__5485 (
            .O(N__30237),
            .I(N__30228));
    InMux I__5484 (
            .O(N__30236),
            .I(N__30225));
    Span4Mux_h I__5483 (
            .O(N__30231),
            .I(N__30222));
    Span4Mux_v I__5482 (
            .O(N__30228),
            .I(N__30217));
    LocalMux I__5481 (
            .O(N__30225),
            .I(N__30217));
    Odrv4 I__5480 (
            .O(N__30222),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    Odrv4 I__5479 (
            .O(N__30217),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    InMux I__5478 (
            .O(N__30212),
            .I(N__30209));
    LocalMux I__5477 (
            .O(N__30209),
            .I(N__30206));
    Span4Mux_h I__5476 (
            .O(N__30206),
            .I(N__30203));
    Span4Mux_v I__5475 (
            .O(N__30203),
            .I(N__30199));
    InMux I__5474 (
            .O(N__30202),
            .I(N__30196));
    Span4Mux_v I__5473 (
            .O(N__30199),
            .I(N__30190));
    LocalMux I__5472 (
            .O(N__30196),
            .I(N__30190));
    InMux I__5471 (
            .O(N__30195),
            .I(N__30187));
    Odrv4 I__5470 (
            .O(N__30190),
            .I(\current_shift_inst.un4_control_input1_20 ));
    LocalMux I__5469 (
            .O(N__30187),
            .I(\current_shift_inst.un4_control_input1_20 ));
    InMux I__5468 (
            .O(N__30182),
            .I(N__30179));
    LocalMux I__5467 (
            .O(N__30179),
            .I(N__30176));
    Span4Mux_v I__5466 (
            .O(N__30176),
            .I(N__30173));
    Odrv4 I__5465 (
            .O(N__30173),
            .I(\current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ));
    CascadeMux I__5464 (
            .O(N__30170),
            .I(N__30165));
    InMux I__5463 (
            .O(N__30169),
            .I(N__30160));
    InMux I__5462 (
            .O(N__30168),
            .I(N__30160));
    InMux I__5461 (
            .O(N__30165),
            .I(N__30156));
    LocalMux I__5460 (
            .O(N__30160),
            .I(N__30153));
    InMux I__5459 (
            .O(N__30159),
            .I(N__30150));
    LocalMux I__5458 (
            .O(N__30156),
            .I(N__30147));
    Span4Mux_v I__5457 (
            .O(N__30153),
            .I(N__30142));
    LocalMux I__5456 (
            .O(N__30150),
            .I(N__30142));
    Span12Mux_h I__5455 (
            .O(N__30147),
            .I(N__30139));
    Span4Mux_h I__5454 (
            .O(N__30142),
            .I(N__30136));
    Odrv12 I__5453 (
            .O(N__30139),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    Odrv4 I__5452 (
            .O(N__30136),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    InMux I__5451 (
            .O(N__30131),
            .I(N__30127));
    InMux I__5450 (
            .O(N__30130),
            .I(N__30123));
    LocalMux I__5449 (
            .O(N__30127),
            .I(N__30120));
    InMux I__5448 (
            .O(N__30126),
            .I(N__30117));
    LocalMux I__5447 (
            .O(N__30123),
            .I(\current_shift_inst.un4_control_input1_21 ));
    Odrv4 I__5446 (
            .O(N__30120),
            .I(\current_shift_inst.un4_control_input1_21 ));
    LocalMux I__5445 (
            .O(N__30117),
            .I(\current_shift_inst.un4_control_input1_21 ));
    CascadeMux I__5444 (
            .O(N__30110),
            .I(N__30107));
    InMux I__5443 (
            .O(N__30107),
            .I(N__30104));
    LocalMux I__5442 (
            .O(N__30104),
            .I(N__30101));
    Span4Mux_v I__5441 (
            .O(N__30101),
            .I(N__30098));
    Odrv4 I__5440 (
            .O(N__30098),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ));
    InMux I__5439 (
            .O(N__30095),
            .I(N__30091));
    InMux I__5438 (
            .O(N__30094),
            .I(N__30087));
    LocalMux I__5437 (
            .O(N__30091),
            .I(N__30084));
    InMux I__5436 (
            .O(N__30090),
            .I(N__30081));
    LocalMux I__5435 (
            .O(N__30087),
            .I(\current_shift_inst.un4_control_input1_24 ));
    Odrv4 I__5434 (
            .O(N__30084),
            .I(\current_shift_inst.un4_control_input1_24 ));
    LocalMux I__5433 (
            .O(N__30081),
            .I(\current_shift_inst.un4_control_input1_24 ));
    InMux I__5432 (
            .O(N__30074),
            .I(N__30070));
    CascadeMux I__5431 (
            .O(N__30073),
            .I(N__30066));
    LocalMux I__5430 (
            .O(N__30070),
            .I(N__30063));
    InMux I__5429 (
            .O(N__30069),
            .I(N__30060));
    InMux I__5428 (
            .O(N__30066),
            .I(N__30057));
    Span4Mux_h I__5427 (
            .O(N__30063),
            .I(N__30053));
    LocalMux I__5426 (
            .O(N__30060),
            .I(N__30050));
    LocalMux I__5425 (
            .O(N__30057),
            .I(N__30047));
    InMux I__5424 (
            .O(N__30056),
            .I(N__30044));
    Span4Mux_h I__5423 (
            .O(N__30053),
            .I(N__30041));
    Span4Mux_h I__5422 (
            .O(N__30050),
            .I(N__30038));
    Span4Mux_v I__5421 (
            .O(N__30047),
            .I(N__30033));
    LocalMux I__5420 (
            .O(N__30044),
            .I(N__30033));
    Odrv4 I__5419 (
            .O(N__30041),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv4 I__5418 (
            .O(N__30038),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv4 I__5417 (
            .O(N__30033),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    InMux I__5416 (
            .O(N__30026),
            .I(N__30023));
    LocalMux I__5415 (
            .O(N__30023),
            .I(N__30020));
    Span4Mux_v I__5414 (
            .O(N__30020),
            .I(N__30017));
    Odrv4 I__5413 (
            .O(N__30017),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ));
    CascadeMux I__5412 (
            .O(N__30014),
            .I(N__30011));
    InMux I__5411 (
            .O(N__30011),
            .I(N__30008));
    LocalMux I__5410 (
            .O(N__30008),
            .I(N__30002));
    InMux I__5409 (
            .O(N__30007),
            .I(N__29999));
    InMux I__5408 (
            .O(N__30006),
            .I(N__29996));
    InMux I__5407 (
            .O(N__30005),
            .I(N__29993));
    Span4Mux_v I__5406 (
            .O(N__30002),
            .I(N__29990));
    LocalMux I__5405 (
            .O(N__29999),
            .I(N__29987));
    LocalMux I__5404 (
            .O(N__29996),
            .I(N__29982));
    LocalMux I__5403 (
            .O(N__29993),
            .I(N__29982));
    Span4Mux_h I__5402 (
            .O(N__29990),
            .I(N__29977));
    Span4Mux_v I__5401 (
            .O(N__29987),
            .I(N__29977));
    Span4Mux_v I__5400 (
            .O(N__29982),
            .I(N__29974));
    Odrv4 I__5399 (
            .O(N__29977),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    Odrv4 I__5398 (
            .O(N__29974),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    InMux I__5397 (
            .O(N__29969),
            .I(N__29966));
    LocalMux I__5396 (
            .O(N__29966),
            .I(N__29961));
    InMux I__5395 (
            .O(N__29965),
            .I(N__29958));
    InMux I__5394 (
            .O(N__29964),
            .I(N__29955));
    Odrv4 I__5393 (
            .O(N__29961),
            .I(\current_shift_inst.un4_control_input1_19 ));
    LocalMux I__5392 (
            .O(N__29958),
            .I(\current_shift_inst.un4_control_input1_19 ));
    LocalMux I__5391 (
            .O(N__29955),
            .I(\current_shift_inst.un4_control_input1_19 ));
    CascadeMux I__5390 (
            .O(N__29948),
            .I(N__29945));
    InMux I__5389 (
            .O(N__29945),
            .I(N__29942));
    LocalMux I__5388 (
            .O(N__29942),
            .I(N__29939));
    Span4Mux_v I__5387 (
            .O(N__29939),
            .I(N__29936));
    Odrv4 I__5386 (
            .O(N__29936),
            .I(\current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ));
    CascadeMux I__5385 (
            .O(N__29933),
            .I(N__29930));
    InMux I__5384 (
            .O(N__29930),
            .I(N__29918));
    InMux I__5383 (
            .O(N__29929),
            .I(N__29918));
    InMux I__5382 (
            .O(N__29928),
            .I(N__29918));
    InMux I__5381 (
            .O(N__29927),
            .I(N__29918));
    LocalMux I__5380 (
            .O(N__29918),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    CascadeMux I__5379 (
            .O(N__29915),
            .I(N__29911));
    InMux I__5378 (
            .O(N__29914),
            .I(N__29903));
    InMux I__5377 (
            .O(N__29911),
            .I(N__29903));
    InMux I__5376 (
            .O(N__29910),
            .I(N__29903));
    LocalMux I__5375 (
            .O(N__29903),
            .I(N__29900));
    Span4Mux_v I__5374 (
            .O(N__29900),
            .I(N__29897));
    Span4Mux_h I__5373 (
            .O(N__29897),
            .I(N__29894));
    Span4Mux_h I__5372 (
            .O(N__29894),
            .I(N__29891));
    Odrv4 I__5371 (
            .O(N__29891),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    CEMux I__5370 (
            .O(N__29888),
            .I(N__29883));
    CEMux I__5369 (
            .O(N__29887),
            .I(N__29879));
    CEMux I__5368 (
            .O(N__29886),
            .I(N__29876));
    LocalMux I__5367 (
            .O(N__29883),
            .I(N__29872));
    CEMux I__5366 (
            .O(N__29882),
            .I(N__29869));
    LocalMux I__5365 (
            .O(N__29879),
            .I(N__29866));
    LocalMux I__5364 (
            .O(N__29876),
            .I(N__29863));
    CEMux I__5363 (
            .O(N__29875),
            .I(N__29860));
    Span4Mux_h I__5362 (
            .O(N__29872),
            .I(N__29857));
    LocalMux I__5361 (
            .O(N__29869),
            .I(N__29854));
    Span4Mux_v I__5360 (
            .O(N__29866),
            .I(N__29847));
    Span4Mux_v I__5359 (
            .O(N__29863),
            .I(N__29847));
    LocalMux I__5358 (
            .O(N__29860),
            .I(N__29847));
    Span4Mux_v I__5357 (
            .O(N__29857),
            .I(N__29844));
    Span4Mux_v I__5356 (
            .O(N__29854),
            .I(N__29841));
    Span4Mux_h I__5355 (
            .O(N__29847),
            .I(N__29838));
    Span4Mux_v I__5354 (
            .O(N__29844),
            .I(N__29835));
    Span4Mux_h I__5353 (
            .O(N__29841),
            .I(N__29830));
    Span4Mux_h I__5352 (
            .O(N__29838),
            .I(N__29830));
    Odrv4 I__5351 (
            .O(N__29835),
            .I(\delay_measurement_inst.delay_hc_timer.N_198_i ));
    Odrv4 I__5350 (
            .O(N__29830),
            .I(\delay_measurement_inst.delay_hc_timer.N_198_i ));
    CascadeMux I__5349 (
            .O(N__29825),
            .I(N__29822));
    InMux I__5348 (
            .O(N__29822),
            .I(N__29819));
    LocalMux I__5347 (
            .O(N__29819),
            .I(\current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ));
    CascadeMux I__5346 (
            .O(N__29816),
            .I(N__29812));
    CascadeMux I__5345 (
            .O(N__29815),
            .I(N__29809));
    InMux I__5344 (
            .O(N__29812),
            .I(N__29806));
    InMux I__5343 (
            .O(N__29809),
            .I(N__29803));
    LocalMux I__5342 (
            .O(N__29806),
            .I(N__29799));
    LocalMux I__5341 (
            .O(N__29803),
            .I(N__29796));
    InMux I__5340 (
            .O(N__29802),
            .I(N__29793));
    Span4Mux_v I__5339 (
            .O(N__29799),
            .I(N__29788));
    Span4Mux_h I__5338 (
            .O(N__29796),
            .I(N__29788));
    LocalMux I__5337 (
            .O(N__29793),
            .I(N__29785));
    Span4Mux_h I__5336 (
            .O(N__29788),
            .I(N__29781));
    Span4Mux_h I__5335 (
            .O(N__29785),
            .I(N__29778));
    InMux I__5334 (
            .O(N__29784),
            .I(N__29775));
    Odrv4 I__5333 (
            .O(N__29781),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    Odrv4 I__5332 (
            .O(N__29778),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    LocalMux I__5331 (
            .O(N__29775),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    InMux I__5330 (
            .O(N__29768),
            .I(N__29764));
    InMux I__5329 (
            .O(N__29767),
            .I(N__29761));
    LocalMux I__5328 (
            .O(N__29764),
            .I(N__29757));
    LocalMux I__5327 (
            .O(N__29761),
            .I(N__29754));
    InMux I__5326 (
            .O(N__29760),
            .I(N__29751));
    Odrv4 I__5325 (
            .O(N__29757),
            .I(\current_shift_inst.un4_control_input1_4 ));
    Odrv4 I__5324 (
            .O(N__29754),
            .I(\current_shift_inst.un4_control_input1_4 ));
    LocalMux I__5323 (
            .O(N__29751),
            .I(\current_shift_inst.un4_control_input1_4 ));
    InMux I__5322 (
            .O(N__29744),
            .I(N__29741));
    LocalMux I__5321 (
            .O(N__29741),
            .I(N__29738));
    Odrv12 I__5320 (
            .O(N__29738),
            .I(\current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ));
    CascadeMux I__5319 (
            .O(N__29735),
            .I(N__29732));
    InMux I__5318 (
            .O(N__29732),
            .I(N__29729));
    LocalMux I__5317 (
            .O(N__29729),
            .I(N__29726));
    Span4Mux_v I__5316 (
            .O(N__29726),
            .I(N__29723));
    Odrv4 I__5315 (
            .O(N__29723),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ));
    CascadeMux I__5314 (
            .O(N__29720),
            .I(N__29716));
    InMux I__5313 (
            .O(N__29719),
            .I(N__29713));
    InMux I__5312 (
            .O(N__29716),
            .I(N__29710));
    LocalMux I__5311 (
            .O(N__29713),
            .I(N__29706));
    LocalMux I__5310 (
            .O(N__29710),
            .I(N__29703));
    InMux I__5309 (
            .O(N__29709),
            .I(N__29700));
    Odrv4 I__5308 (
            .O(N__29706),
            .I(\current_shift_inst.un4_control_input1_8 ));
    Odrv4 I__5307 (
            .O(N__29703),
            .I(\current_shift_inst.un4_control_input1_8 ));
    LocalMux I__5306 (
            .O(N__29700),
            .I(\current_shift_inst.un4_control_input1_8 ));
    CascadeMux I__5305 (
            .O(N__29693),
            .I(N__29688));
    InMux I__5304 (
            .O(N__29692),
            .I(N__29685));
    InMux I__5303 (
            .O(N__29691),
            .I(N__29682));
    InMux I__5302 (
            .O(N__29688),
            .I(N__29679));
    LocalMux I__5301 (
            .O(N__29685),
            .I(N__29676));
    LocalMux I__5300 (
            .O(N__29682),
            .I(N__29672));
    LocalMux I__5299 (
            .O(N__29679),
            .I(N__29669));
    Span4Mux_v I__5298 (
            .O(N__29676),
            .I(N__29666));
    InMux I__5297 (
            .O(N__29675),
            .I(N__29663));
    Span4Mux_v I__5296 (
            .O(N__29672),
            .I(N__29660));
    Span4Mux_h I__5295 (
            .O(N__29669),
            .I(N__29653));
    Span4Mux_h I__5294 (
            .O(N__29666),
            .I(N__29653));
    LocalMux I__5293 (
            .O(N__29663),
            .I(N__29653));
    Odrv4 I__5292 (
            .O(N__29660),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    Odrv4 I__5291 (
            .O(N__29653),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    InMux I__5290 (
            .O(N__29648),
            .I(N__29645));
    LocalMux I__5289 (
            .O(N__29645),
            .I(N__29642));
    Span12Mux_v I__5288 (
            .O(N__29642),
            .I(N__29639));
    Odrv12 I__5287 (
            .O(N__29639),
            .I(\current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ));
    CascadeMux I__5286 (
            .O(N__29636),
            .I(N__29632));
    CascadeMux I__5285 (
            .O(N__29635),
            .I(N__29629));
    InMux I__5284 (
            .O(N__29632),
            .I(N__29625));
    InMux I__5283 (
            .O(N__29629),
            .I(N__29622));
    InMux I__5282 (
            .O(N__29628),
            .I(N__29619));
    LocalMux I__5281 (
            .O(N__29625),
            .I(N__29616));
    LocalMux I__5280 (
            .O(N__29622),
            .I(N__29613));
    LocalMux I__5279 (
            .O(N__29619),
            .I(N__29610));
    Span4Mux_h I__5278 (
            .O(N__29616),
            .I(N__29607));
    Span4Mux_h I__5277 (
            .O(N__29613),
            .I(N__29604));
    Span4Mux_h I__5276 (
            .O(N__29610),
            .I(N__29601));
    Span4Mux_v I__5275 (
            .O(N__29607),
            .I(N__29595));
    Span4Mux_h I__5274 (
            .O(N__29604),
            .I(N__29595));
    Span4Mux_v I__5273 (
            .O(N__29601),
            .I(N__29592));
    InMux I__5272 (
            .O(N__29600),
            .I(N__29589));
    Odrv4 I__5271 (
            .O(N__29595),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    Odrv4 I__5270 (
            .O(N__29592),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    LocalMux I__5269 (
            .O(N__29589),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    InMux I__5268 (
            .O(N__29582),
            .I(N__29579));
    LocalMux I__5267 (
            .O(N__29579),
            .I(N__29576));
    Span4Mux_h I__5266 (
            .O(N__29576),
            .I(N__29571));
    InMux I__5265 (
            .O(N__29575),
            .I(N__29568));
    InMux I__5264 (
            .O(N__29574),
            .I(N__29565));
    Span4Mux_v I__5263 (
            .O(N__29571),
            .I(N__29560));
    LocalMux I__5262 (
            .O(N__29568),
            .I(N__29560));
    LocalMux I__5261 (
            .O(N__29565),
            .I(N__29557));
    Odrv4 I__5260 (
            .O(N__29560),
            .I(\current_shift_inst.un4_control_input1_7 ));
    Odrv4 I__5259 (
            .O(N__29557),
            .I(\current_shift_inst.un4_control_input1_7 ));
    CascadeMux I__5258 (
            .O(N__29552),
            .I(N__29549));
    InMux I__5257 (
            .O(N__29549),
            .I(N__29546));
    LocalMux I__5256 (
            .O(N__29546),
            .I(N__29543));
    Sp12to4 I__5255 (
            .O(N__29543),
            .I(N__29540));
    Odrv12 I__5254 (
            .O(N__29540),
            .I(\current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ));
    CascadeMux I__5253 (
            .O(N__29537),
            .I(N__29534));
    InMux I__5252 (
            .O(N__29534),
            .I(N__29529));
    InMux I__5251 (
            .O(N__29533),
            .I(N__29526));
    InMux I__5250 (
            .O(N__29532),
            .I(N__29523));
    LocalMux I__5249 (
            .O(N__29529),
            .I(N__29520));
    LocalMux I__5248 (
            .O(N__29526),
            .I(N__29516));
    LocalMux I__5247 (
            .O(N__29523),
            .I(N__29513));
    Span4Mux_h I__5246 (
            .O(N__29520),
            .I(N__29510));
    InMux I__5245 (
            .O(N__29519),
            .I(N__29507));
    Span4Mux_h I__5244 (
            .O(N__29516),
            .I(N__29504));
    Span4Mux_v I__5243 (
            .O(N__29513),
            .I(N__29501));
    Span4Mux_h I__5242 (
            .O(N__29510),
            .I(N__29496));
    LocalMux I__5241 (
            .O(N__29507),
            .I(N__29496));
    Odrv4 I__5240 (
            .O(N__29504),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    Odrv4 I__5239 (
            .O(N__29501),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    Odrv4 I__5238 (
            .O(N__29496),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    InMux I__5237 (
            .O(N__29489),
            .I(N__29485));
    CascadeMux I__5236 (
            .O(N__29488),
            .I(N__29482));
    LocalMux I__5235 (
            .O(N__29485),
            .I(N__29479));
    InMux I__5234 (
            .O(N__29482),
            .I(N__29475));
    Span4Mux_h I__5233 (
            .O(N__29479),
            .I(N__29472));
    InMux I__5232 (
            .O(N__29478),
            .I(N__29469));
    LocalMux I__5231 (
            .O(N__29475),
            .I(\current_shift_inst.un4_control_input1_17 ));
    Odrv4 I__5230 (
            .O(N__29472),
            .I(\current_shift_inst.un4_control_input1_17 ));
    LocalMux I__5229 (
            .O(N__29469),
            .I(\current_shift_inst.un4_control_input1_17 ));
    CascadeMux I__5228 (
            .O(N__29462),
            .I(N__29459));
    InMux I__5227 (
            .O(N__29459),
            .I(N__29456));
    LocalMux I__5226 (
            .O(N__29456),
            .I(N__29453));
    Span4Mux_h I__5225 (
            .O(N__29453),
            .I(N__29450));
    Odrv4 I__5224 (
            .O(N__29450),
            .I(\current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ));
    CascadeMux I__5223 (
            .O(N__29447),
            .I(N__29443));
    InMux I__5222 (
            .O(N__29446),
            .I(N__29440));
    InMux I__5221 (
            .O(N__29443),
            .I(N__29437));
    LocalMux I__5220 (
            .O(N__29440),
            .I(N__29434));
    LocalMux I__5219 (
            .O(N__29437),
            .I(N__29431));
    Span4Mux_v I__5218 (
            .O(N__29434),
            .I(N__29428));
    Span4Mux_v I__5217 (
            .O(N__29431),
            .I(N__29425));
    Odrv4 I__5216 (
            .O(N__29428),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    Odrv4 I__5215 (
            .O(N__29425),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    InMux I__5214 (
            .O(N__29420),
            .I(\current_shift_inst.un38_control_input_cry_28_s0 ));
    InMux I__5213 (
            .O(N__29417),
            .I(\current_shift_inst.un38_control_input_cry_29_s0 ));
    InMux I__5212 (
            .O(N__29414),
            .I(N__29411));
    LocalMux I__5211 (
            .O(N__29411),
            .I(N__29408));
    Span4Mux_h I__5210 (
            .O(N__29408),
            .I(N__29405));
    Odrv4 I__5209 (
            .O(N__29405),
            .I(\current_shift_inst.un38_control_input_axb_31_s0 ));
    InMux I__5208 (
            .O(N__29402),
            .I(N__29399));
    LocalMux I__5207 (
            .O(N__29399),
            .I(N__29396));
    Odrv4 I__5206 (
            .O(N__29396),
            .I(\current_shift_inst.un38_control_input_0_s1_31 ));
    InMux I__5205 (
            .O(N__29393),
            .I(\current_shift_inst.un38_control_input_cry_30_s0 ));
    InMux I__5204 (
            .O(N__29390),
            .I(N__29387));
    LocalMux I__5203 (
            .O(N__29387),
            .I(N__29384));
    Span4Mux_v I__5202 (
            .O(N__29384),
            .I(N__29381));
    Odrv4 I__5201 (
            .O(N__29381),
            .I(\current_shift_inst.control_input_axb_11 ));
    InMux I__5200 (
            .O(N__29378),
            .I(N__29375));
    LocalMux I__5199 (
            .O(N__29375),
            .I(\current_shift_inst.un38_control_input_0_s1_28 ));
    InMux I__5198 (
            .O(N__29372),
            .I(N__29369));
    LocalMux I__5197 (
            .O(N__29369),
            .I(\current_shift_inst.un38_control_input_0_s0_28 ));
    InMux I__5196 (
            .O(N__29366),
            .I(N__29363));
    LocalMux I__5195 (
            .O(N__29363),
            .I(N__29360));
    Span4Mux_h I__5194 (
            .O(N__29360),
            .I(N__29357));
    Odrv4 I__5193 (
            .O(N__29357),
            .I(\current_shift_inst.control_input_axb_8 ));
    InMux I__5192 (
            .O(N__29354),
            .I(N__29351));
    LocalMux I__5191 (
            .O(N__29351),
            .I(\current_shift_inst.un38_control_input_0_s1_29 ));
    InMux I__5190 (
            .O(N__29348),
            .I(N__29345));
    LocalMux I__5189 (
            .O(N__29345),
            .I(\current_shift_inst.un38_control_input_0_s0_29 ));
    InMux I__5188 (
            .O(N__29342),
            .I(N__29339));
    LocalMux I__5187 (
            .O(N__29339),
            .I(N__29336));
    Span4Mux_h I__5186 (
            .O(N__29336),
            .I(N__29333));
    Odrv4 I__5185 (
            .O(N__29333),
            .I(\current_shift_inst.control_input_axb_9 ));
    InMux I__5184 (
            .O(N__29330),
            .I(N__29327));
    LocalMux I__5183 (
            .O(N__29327),
            .I(\current_shift_inst.un38_control_input_0_s1_30 ));
    InMux I__5182 (
            .O(N__29324),
            .I(N__29321));
    LocalMux I__5181 (
            .O(N__29321),
            .I(\current_shift_inst.un38_control_input_0_s0_30 ));
    CascadeMux I__5180 (
            .O(N__29318),
            .I(N__29315));
    InMux I__5179 (
            .O(N__29315),
            .I(N__29298));
    InMux I__5178 (
            .O(N__29314),
            .I(N__29291));
    InMux I__5177 (
            .O(N__29313),
            .I(N__29291));
    InMux I__5176 (
            .O(N__29312),
            .I(N__29291));
    InMux I__5175 (
            .O(N__29311),
            .I(N__29278));
    InMux I__5174 (
            .O(N__29310),
            .I(N__29278));
    InMux I__5173 (
            .O(N__29309),
            .I(N__29278));
    InMux I__5172 (
            .O(N__29308),
            .I(N__29278));
    InMux I__5171 (
            .O(N__29307),
            .I(N__29278));
    InMux I__5170 (
            .O(N__29306),
            .I(N__29278));
    InMux I__5169 (
            .O(N__29305),
            .I(N__29271));
    InMux I__5168 (
            .O(N__29304),
            .I(N__29271));
    InMux I__5167 (
            .O(N__29303),
            .I(N__29271));
    InMux I__5166 (
            .O(N__29302),
            .I(N__29266));
    InMux I__5165 (
            .O(N__29301),
            .I(N__29266));
    LocalMux I__5164 (
            .O(N__29298),
            .I(N__29263));
    LocalMux I__5163 (
            .O(N__29291),
            .I(N__29260));
    LocalMux I__5162 (
            .O(N__29278),
            .I(N__29257));
    LocalMux I__5161 (
            .O(N__29271),
            .I(N__29252));
    LocalMux I__5160 (
            .O(N__29266),
            .I(N__29252));
    Span4Mux_h I__5159 (
            .O(N__29263),
            .I(N__29249));
    Span4Mux_h I__5158 (
            .O(N__29260),
            .I(N__29246));
    Span4Mux_v I__5157 (
            .O(N__29257),
            .I(N__29243));
    Span4Mux_v I__5156 (
            .O(N__29252),
            .I(N__29240));
    Odrv4 I__5155 (
            .O(N__29249),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__5154 (
            .O(N__29246),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__5153 (
            .O(N__29243),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__5152 (
            .O(N__29240),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    InMux I__5151 (
            .O(N__29231),
            .I(N__29228));
    LocalMux I__5150 (
            .O(N__29228),
            .I(N__29225));
    Span4Mux_v I__5149 (
            .O(N__29225),
            .I(N__29222));
    Odrv4 I__5148 (
            .O(N__29222),
            .I(\current_shift_inst.control_input_axb_10 ));
    CEMux I__5147 (
            .O(N__29219),
            .I(N__29214));
    CEMux I__5146 (
            .O(N__29218),
            .I(N__29211));
    CEMux I__5145 (
            .O(N__29217),
            .I(N__29207));
    LocalMux I__5144 (
            .O(N__29214),
            .I(N__29204));
    LocalMux I__5143 (
            .O(N__29211),
            .I(N__29201));
    CEMux I__5142 (
            .O(N__29210),
            .I(N__29198));
    LocalMux I__5141 (
            .O(N__29207),
            .I(N__29195));
    Span4Mux_v I__5140 (
            .O(N__29204),
            .I(N__29192));
    Span4Mux_v I__5139 (
            .O(N__29201),
            .I(N__29189));
    LocalMux I__5138 (
            .O(N__29198),
            .I(N__29186));
    Span4Mux_h I__5137 (
            .O(N__29195),
            .I(N__29183));
    Span4Mux_h I__5136 (
            .O(N__29192),
            .I(N__29180));
    Span4Mux_h I__5135 (
            .O(N__29189),
            .I(N__29177));
    Span4Mux_h I__5134 (
            .O(N__29186),
            .I(N__29174));
    Span4Mux_v I__5133 (
            .O(N__29183),
            .I(N__29171));
    Span4Mux_v I__5132 (
            .O(N__29180),
            .I(N__29164));
    Span4Mux_v I__5131 (
            .O(N__29177),
            .I(N__29164));
    Span4Mux_v I__5130 (
            .O(N__29174),
            .I(N__29164));
    Odrv4 I__5129 (
            .O(N__29171),
            .I(\delay_measurement_inst.delay_hc_timer.N_199_i ));
    Odrv4 I__5128 (
            .O(N__29164),
            .I(\delay_measurement_inst.delay_hc_timer.N_199_i ));
    InMux I__5127 (
            .O(N__29159),
            .I(N__29153));
    InMux I__5126 (
            .O(N__29158),
            .I(N__29153));
    LocalMux I__5125 (
            .O(N__29153),
            .I(N__29150));
    Span4Mux_h I__5124 (
            .O(N__29150),
            .I(N__29147));
    Span4Mux_h I__5123 (
            .O(N__29147),
            .I(N__29144));
    Span4Mux_h I__5122 (
            .O(N__29144),
            .I(N__29139));
    InMux I__5121 (
            .O(N__29143),
            .I(N__29136));
    InMux I__5120 (
            .O(N__29142),
            .I(N__29133));
    Span4Mux_v I__5119 (
            .O(N__29139),
            .I(N__29130));
    LocalMux I__5118 (
            .O(N__29136),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    LocalMux I__5117 (
            .O(N__29133),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    Odrv4 I__5116 (
            .O(N__29130),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    InMux I__5115 (
            .O(N__29123),
            .I(N__29091));
    InMux I__5114 (
            .O(N__29122),
            .I(N__29091));
    InMux I__5113 (
            .O(N__29121),
            .I(N__29091));
    InMux I__5112 (
            .O(N__29120),
            .I(N__29091));
    InMux I__5111 (
            .O(N__29119),
            .I(N__29082));
    InMux I__5110 (
            .O(N__29118),
            .I(N__29082));
    InMux I__5109 (
            .O(N__29117),
            .I(N__29082));
    InMux I__5108 (
            .O(N__29116),
            .I(N__29082));
    InMux I__5107 (
            .O(N__29115),
            .I(N__29073));
    InMux I__5106 (
            .O(N__29114),
            .I(N__29073));
    InMux I__5105 (
            .O(N__29113),
            .I(N__29073));
    InMux I__5104 (
            .O(N__29112),
            .I(N__29073));
    InMux I__5103 (
            .O(N__29111),
            .I(N__29064));
    InMux I__5102 (
            .O(N__29110),
            .I(N__29064));
    InMux I__5101 (
            .O(N__29109),
            .I(N__29064));
    InMux I__5100 (
            .O(N__29108),
            .I(N__29064));
    InMux I__5099 (
            .O(N__29107),
            .I(N__29049));
    InMux I__5098 (
            .O(N__29106),
            .I(N__29049));
    InMux I__5097 (
            .O(N__29105),
            .I(N__29049));
    InMux I__5096 (
            .O(N__29104),
            .I(N__29049));
    InMux I__5095 (
            .O(N__29103),
            .I(N__29040));
    InMux I__5094 (
            .O(N__29102),
            .I(N__29040));
    InMux I__5093 (
            .O(N__29101),
            .I(N__29040));
    InMux I__5092 (
            .O(N__29100),
            .I(N__29040));
    LocalMux I__5091 (
            .O(N__29091),
            .I(N__29031));
    LocalMux I__5090 (
            .O(N__29082),
            .I(N__29031));
    LocalMux I__5089 (
            .O(N__29073),
            .I(N__29031));
    LocalMux I__5088 (
            .O(N__29064),
            .I(N__29031));
    InMux I__5087 (
            .O(N__29063),
            .I(N__29026));
    InMux I__5086 (
            .O(N__29062),
            .I(N__29026));
    InMux I__5085 (
            .O(N__29061),
            .I(N__29017));
    InMux I__5084 (
            .O(N__29060),
            .I(N__29017));
    InMux I__5083 (
            .O(N__29059),
            .I(N__29017));
    InMux I__5082 (
            .O(N__29058),
            .I(N__29017));
    LocalMux I__5081 (
            .O(N__29049),
            .I(N__29010));
    LocalMux I__5080 (
            .O(N__29040),
            .I(N__29010));
    Span4Mux_v I__5079 (
            .O(N__29031),
            .I(N__29010));
    LocalMux I__5078 (
            .O(N__29026),
            .I(N__29005));
    LocalMux I__5077 (
            .O(N__29017),
            .I(N__29005));
    Span4Mux_h I__5076 (
            .O(N__29010),
            .I(N__29002));
    Span12Mux_h I__5075 (
            .O(N__29005),
            .I(N__28999));
    Span4Mux_v I__5074 (
            .O(N__29002),
            .I(N__28996));
    Odrv12 I__5073 (
            .O(N__28999),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__5072 (
            .O(N__28996),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    InMux I__5071 (
            .O(N__28991),
            .I(N__28988));
    LocalMux I__5070 (
            .O(N__28988),
            .I(N__28985));
    Span4Mux_h I__5069 (
            .O(N__28985),
            .I(N__28982));
    Odrv4 I__5068 (
            .O(N__28982),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ));
    InMux I__5067 (
            .O(N__28979),
            .I(N__28976));
    LocalMux I__5066 (
            .O(N__28976),
            .I(N__28973));
    Odrv4 I__5065 (
            .O(N__28973),
            .I(\current_shift_inst.un38_control_input_0_s0_21 ));
    InMux I__5064 (
            .O(N__28970),
            .I(\current_shift_inst.un38_control_input_cry_20_s0 ));
    InMux I__5063 (
            .O(N__28967),
            .I(N__28964));
    LocalMux I__5062 (
            .O(N__28964),
            .I(N__28961));
    Odrv12 I__5061 (
            .O(N__28961),
            .I(\current_shift_inst.un38_control_input_0_s0_22 ));
    InMux I__5060 (
            .O(N__28958),
            .I(\current_shift_inst.un38_control_input_cry_21_s0 ));
    InMux I__5059 (
            .O(N__28955),
            .I(N__28952));
    LocalMux I__5058 (
            .O(N__28952),
            .I(N__28949));
    Odrv4 I__5057 (
            .O(N__28949),
            .I(\current_shift_inst.un38_control_input_0_s0_23 ));
    InMux I__5056 (
            .O(N__28946),
            .I(\current_shift_inst.un38_control_input_cry_22_s0 ));
    CascadeMux I__5055 (
            .O(N__28943),
            .I(N__28940));
    InMux I__5054 (
            .O(N__28940),
            .I(N__28937));
    LocalMux I__5053 (
            .O(N__28937),
            .I(N__28934));
    Span4Mux_v I__5052 (
            .O(N__28934),
            .I(N__28931));
    Odrv4 I__5051 (
            .O(N__28931),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ));
    InMux I__5050 (
            .O(N__28928),
            .I(N__28925));
    LocalMux I__5049 (
            .O(N__28925),
            .I(N__28922));
    Span4Mux_v I__5048 (
            .O(N__28922),
            .I(N__28919));
    Span4Mux_h I__5047 (
            .O(N__28919),
            .I(N__28916));
    Odrv4 I__5046 (
            .O(N__28916),
            .I(\current_shift_inst.un38_control_input_0_s0_24 ));
    InMux I__5045 (
            .O(N__28913),
            .I(bfn_12_16_0_));
    InMux I__5044 (
            .O(N__28910),
            .I(N__28907));
    LocalMux I__5043 (
            .O(N__28907),
            .I(N__28904));
    Span4Mux_v I__5042 (
            .O(N__28904),
            .I(N__28901));
    Odrv4 I__5041 (
            .O(N__28901),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ));
    InMux I__5040 (
            .O(N__28898),
            .I(N__28895));
    LocalMux I__5039 (
            .O(N__28895),
            .I(N__28892));
    Span4Mux_v I__5038 (
            .O(N__28892),
            .I(N__28889));
    Span4Mux_h I__5037 (
            .O(N__28889),
            .I(N__28886));
    Odrv4 I__5036 (
            .O(N__28886),
            .I(\current_shift_inst.un38_control_input_0_s0_25 ));
    InMux I__5035 (
            .O(N__28883),
            .I(\current_shift_inst.un38_control_input_cry_24_s0 ));
    CascadeMux I__5034 (
            .O(N__28880),
            .I(N__28877));
    InMux I__5033 (
            .O(N__28877),
            .I(N__28874));
    LocalMux I__5032 (
            .O(N__28874),
            .I(N__28871));
    Span4Mux_v I__5031 (
            .O(N__28871),
            .I(N__28868));
    Odrv4 I__5030 (
            .O(N__28868),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ));
    InMux I__5029 (
            .O(N__28865),
            .I(N__28862));
    LocalMux I__5028 (
            .O(N__28862),
            .I(N__28859));
    Span4Mux_h I__5027 (
            .O(N__28859),
            .I(N__28856));
    Odrv4 I__5026 (
            .O(N__28856),
            .I(\current_shift_inst.un38_control_input_0_s0_26 ));
    InMux I__5025 (
            .O(N__28853),
            .I(\current_shift_inst.un38_control_input_cry_25_s0 ));
    InMux I__5024 (
            .O(N__28850),
            .I(N__28847));
    LocalMux I__5023 (
            .O(N__28847),
            .I(N__28844));
    Span4Mux_v I__5022 (
            .O(N__28844),
            .I(N__28841));
    Odrv4 I__5021 (
            .O(N__28841),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ));
    InMux I__5020 (
            .O(N__28838),
            .I(N__28835));
    LocalMux I__5019 (
            .O(N__28835),
            .I(N__28832));
    Span4Mux_h I__5018 (
            .O(N__28832),
            .I(N__28829));
    Odrv4 I__5017 (
            .O(N__28829),
            .I(\current_shift_inst.un38_control_input_0_s0_27 ));
    InMux I__5016 (
            .O(N__28826),
            .I(\current_shift_inst.un38_control_input_cry_26_s0 ));
    CascadeMux I__5015 (
            .O(N__28823),
            .I(N__28820));
    InMux I__5014 (
            .O(N__28820),
            .I(N__28817));
    LocalMux I__5013 (
            .O(N__28817),
            .I(N__28814));
    Span4Mux_v I__5012 (
            .O(N__28814),
            .I(N__28811));
    Odrv4 I__5011 (
            .O(N__28811),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ));
    InMux I__5010 (
            .O(N__28808),
            .I(\current_shift_inst.un38_control_input_cry_27_s0 ));
    InMux I__5009 (
            .O(N__28805),
            .I(N__28802));
    LocalMux I__5008 (
            .O(N__28802),
            .I(N__28799));
    Odrv4 I__5007 (
            .O(N__28799),
            .I(\current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ));
    InMux I__5006 (
            .O(N__28796),
            .I(N__28793));
    LocalMux I__5005 (
            .O(N__28793),
            .I(N__28790));
    Odrv4 I__5004 (
            .O(N__28790),
            .I(\current_shift_inst.un38_control_input_0_s0_20 ));
    InMux I__5003 (
            .O(N__28787),
            .I(\current_shift_inst.un38_control_input_cry_19_s0 ));
    InMux I__5002 (
            .O(N__28784),
            .I(N__28781));
    LocalMux I__5001 (
            .O(N__28781),
            .I(N__28778));
    Span4Mux_h I__5000 (
            .O(N__28778),
            .I(N__28775));
    Odrv4 I__4999 (
            .O(N__28775),
            .I(\current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ));
    CascadeMux I__4998 (
            .O(N__28772),
            .I(N__28769));
    InMux I__4997 (
            .O(N__28769),
            .I(N__28766));
    LocalMux I__4996 (
            .O(N__28766),
            .I(N__28763));
    Span4Mux_v I__4995 (
            .O(N__28763),
            .I(N__28760));
    Span4Mux_h I__4994 (
            .O(N__28760),
            .I(N__28757));
    Odrv4 I__4993 (
            .O(N__28757),
            .I(\current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ));
    InMux I__4992 (
            .O(N__28754),
            .I(N__28751));
    LocalMux I__4991 (
            .O(N__28751),
            .I(N__28748));
    Odrv4 I__4990 (
            .O(N__28748),
            .I(\current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ));
    InMux I__4989 (
            .O(N__28745),
            .I(N__28740));
    InMux I__4988 (
            .O(N__28744),
            .I(N__28736));
    InMux I__4987 (
            .O(N__28743),
            .I(N__28733));
    LocalMux I__4986 (
            .O(N__28740),
            .I(N__28730));
    CascadeMux I__4985 (
            .O(N__28739),
            .I(N__28727));
    LocalMux I__4984 (
            .O(N__28736),
            .I(N__28724));
    LocalMux I__4983 (
            .O(N__28733),
            .I(N__28721));
    Span4Mux_h I__4982 (
            .O(N__28730),
            .I(N__28718));
    InMux I__4981 (
            .O(N__28727),
            .I(N__28715));
    Odrv4 I__4980 (
            .O(N__28724),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    Odrv12 I__4979 (
            .O(N__28721),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    Odrv4 I__4978 (
            .O(N__28718),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    LocalMux I__4977 (
            .O(N__28715),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    InMux I__4976 (
            .O(N__28706),
            .I(N__28702));
    InMux I__4975 (
            .O(N__28705),
            .I(N__28698));
    LocalMux I__4974 (
            .O(N__28702),
            .I(N__28695));
    InMux I__4973 (
            .O(N__28701),
            .I(N__28692));
    LocalMux I__4972 (
            .O(N__28698),
            .I(N__28689));
    Span4Mux_h I__4971 (
            .O(N__28695),
            .I(N__28686));
    LocalMux I__4970 (
            .O(N__28692),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    Odrv4 I__4969 (
            .O(N__28689),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    Odrv4 I__4968 (
            .O(N__28686),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    CascadeMux I__4967 (
            .O(N__28679),
            .I(N__28676));
    InMux I__4966 (
            .O(N__28676),
            .I(N__28673));
    LocalMux I__4965 (
            .O(N__28673),
            .I(N__28670));
    Odrv4 I__4964 (
            .O(N__28670),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ));
    InMux I__4963 (
            .O(N__28667),
            .I(N__28663));
    InMux I__4962 (
            .O(N__28666),
            .I(N__28659));
    LocalMux I__4961 (
            .O(N__28663),
            .I(N__28656));
    InMux I__4960 (
            .O(N__28662),
            .I(N__28653));
    LocalMux I__4959 (
            .O(N__28659),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    Odrv4 I__4958 (
            .O(N__28656),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    LocalMux I__4957 (
            .O(N__28653),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    InMux I__4956 (
            .O(N__28646),
            .I(N__28642));
    InMux I__4955 (
            .O(N__28645),
            .I(N__28637));
    LocalMux I__4954 (
            .O(N__28642),
            .I(N__28634));
    InMux I__4953 (
            .O(N__28641),
            .I(N__28631));
    InMux I__4952 (
            .O(N__28640),
            .I(N__28628));
    LocalMux I__4951 (
            .O(N__28637),
            .I(N__28625));
    Span4Mux_v I__4950 (
            .O(N__28634),
            .I(N__28620));
    LocalMux I__4949 (
            .O(N__28631),
            .I(N__28620));
    LocalMux I__4948 (
            .O(N__28628),
            .I(N__28617));
    Span12Mux_v I__4947 (
            .O(N__28625),
            .I(N__28614));
    Span4Mux_h I__4946 (
            .O(N__28620),
            .I(N__28609));
    Span4Mux_v I__4945 (
            .O(N__28617),
            .I(N__28609));
    Odrv12 I__4944 (
            .O(N__28614),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    Odrv4 I__4943 (
            .O(N__28609),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    CascadeMux I__4942 (
            .O(N__28604),
            .I(N__28601));
    InMux I__4941 (
            .O(N__28601),
            .I(N__28595));
    InMux I__4940 (
            .O(N__28600),
            .I(N__28595));
    LocalMux I__4939 (
            .O(N__28595),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ));
    InMux I__4938 (
            .O(N__28592),
            .I(N__28588));
    InMux I__4937 (
            .O(N__28591),
            .I(N__28585));
    LocalMux I__4936 (
            .O(N__28588),
            .I(N__28581));
    LocalMux I__4935 (
            .O(N__28585),
            .I(N__28578));
    InMux I__4934 (
            .O(N__28584),
            .I(N__28574));
    Span4Mux_h I__4933 (
            .O(N__28581),
            .I(N__28571));
    Span4Mux_v I__4932 (
            .O(N__28578),
            .I(N__28568));
    InMux I__4931 (
            .O(N__28577),
            .I(N__28565));
    LocalMux I__4930 (
            .O(N__28574),
            .I(N__28562));
    Span4Mux_v I__4929 (
            .O(N__28571),
            .I(N__28559));
    Span4Mux_h I__4928 (
            .O(N__28568),
            .I(N__28554));
    LocalMux I__4927 (
            .O(N__28565),
            .I(N__28554));
    Span4Mux_h I__4926 (
            .O(N__28562),
            .I(N__28551));
    Span4Mux_v I__4925 (
            .O(N__28559),
            .I(N__28548));
    Span4Mux_v I__4924 (
            .O(N__28554),
            .I(N__28545));
    Odrv4 I__4923 (
            .O(N__28551),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    Odrv4 I__4922 (
            .O(N__28548),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    Odrv4 I__4921 (
            .O(N__28545),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    InMux I__4920 (
            .O(N__28538),
            .I(N__28535));
    LocalMux I__4919 (
            .O(N__28535),
            .I(N__28531));
    InMux I__4918 (
            .O(N__28534),
            .I(N__28527));
    Span4Mux_v I__4917 (
            .O(N__28531),
            .I(N__28524));
    InMux I__4916 (
            .O(N__28530),
            .I(N__28521));
    LocalMux I__4915 (
            .O(N__28527),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    Odrv4 I__4914 (
            .O(N__28524),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    LocalMux I__4913 (
            .O(N__28521),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    CEMux I__4912 (
            .O(N__28514),
            .I(N__28475));
    CEMux I__4911 (
            .O(N__28513),
            .I(N__28475));
    CEMux I__4910 (
            .O(N__28512),
            .I(N__28475));
    CEMux I__4909 (
            .O(N__28511),
            .I(N__28475));
    CEMux I__4908 (
            .O(N__28510),
            .I(N__28475));
    CEMux I__4907 (
            .O(N__28509),
            .I(N__28475));
    CEMux I__4906 (
            .O(N__28508),
            .I(N__28475));
    CEMux I__4905 (
            .O(N__28507),
            .I(N__28475));
    CEMux I__4904 (
            .O(N__28506),
            .I(N__28475));
    CEMux I__4903 (
            .O(N__28505),
            .I(N__28475));
    CEMux I__4902 (
            .O(N__28504),
            .I(N__28475));
    CEMux I__4901 (
            .O(N__28503),
            .I(N__28475));
    CEMux I__4900 (
            .O(N__28502),
            .I(N__28475));
    GlobalMux I__4899 (
            .O(N__28475),
            .I(N__28472));
    gio2CtrlBuf I__4898 (
            .O(N__28472),
            .I(\phase_controller_inst2.stoper_hc.un1_start_g ));
    InMux I__4897 (
            .O(N__28469),
            .I(N__28466));
    LocalMux I__4896 (
            .O(N__28466),
            .I(N__28463));
    Span4Mux_h I__4895 (
            .O(N__28463),
            .I(N__28459));
    InMux I__4894 (
            .O(N__28462),
            .I(N__28456));
    Odrv4 I__4893 (
            .O(N__28459),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ));
    LocalMux I__4892 (
            .O(N__28456),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ));
    InMux I__4891 (
            .O(N__28451),
            .I(N__28446));
    InMux I__4890 (
            .O(N__28450),
            .I(N__28443));
    InMux I__4889 (
            .O(N__28449),
            .I(N__28440));
    LocalMux I__4888 (
            .O(N__28446),
            .I(N__28437));
    LocalMux I__4887 (
            .O(N__28443),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    LocalMux I__4886 (
            .O(N__28440),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    Odrv4 I__4885 (
            .O(N__28437),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    CascadeMux I__4884 (
            .O(N__28430),
            .I(N__28427));
    InMux I__4883 (
            .O(N__28427),
            .I(N__28423));
    CascadeMux I__4882 (
            .O(N__28426),
            .I(N__28419));
    LocalMux I__4881 (
            .O(N__28423),
            .I(N__28416));
    InMux I__4880 (
            .O(N__28422),
            .I(N__28413));
    InMux I__4879 (
            .O(N__28419),
            .I(N__28410));
    Span4Mux_h I__4878 (
            .O(N__28416),
            .I(N__28407));
    LocalMux I__4877 (
            .O(N__28413),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    LocalMux I__4876 (
            .O(N__28410),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    Odrv4 I__4875 (
            .O(N__28407),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    InMux I__4874 (
            .O(N__28400),
            .I(N__28397));
    LocalMux I__4873 (
            .O(N__28397),
            .I(N__28394));
    Span4Mux_v I__4872 (
            .O(N__28394),
            .I(N__28390));
    InMux I__4871 (
            .O(N__28393),
            .I(N__28387));
    Odrv4 I__4870 (
            .O(N__28390),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ));
    LocalMux I__4869 (
            .O(N__28387),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ));
    CascadeMux I__4868 (
            .O(N__28382),
            .I(N__28379));
    InMux I__4867 (
            .O(N__28379),
            .I(N__28376));
    LocalMux I__4866 (
            .O(N__28376),
            .I(N__28373));
    Span4Mux_h I__4865 (
            .O(N__28373),
            .I(N__28370));
    Odrv4 I__4864 (
            .O(N__28370),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ));
    InMux I__4863 (
            .O(N__28367),
            .I(N__28363));
    InMux I__4862 (
            .O(N__28366),
            .I(N__28360));
    LocalMux I__4861 (
            .O(N__28363),
            .I(N__28357));
    LocalMux I__4860 (
            .O(N__28360),
            .I(N__28354));
    Span4Mux_h I__4859 (
            .O(N__28357),
            .I(N__28351));
    Span4Mux_v I__4858 (
            .O(N__28354),
            .I(N__28348));
    Odrv4 I__4857 (
            .O(N__28351),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    Odrv4 I__4856 (
            .O(N__28348),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    CascadeMux I__4855 (
            .O(N__28343),
            .I(N__28340));
    InMux I__4854 (
            .O(N__28340),
            .I(N__28337));
    LocalMux I__4853 (
            .O(N__28337),
            .I(N__28334));
    Odrv4 I__4852 (
            .O(N__28334),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2 ));
    CascadeMux I__4851 (
            .O(N__28331),
            .I(N__28327));
    InMux I__4850 (
            .O(N__28330),
            .I(N__28321));
    InMux I__4849 (
            .O(N__28327),
            .I(N__28321));
    InMux I__4848 (
            .O(N__28326),
            .I(N__28318));
    LocalMux I__4847 (
            .O(N__28321),
            .I(N__28314));
    LocalMux I__4846 (
            .O(N__28318),
            .I(N__28311));
    InMux I__4845 (
            .O(N__28317),
            .I(N__28308));
    Odrv4 I__4844 (
            .O(N__28314),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    Odrv4 I__4843 (
            .O(N__28311),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    LocalMux I__4842 (
            .O(N__28308),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    InMux I__4841 (
            .O(N__28301),
            .I(N__28298));
    LocalMux I__4840 (
            .O(N__28298),
            .I(N__28294));
    InMux I__4839 (
            .O(N__28297),
            .I(N__28291));
    Span4Mux_h I__4838 (
            .O(N__28294),
            .I(N__28288));
    LocalMux I__4837 (
            .O(N__28291),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    Odrv4 I__4836 (
            .O(N__28288),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    InMux I__4835 (
            .O(N__28283),
            .I(N__28280));
    LocalMux I__4834 (
            .O(N__28280),
            .I(N__28274));
    InMux I__4833 (
            .O(N__28279),
            .I(N__28267));
    InMux I__4832 (
            .O(N__28278),
            .I(N__28267));
    InMux I__4831 (
            .O(N__28277),
            .I(N__28267));
    Odrv12 I__4830 (
            .O(N__28274),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    LocalMux I__4829 (
            .O(N__28267),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    CascadeMux I__4828 (
            .O(N__28262),
            .I(N__28258));
    InMux I__4827 (
            .O(N__28261),
            .I(N__28247));
    InMux I__4826 (
            .O(N__28258),
            .I(N__28247));
    InMux I__4825 (
            .O(N__28257),
            .I(N__28247));
    InMux I__4824 (
            .O(N__28256),
            .I(N__28247));
    LocalMux I__4823 (
            .O(N__28247),
            .I(N__28244));
    Span4Mux_h I__4822 (
            .O(N__28244),
            .I(N__28241));
    Odrv4 I__4821 (
            .O(N__28241),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    InMux I__4820 (
            .O(N__28238),
            .I(N__28234));
    InMux I__4819 (
            .O(N__28237),
            .I(N__28231));
    LocalMux I__4818 (
            .O(N__28234),
            .I(N__28228));
    LocalMux I__4817 (
            .O(N__28231),
            .I(N__28225));
    Span4Mux_h I__4816 (
            .O(N__28228),
            .I(N__28222));
    Span4Mux_h I__4815 (
            .O(N__28225),
            .I(N__28219));
    Odrv4 I__4814 (
            .O(N__28222),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ));
    Odrv4 I__4813 (
            .O(N__28219),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ));
    CascadeMux I__4812 (
            .O(N__28214),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0_cascade_ ));
    InMux I__4811 (
            .O(N__28211),
            .I(N__28204));
    InMux I__4810 (
            .O(N__28210),
            .I(N__28204));
    InMux I__4809 (
            .O(N__28209),
            .I(N__28201));
    LocalMux I__4808 (
            .O(N__28204),
            .I(N__28198));
    LocalMux I__4807 (
            .O(N__28201),
            .I(N__28193));
    Span4Mux_v I__4806 (
            .O(N__28198),
            .I(N__28190));
    InMux I__4805 (
            .O(N__28197),
            .I(N__28185));
    InMux I__4804 (
            .O(N__28196),
            .I(N__28185));
    Odrv12 I__4803 (
            .O(N__28193),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    Odrv4 I__4802 (
            .O(N__28190),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    LocalMux I__4801 (
            .O(N__28185),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    InMux I__4800 (
            .O(N__28178),
            .I(N__28175));
    LocalMux I__4799 (
            .O(N__28175),
            .I(N__28170));
    InMux I__4798 (
            .O(N__28174),
            .I(N__28167));
    InMux I__4797 (
            .O(N__28173),
            .I(N__28163));
    Span4Mux_v I__4796 (
            .O(N__28170),
            .I(N__28158));
    LocalMux I__4795 (
            .O(N__28167),
            .I(N__28158));
    InMux I__4794 (
            .O(N__28166),
            .I(N__28155));
    LocalMux I__4793 (
            .O(N__28163),
            .I(N__28152));
    Span4Mux_h I__4792 (
            .O(N__28158),
            .I(N__28149));
    LocalMux I__4791 (
            .O(N__28155),
            .I(N__28146));
    Span4Mux_v I__4790 (
            .O(N__28152),
            .I(N__28143));
    Span4Mux_v I__4789 (
            .O(N__28149),
            .I(N__28140));
    Span4Mux_v I__4788 (
            .O(N__28146),
            .I(N__28137));
    Odrv4 I__4787 (
            .O(N__28143),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    Odrv4 I__4786 (
            .O(N__28140),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    Odrv4 I__4785 (
            .O(N__28137),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    InMux I__4784 (
            .O(N__28130),
            .I(N__28127));
    LocalMux I__4783 (
            .O(N__28127),
            .I(N__28122));
    InMux I__4782 (
            .O(N__28126),
            .I(N__28119));
    InMux I__4781 (
            .O(N__28125),
            .I(N__28116));
    Span4Mux_v I__4780 (
            .O(N__28122),
            .I(N__28113));
    LocalMux I__4779 (
            .O(N__28119),
            .I(N__28110));
    LocalMux I__4778 (
            .O(N__28116),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    Odrv4 I__4777 (
            .O(N__28113),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    Odrv4 I__4776 (
            .O(N__28110),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    InMux I__4775 (
            .O(N__28103),
            .I(N__28100));
    LocalMux I__4774 (
            .O(N__28100),
            .I(N__28097));
    Span4Mux_v I__4773 (
            .O(N__28097),
            .I(N__28094));
    Odrv4 I__4772 (
            .O(N__28094),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ));
    InMux I__4771 (
            .O(N__28091),
            .I(N__28084));
    InMux I__4770 (
            .O(N__28090),
            .I(N__28084));
    InMux I__4769 (
            .O(N__28089),
            .I(N__28081));
    LocalMux I__4768 (
            .O(N__28084),
            .I(N__28078));
    LocalMux I__4767 (
            .O(N__28081),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ));
    Odrv4 I__4766 (
            .O(N__28078),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ));
    CascadeMux I__4765 (
            .O(N__28073),
            .I(N__28070));
    InMux I__4764 (
            .O(N__28070),
            .I(N__28064));
    InMux I__4763 (
            .O(N__28069),
            .I(N__28064));
    LocalMux I__4762 (
            .O(N__28064),
            .I(N__28061));
    Span4Mux_h I__4761 (
            .O(N__28061),
            .I(N__28058));
    Span4Mux_h I__4760 (
            .O(N__28058),
            .I(N__28055));
    Odrv4 I__4759 (
            .O(N__28055),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ));
    CascadeMux I__4758 (
            .O(N__28052),
            .I(N__28048));
    InMux I__4757 (
            .O(N__28051),
            .I(N__28043));
    InMux I__4756 (
            .O(N__28048),
            .I(N__28043));
    LocalMux I__4755 (
            .O(N__28043),
            .I(N__28039));
    InMux I__4754 (
            .O(N__28042),
            .I(N__28036));
    Span4Mux_h I__4753 (
            .O(N__28039),
            .I(N__28033));
    LocalMux I__4752 (
            .O(N__28036),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ));
    Odrv4 I__4751 (
            .O(N__28033),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ));
    InMux I__4750 (
            .O(N__28028),
            .I(N__28022));
    InMux I__4749 (
            .O(N__28027),
            .I(N__28022));
    LocalMux I__4748 (
            .O(N__28022),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ));
    CascadeMux I__4747 (
            .O(N__28019),
            .I(N__28016));
    InMux I__4746 (
            .O(N__28016),
            .I(N__28013));
    LocalMux I__4745 (
            .O(N__28013),
            .I(N__28010));
    Span4Mux_h I__4744 (
            .O(N__28010),
            .I(N__28007));
    Odrv4 I__4743 (
            .O(N__28007),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt28 ));
    CascadeMux I__4742 (
            .O(N__28004),
            .I(N__28001));
    InMux I__4741 (
            .O(N__28001),
            .I(N__27998));
    LocalMux I__4740 (
            .O(N__27998),
            .I(N__27995));
    Span4Mux_h I__4739 (
            .O(N__27995),
            .I(N__27992));
    Odrv4 I__4738 (
            .O(N__27992),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt24 ));
    InMux I__4737 (
            .O(N__27989),
            .I(N__27984));
    InMux I__4736 (
            .O(N__27988),
            .I(N__27979));
    InMux I__4735 (
            .O(N__27987),
            .I(N__27979));
    LocalMux I__4734 (
            .O(N__27984),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ));
    LocalMux I__4733 (
            .O(N__27979),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ));
    CascadeMux I__4732 (
            .O(N__27974),
            .I(N__27971));
    InMux I__4731 (
            .O(N__27971),
            .I(N__27964));
    InMux I__4730 (
            .O(N__27970),
            .I(N__27964));
    InMux I__4729 (
            .O(N__27969),
            .I(N__27961));
    LocalMux I__4728 (
            .O(N__27964),
            .I(N__27958));
    LocalMux I__4727 (
            .O(N__27961),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ));
    Odrv4 I__4726 (
            .O(N__27958),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ));
    InMux I__4725 (
            .O(N__27953),
            .I(N__27950));
    LocalMux I__4724 (
            .O(N__27950),
            .I(N__27947));
    Span4Mux_h I__4723 (
            .O(N__27947),
            .I(N__27944));
    Odrv4 I__4722 (
            .O(N__27944),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ));
    InMux I__4721 (
            .O(N__27941),
            .I(N__27935));
    InMux I__4720 (
            .O(N__27940),
            .I(N__27935));
    LocalMux I__4719 (
            .O(N__27935),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ));
    CascadeMux I__4718 (
            .O(N__27932),
            .I(N__27928));
    InMux I__4717 (
            .O(N__27931),
            .I(N__27923));
    InMux I__4716 (
            .O(N__27928),
            .I(N__27923));
    LocalMux I__4715 (
            .O(N__27923),
            .I(N__27919));
    InMux I__4714 (
            .O(N__27922),
            .I(N__27916));
    Span4Mux_h I__4713 (
            .O(N__27919),
            .I(N__27913));
    LocalMux I__4712 (
            .O(N__27916),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ));
    Odrv4 I__4711 (
            .O(N__27913),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ));
    InMux I__4710 (
            .O(N__27908),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ));
    InMux I__4709 (
            .O(N__27905),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ));
    InMux I__4708 (
            .O(N__27902),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ));
    InMux I__4707 (
            .O(N__27899),
            .I(N__27889));
    InMux I__4706 (
            .O(N__27898),
            .I(N__27889));
    InMux I__4705 (
            .O(N__27897),
            .I(N__27889));
    InMux I__4704 (
            .O(N__27896),
            .I(N__27886));
    LocalMux I__4703 (
            .O(N__27889),
            .I(N__27883));
    LocalMux I__4702 (
            .O(N__27886),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    Odrv4 I__4701 (
            .O(N__27883),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    InMux I__4700 (
            .O(N__27878),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ));
    InMux I__4699 (
            .O(N__27875),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ));
    CascadeMux I__4698 (
            .O(N__27872),
            .I(N__27867));
    CascadeMux I__4697 (
            .O(N__27871),
            .I(N__27864));
    InMux I__4696 (
            .O(N__27870),
            .I(N__27857));
    InMux I__4695 (
            .O(N__27867),
            .I(N__27857));
    InMux I__4694 (
            .O(N__27864),
            .I(N__27857));
    LocalMux I__4693 (
            .O(N__27857),
            .I(N__27853));
    InMux I__4692 (
            .O(N__27856),
            .I(N__27850));
    Span4Mux_h I__4691 (
            .O(N__27853),
            .I(N__27847));
    LocalMux I__4690 (
            .O(N__27850),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    Odrv4 I__4689 (
            .O(N__27847),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    InMux I__4688 (
            .O(N__27842),
            .I(N__27839));
    LocalMux I__4687 (
            .O(N__27839),
            .I(N__27836));
    Span4Mux_v I__4686 (
            .O(N__27836),
            .I(N__27831));
    InMux I__4685 (
            .O(N__27835),
            .I(N__27828));
    InMux I__4684 (
            .O(N__27834),
            .I(N__27825));
    Odrv4 I__4683 (
            .O(N__27831),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ));
    LocalMux I__4682 (
            .O(N__27828),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ));
    LocalMux I__4681 (
            .O(N__27825),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ));
    InMux I__4680 (
            .O(N__27818),
            .I(N__27815));
    LocalMux I__4679 (
            .O(N__27815),
            .I(N__27810));
    InMux I__4678 (
            .O(N__27814),
            .I(N__27807));
    InMux I__4677 (
            .O(N__27813),
            .I(N__27804));
    Span4Mux_h I__4676 (
            .O(N__27810),
            .I(N__27799));
    LocalMux I__4675 (
            .O(N__27807),
            .I(N__27799));
    LocalMux I__4674 (
            .O(N__27804),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__4673 (
            .O(N__27799),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__4672 (
            .O(N__27794),
            .I(N__27790));
    InMux I__4671 (
            .O(N__27793),
            .I(N__27787));
    LocalMux I__4670 (
            .O(N__27790),
            .I(N__27784));
    LocalMux I__4669 (
            .O(N__27787),
            .I(N__27781));
    Odrv12 I__4668 (
            .O(N__27784),
            .I(\phase_controller_inst2.state_RNIG7JFZ0Z_2 ));
    Odrv12 I__4667 (
            .O(N__27781),
            .I(\phase_controller_inst2.state_RNIG7JFZ0Z_2 ));
    InMux I__4666 (
            .O(N__27776),
            .I(N__27769));
    InMux I__4665 (
            .O(N__27775),
            .I(N__27769));
    InMux I__4664 (
            .O(N__27774),
            .I(N__27766));
    LocalMux I__4663 (
            .O(N__27769),
            .I(N__27763));
    LocalMux I__4662 (
            .O(N__27766),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv4 I__4661 (
            .O(N__27763),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__4660 (
            .O(N__27758),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ));
    InMux I__4659 (
            .O(N__27755),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ));
    InMux I__4658 (
            .O(N__27752),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__4657 (
            .O(N__27749),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ));
    InMux I__4656 (
            .O(N__27746),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ));
    CascadeMux I__4655 (
            .O(N__27743),
            .I(N__27740));
    InMux I__4654 (
            .O(N__27740),
            .I(N__27736));
    InMux I__4653 (
            .O(N__27739),
            .I(N__27732));
    LocalMux I__4652 (
            .O(N__27736),
            .I(N__27729));
    InMux I__4651 (
            .O(N__27735),
            .I(N__27726));
    LocalMux I__4650 (
            .O(N__27732),
            .I(N__27723));
    Span4Mux_h I__4649 (
            .O(N__27729),
            .I(N__27720));
    LocalMux I__4648 (
            .O(N__27726),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    Odrv4 I__4647 (
            .O(N__27723),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    Odrv4 I__4646 (
            .O(N__27720),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    InMux I__4645 (
            .O(N__27713),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ));
    InMux I__4644 (
            .O(N__27710),
            .I(N__27706));
    InMux I__4643 (
            .O(N__27709),
            .I(N__27703));
    LocalMux I__4642 (
            .O(N__27706),
            .I(N__27699));
    LocalMux I__4641 (
            .O(N__27703),
            .I(N__27696));
    InMux I__4640 (
            .O(N__27702),
            .I(N__27693));
    Span4Mux_v I__4639 (
            .O(N__27699),
            .I(N__27690));
    Span4Mux_h I__4638 (
            .O(N__27696),
            .I(N__27687));
    LocalMux I__4637 (
            .O(N__27693),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    Odrv4 I__4636 (
            .O(N__27690),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    Odrv4 I__4635 (
            .O(N__27687),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    InMux I__4634 (
            .O(N__27680),
            .I(bfn_12_9_0_));
    CascadeMux I__4633 (
            .O(N__27677),
            .I(N__27673));
    InMux I__4632 (
            .O(N__27676),
            .I(N__27668));
    InMux I__4631 (
            .O(N__27673),
            .I(N__27668));
    LocalMux I__4630 (
            .O(N__27668),
            .I(N__27664));
    InMux I__4629 (
            .O(N__27667),
            .I(N__27661));
    Span4Mux_h I__4628 (
            .O(N__27664),
            .I(N__27658));
    LocalMux I__4627 (
            .O(N__27661),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ));
    Odrv4 I__4626 (
            .O(N__27658),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ));
    InMux I__4625 (
            .O(N__27653),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ));
    InMux I__4624 (
            .O(N__27650),
            .I(N__27646));
    InMux I__4623 (
            .O(N__27649),
            .I(N__27643));
    LocalMux I__4622 (
            .O(N__27646),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__4621 (
            .O(N__27643),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__4620 (
            .O(N__27638),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__4619 (
            .O(N__27635),
            .I(N__27631));
    InMux I__4618 (
            .O(N__27634),
            .I(N__27628));
    LocalMux I__4617 (
            .O(N__27631),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__4616 (
            .O(N__27628),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__4615 (
            .O(N__27623),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__4614 (
            .O(N__27620),
            .I(N__27616));
    InMux I__4613 (
            .O(N__27619),
            .I(N__27613));
    LocalMux I__4612 (
            .O(N__27616),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    LocalMux I__4611 (
            .O(N__27613),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__4610 (
            .O(N__27608),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__4609 (
            .O(N__27605),
            .I(N__27601));
    InMux I__4608 (
            .O(N__27604),
            .I(N__27598));
    LocalMux I__4607 (
            .O(N__27601),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    LocalMux I__4606 (
            .O(N__27598),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__4605 (
            .O(N__27593),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__4604 (
            .O(N__27590),
            .I(N__27586));
    InMux I__4603 (
            .O(N__27589),
            .I(N__27583));
    LocalMux I__4602 (
            .O(N__27586),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__4601 (
            .O(N__27583),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__4600 (
            .O(N__27578),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__4599 (
            .O(N__27575),
            .I(N__27571));
    InMux I__4598 (
            .O(N__27574),
            .I(N__27568));
    LocalMux I__4597 (
            .O(N__27571),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__4596 (
            .O(N__27568),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__4595 (
            .O(N__27563),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ));
    InMux I__4594 (
            .O(N__27560),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ));
    InMux I__4593 (
            .O(N__27557),
            .I(bfn_12_8_0_));
    CascadeMux I__4592 (
            .O(N__27554),
            .I(N__27550));
    InMux I__4591 (
            .O(N__27553),
            .I(N__27544));
    InMux I__4590 (
            .O(N__27550),
            .I(N__27544));
    InMux I__4589 (
            .O(N__27549),
            .I(N__27541));
    LocalMux I__4588 (
            .O(N__27544),
            .I(N__27538));
    LocalMux I__4587 (
            .O(N__27541),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv4 I__4586 (
            .O(N__27538),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__4585 (
            .O(N__27533),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ));
    InMux I__4584 (
            .O(N__27530),
            .I(N__27526));
    InMux I__4583 (
            .O(N__27529),
            .I(N__27523));
    LocalMux I__4582 (
            .O(N__27526),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__4581 (
            .O(N__27523),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__4580 (
            .O(N__27518),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ));
    CascadeMux I__4579 (
            .O(N__27515),
            .I(N__27512));
    InMux I__4578 (
            .O(N__27512),
            .I(N__27509));
    LocalMux I__4577 (
            .O(N__27509),
            .I(N__27506));
    Odrv4 I__4576 (
            .O(N__27506),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28 ));
    InMux I__4575 (
            .O(N__27503),
            .I(N__27499));
    InMux I__4574 (
            .O(N__27502),
            .I(N__27496));
    LocalMux I__4573 (
            .O(N__27499),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__4572 (
            .O(N__27496),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__4571 (
            .O(N__27491),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__4570 (
            .O(N__27488),
            .I(N__27484));
    InMux I__4569 (
            .O(N__27487),
            .I(N__27481));
    LocalMux I__4568 (
            .O(N__27484),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__4567 (
            .O(N__27481),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__4566 (
            .O(N__27476),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__4565 (
            .O(N__27473),
            .I(N__27469));
    InMux I__4564 (
            .O(N__27472),
            .I(N__27466));
    LocalMux I__4563 (
            .O(N__27469),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__4562 (
            .O(N__27466),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__4561 (
            .O(N__27461),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__4560 (
            .O(N__27458),
            .I(N__27454));
    InMux I__4559 (
            .O(N__27457),
            .I(N__27451));
    LocalMux I__4558 (
            .O(N__27454),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__4557 (
            .O(N__27451),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__4556 (
            .O(N__27446),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__4555 (
            .O(N__27443),
            .I(N__27439));
    InMux I__4554 (
            .O(N__27442),
            .I(N__27436));
    LocalMux I__4553 (
            .O(N__27439),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__4552 (
            .O(N__27436),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__4551 (
            .O(N__27431),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__4550 (
            .O(N__27428),
            .I(N__27424));
    InMux I__4549 (
            .O(N__27427),
            .I(N__27421));
    LocalMux I__4548 (
            .O(N__27424),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__4547 (
            .O(N__27421),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__4546 (
            .O(N__27416),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__4545 (
            .O(N__27413),
            .I(N__27409));
    InMux I__4544 (
            .O(N__27412),
            .I(N__27406));
    LocalMux I__4543 (
            .O(N__27409),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__4542 (
            .O(N__27406),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__4541 (
            .O(N__27401),
            .I(bfn_12_7_0_));
    InMux I__4540 (
            .O(N__27398),
            .I(N__27395));
    LocalMux I__4539 (
            .O(N__27395),
            .I(\pwm_generator_inst.counter_i_9 ));
    InMux I__4538 (
            .O(N__27392),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    IoInMux I__4537 (
            .O(N__27389),
            .I(N__27386));
    LocalMux I__4536 (
            .O(N__27386),
            .I(N__27383));
    IoSpan4Mux I__4535 (
            .O(N__27383),
            .I(N__27380));
    Sp12to4 I__4534 (
            .O(N__27380),
            .I(N__27377));
    Span12Mux_s9_v I__4533 (
            .O(N__27377),
            .I(N__27374));
    Span12Mux_h I__4532 (
            .O(N__27374),
            .I(N__27371));
    Span12Mux_v I__4531 (
            .O(N__27371),
            .I(N__27368));
    Odrv12 I__4530 (
            .O(N__27368),
            .I(pwm_output_c));
    IoInMux I__4529 (
            .O(N__27365),
            .I(N__27362));
    LocalMux I__4528 (
            .O(N__27362),
            .I(N__27359));
    Span12Mux_s3_v I__4527 (
            .O(N__27359),
            .I(N__27356));
    Odrv12 I__4526 (
            .O(N__27356),
            .I(s3_phy_c));
    InMux I__4525 (
            .O(N__27353),
            .I(N__27350));
    LocalMux I__4524 (
            .O(N__27350),
            .I(N__27347));
    Span4Mux_v I__4523 (
            .O(N__27347),
            .I(N__27344));
    Odrv4 I__4522 (
            .O(N__27344),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ));
    InMux I__4521 (
            .O(N__27341),
            .I(N__27335));
    InMux I__4520 (
            .O(N__27340),
            .I(N__27335));
    LocalMux I__4519 (
            .O(N__27335),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ));
    InMux I__4518 (
            .O(N__27332),
            .I(N__27329));
    LocalMux I__4517 (
            .O(N__27329),
            .I(N__27324));
    InMux I__4516 (
            .O(N__27328),
            .I(N__27321));
    InMux I__4515 (
            .O(N__27327),
            .I(N__27318));
    Span4Mux_h I__4514 (
            .O(N__27324),
            .I(N__27315));
    LocalMux I__4513 (
            .O(N__27321),
            .I(N__27312));
    LocalMux I__4512 (
            .O(N__27318),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    Odrv4 I__4511 (
            .O(N__27315),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    Odrv4 I__4510 (
            .O(N__27312),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    InMux I__4509 (
            .O(N__27305),
            .I(N__27302));
    LocalMux I__4508 (
            .O(N__27302),
            .I(N__27298));
    InMux I__4507 (
            .O(N__27301),
            .I(N__27293));
    Span4Mux_h I__4506 (
            .O(N__27298),
            .I(N__27290));
    InMux I__4505 (
            .O(N__27297),
            .I(N__27285));
    InMux I__4504 (
            .O(N__27296),
            .I(N__27285));
    LocalMux I__4503 (
            .O(N__27293),
            .I(N__27282));
    Span4Mux_v I__4502 (
            .O(N__27290),
            .I(N__27277));
    LocalMux I__4501 (
            .O(N__27285),
            .I(N__27277));
    Span4Mux_v I__4500 (
            .O(N__27282),
            .I(N__27274));
    Span4Mux_h I__4499 (
            .O(N__27277),
            .I(N__27271));
    Odrv4 I__4498 (
            .O(N__27274),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    Odrv4 I__4497 (
            .O(N__27271),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    CascadeMux I__4496 (
            .O(N__27266),
            .I(N__27263));
    InMux I__4495 (
            .O(N__27263),
            .I(N__27260));
    LocalMux I__4494 (
            .O(N__27260),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ));
    InMux I__4493 (
            .O(N__27257),
            .I(N__27254));
    LocalMux I__4492 (
            .O(N__27254),
            .I(\pwm_generator_inst.counter_i_0 ));
    InMux I__4491 (
            .O(N__27251),
            .I(N__27248));
    LocalMux I__4490 (
            .O(N__27248),
            .I(\pwm_generator_inst.counter_i_1 ));
    InMux I__4489 (
            .O(N__27245),
            .I(N__27242));
    LocalMux I__4488 (
            .O(N__27242),
            .I(\pwm_generator_inst.counter_i_2 ));
    InMux I__4487 (
            .O(N__27239),
            .I(N__27236));
    LocalMux I__4486 (
            .O(N__27236),
            .I(\pwm_generator_inst.counter_i_3 ));
    InMux I__4485 (
            .O(N__27233),
            .I(N__27230));
    LocalMux I__4484 (
            .O(N__27230),
            .I(\pwm_generator_inst.counter_i_4 ));
    InMux I__4483 (
            .O(N__27227),
            .I(N__27224));
    LocalMux I__4482 (
            .O(N__27224),
            .I(\pwm_generator_inst.counter_i_5 ));
    InMux I__4481 (
            .O(N__27221),
            .I(N__27218));
    LocalMux I__4480 (
            .O(N__27218),
            .I(\pwm_generator_inst.counter_i_6 ));
    InMux I__4479 (
            .O(N__27215),
            .I(N__27212));
    LocalMux I__4478 (
            .O(N__27212),
            .I(\pwm_generator_inst.counter_i_7 ));
    InMux I__4477 (
            .O(N__27209),
            .I(N__27206));
    LocalMux I__4476 (
            .O(N__27206),
            .I(\pwm_generator_inst.counter_i_8 ));
    CascadeMux I__4475 (
            .O(N__27203),
            .I(N__27200));
    InMux I__4474 (
            .O(N__27200),
            .I(N__27197));
    LocalMux I__4473 (
            .O(N__27197),
            .I(N__27194));
    Odrv4 I__4472 (
            .O(N__27194),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ));
    InMux I__4471 (
            .O(N__27191),
            .I(N__27184));
    InMux I__4470 (
            .O(N__27190),
            .I(N__27184));
    InMux I__4469 (
            .O(N__27189),
            .I(N__27181));
    LocalMux I__4468 (
            .O(N__27184),
            .I(N__27177));
    LocalMux I__4467 (
            .O(N__27181),
            .I(N__27174));
    InMux I__4466 (
            .O(N__27180),
            .I(N__27171));
    Span4Mux_h I__4465 (
            .O(N__27177),
            .I(N__27168));
    Span4Mux_v I__4464 (
            .O(N__27174),
            .I(N__27163));
    LocalMux I__4463 (
            .O(N__27171),
            .I(N__27163));
    Odrv4 I__4462 (
            .O(N__27168),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    Odrv4 I__4461 (
            .O(N__27163),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    CascadeMux I__4460 (
            .O(N__27158),
            .I(N__27155));
    InMux I__4459 (
            .O(N__27155),
            .I(N__27149));
    InMux I__4458 (
            .O(N__27154),
            .I(N__27149));
    LocalMux I__4457 (
            .O(N__27149),
            .I(N__27145));
    InMux I__4456 (
            .O(N__27148),
            .I(N__27142));
    Odrv4 I__4455 (
            .O(N__27145),
            .I(\current_shift_inst.un4_control_input1_26 ));
    LocalMux I__4454 (
            .O(N__27142),
            .I(\current_shift_inst.un4_control_input1_26 ));
    InMux I__4453 (
            .O(N__27137),
            .I(N__27134));
    LocalMux I__4452 (
            .O(N__27134),
            .I(N__27131));
    Odrv4 I__4451 (
            .O(N__27131),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ));
    InMux I__4450 (
            .O(N__27128),
            .I(N__27123));
    InMux I__4449 (
            .O(N__27127),
            .I(N__27120));
    InMux I__4448 (
            .O(N__27126),
            .I(N__27116));
    LocalMux I__4447 (
            .O(N__27123),
            .I(N__27113));
    LocalMux I__4446 (
            .O(N__27120),
            .I(N__27110));
    InMux I__4445 (
            .O(N__27119),
            .I(N__27107));
    LocalMux I__4444 (
            .O(N__27116),
            .I(N__27104));
    Span4Mux_v I__4443 (
            .O(N__27113),
            .I(N__27097));
    Span4Mux_v I__4442 (
            .O(N__27110),
            .I(N__27097));
    LocalMux I__4441 (
            .O(N__27107),
            .I(N__27097));
    Span4Mux_v I__4440 (
            .O(N__27104),
            .I(N__27094));
    Span4Mux_h I__4439 (
            .O(N__27097),
            .I(N__27091));
    Odrv4 I__4438 (
            .O(N__27094),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    Odrv4 I__4437 (
            .O(N__27091),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    InMux I__4436 (
            .O(N__27086),
            .I(N__27081));
    CascadeMux I__4435 (
            .O(N__27085),
            .I(N__27078));
    CascadeMux I__4434 (
            .O(N__27084),
            .I(N__27075));
    LocalMux I__4433 (
            .O(N__27081),
            .I(N__27072));
    InMux I__4432 (
            .O(N__27078),
            .I(N__27069));
    InMux I__4431 (
            .O(N__27075),
            .I(N__27066));
    Span4Mux_h I__4430 (
            .O(N__27072),
            .I(N__27063));
    LocalMux I__4429 (
            .O(N__27069),
            .I(\current_shift_inst.un4_control_input1_29 ));
    LocalMux I__4428 (
            .O(N__27066),
            .I(\current_shift_inst.un4_control_input1_29 ));
    Odrv4 I__4427 (
            .O(N__27063),
            .I(\current_shift_inst.un4_control_input1_29 ));
    CascadeMux I__4426 (
            .O(N__27056),
            .I(N__27052));
    InMux I__4425 (
            .O(N__27055),
            .I(N__27048));
    InMux I__4424 (
            .O(N__27052),
            .I(N__27045));
    InMux I__4423 (
            .O(N__27051),
            .I(N__27041));
    LocalMux I__4422 (
            .O(N__27048),
            .I(N__27038));
    LocalMux I__4421 (
            .O(N__27045),
            .I(N__27035));
    InMux I__4420 (
            .O(N__27044),
            .I(N__27032));
    LocalMux I__4419 (
            .O(N__27041),
            .I(N__27029));
    Span4Mux_v I__4418 (
            .O(N__27038),
            .I(N__27022));
    Span4Mux_h I__4417 (
            .O(N__27035),
            .I(N__27022));
    LocalMux I__4416 (
            .O(N__27032),
            .I(N__27022));
    Span4Mux_h I__4415 (
            .O(N__27029),
            .I(N__27019));
    Span4Mux_h I__4414 (
            .O(N__27022),
            .I(N__27016));
    Odrv4 I__4413 (
            .O(N__27019),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv4 I__4412 (
            .O(N__27016),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    InMux I__4411 (
            .O(N__27011),
            .I(N__27006));
    InMux I__4410 (
            .O(N__27010),
            .I(N__27003));
    InMux I__4409 (
            .O(N__27009),
            .I(N__27000));
    LocalMux I__4408 (
            .O(N__27006),
            .I(\current_shift_inst.un4_control_input1_25 ));
    LocalMux I__4407 (
            .O(N__27003),
            .I(\current_shift_inst.un4_control_input1_25 ));
    LocalMux I__4406 (
            .O(N__27000),
            .I(\current_shift_inst.un4_control_input1_25 ));
    InMux I__4405 (
            .O(N__26993),
            .I(N__26989));
    InMux I__4404 (
            .O(N__26992),
            .I(N__26978));
    LocalMux I__4403 (
            .O(N__26989),
            .I(N__26973));
    InMux I__4402 (
            .O(N__26988),
            .I(N__26966));
    InMux I__4401 (
            .O(N__26987),
            .I(N__26966));
    InMux I__4400 (
            .O(N__26986),
            .I(N__26966));
    InMux I__4399 (
            .O(N__26985),
            .I(N__26961));
    InMux I__4398 (
            .O(N__26984),
            .I(N__26958));
    InMux I__4397 (
            .O(N__26983),
            .I(N__26951));
    InMux I__4396 (
            .O(N__26982),
            .I(N__26951));
    InMux I__4395 (
            .O(N__26981),
            .I(N__26951));
    LocalMux I__4394 (
            .O(N__26978),
            .I(N__26948));
    InMux I__4393 (
            .O(N__26977),
            .I(N__26943));
    InMux I__4392 (
            .O(N__26976),
            .I(N__26943));
    Span4Mux_v I__4391 (
            .O(N__26973),
            .I(N__26931));
    LocalMux I__4390 (
            .O(N__26966),
            .I(N__26931));
    InMux I__4389 (
            .O(N__26965),
            .I(N__26926));
    InMux I__4388 (
            .O(N__26964),
            .I(N__26926));
    LocalMux I__4387 (
            .O(N__26961),
            .I(N__26923));
    LocalMux I__4386 (
            .O(N__26958),
            .I(N__26912));
    LocalMux I__4385 (
            .O(N__26951),
            .I(N__26912));
    Span4Mux_h I__4384 (
            .O(N__26948),
            .I(N__26912));
    LocalMux I__4383 (
            .O(N__26943),
            .I(N__26912));
    InMux I__4382 (
            .O(N__26942),
            .I(N__26895));
    InMux I__4381 (
            .O(N__26941),
            .I(N__26895));
    InMux I__4380 (
            .O(N__26940),
            .I(N__26895));
    InMux I__4379 (
            .O(N__26939),
            .I(N__26895));
    InMux I__4378 (
            .O(N__26938),
            .I(N__26895));
    InMux I__4377 (
            .O(N__26937),
            .I(N__26895));
    InMux I__4376 (
            .O(N__26936),
            .I(N__26895));
    Span4Mux_v I__4375 (
            .O(N__26931),
            .I(N__26890));
    LocalMux I__4374 (
            .O(N__26926),
            .I(N__26890));
    Span4Mux_h I__4373 (
            .O(N__26923),
            .I(N__26887));
    InMux I__4372 (
            .O(N__26922),
            .I(N__26884));
    InMux I__4371 (
            .O(N__26921),
            .I(N__26881));
    Span4Mux_v I__4370 (
            .O(N__26912),
            .I(N__26878));
    InMux I__4369 (
            .O(N__26911),
            .I(N__26873));
    InMux I__4368 (
            .O(N__26910),
            .I(N__26873));
    LocalMux I__4367 (
            .O(N__26895),
            .I(N__26866));
    Span4Mux_v I__4366 (
            .O(N__26890),
            .I(N__26866));
    Span4Mux_v I__4365 (
            .O(N__26887),
            .I(N__26866));
    LocalMux I__4364 (
            .O(N__26884),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__4363 (
            .O(N__26881),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__4362 (
            .O(N__26878),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__4361 (
            .O(N__26873),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__4360 (
            .O(N__26866),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    InMux I__4359 (
            .O(N__26855),
            .I(N__26852));
    LocalMux I__4358 (
            .O(N__26852),
            .I(N__26849));
    Span4Mux_v I__4357 (
            .O(N__26849),
            .I(N__26846));
    Odrv4 I__4356 (
            .O(N__26846),
            .I(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ));
    InMux I__4355 (
            .O(N__26843),
            .I(N__26840));
    LocalMux I__4354 (
            .O(N__26840),
            .I(N__26837));
    Odrv12 I__4353 (
            .O(N__26837),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ));
    InMux I__4352 (
            .O(N__26834),
            .I(N__26801));
    InMux I__4351 (
            .O(N__26833),
            .I(N__26801));
    InMux I__4350 (
            .O(N__26832),
            .I(N__26801));
    InMux I__4349 (
            .O(N__26831),
            .I(N__26801));
    InMux I__4348 (
            .O(N__26830),
            .I(N__26801));
    InMux I__4347 (
            .O(N__26829),
            .I(N__26801));
    InMux I__4346 (
            .O(N__26828),
            .I(N__26801));
    InMux I__4345 (
            .O(N__26827),
            .I(N__26801));
    InMux I__4344 (
            .O(N__26826),
            .I(N__26784));
    InMux I__4343 (
            .O(N__26825),
            .I(N__26784));
    InMux I__4342 (
            .O(N__26824),
            .I(N__26784));
    InMux I__4341 (
            .O(N__26823),
            .I(N__26784));
    InMux I__4340 (
            .O(N__26822),
            .I(N__26784));
    InMux I__4339 (
            .O(N__26821),
            .I(N__26784));
    InMux I__4338 (
            .O(N__26820),
            .I(N__26784));
    InMux I__4337 (
            .O(N__26819),
            .I(N__26784));
    InMux I__4336 (
            .O(N__26818),
            .I(N__26781));
    LocalMux I__4335 (
            .O(N__26801),
            .I(N__26775));
    LocalMux I__4334 (
            .O(N__26784),
            .I(N__26775));
    LocalMux I__4333 (
            .O(N__26781),
            .I(N__26772));
    InMux I__4332 (
            .O(N__26780),
            .I(N__26769));
    Span4Mux_s3_h I__4331 (
            .O(N__26775),
            .I(N__26766));
    Span4Mux_v I__4330 (
            .O(N__26772),
            .I(N__26763));
    LocalMux I__4329 (
            .O(N__26769),
            .I(N__26760));
    Span4Mux_v I__4328 (
            .O(N__26766),
            .I(N__26757));
    Span4Mux_h I__4327 (
            .O(N__26763),
            .I(N__26754));
    Span4Mux_s3_h I__4326 (
            .O(N__26760),
            .I(N__26751));
    Span4Mux_h I__4325 (
            .O(N__26757),
            .I(N__26748));
    Span4Mux_v I__4324 (
            .O(N__26754),
            .I(N__26743));
    Span4Mux_h I__4323 (
            .O(N__26751),
            .I(N__26743));
    Odrv4 I__4322 (
            .O(N__26748),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv4 I__4321 (
            .O(N__26743),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    InMux I__4320 (
            .O(N__26738),
            .I(N__26735));
    LocalMux I__4319 (
            .O(N__26735),
            .I(N__26732));
    Odrv4 I__4318 (
            .O(N__26732),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ));
    InMux I__4317 (
            .O(N__26729),
            .I(N__26726));
    LocalMux I__4316 (
            .O(N__26726),
            .I(N__26723));
    Odrv4 I__4315 (
            .O(N__26723),
            .I(\current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ));
    InMux I__4314 (
            .O(N__26720),
            .I(N__26717));
    LocalMux I__4313 (
            .O(N__26717),
            .I(N__26714));
    Odrv4 I__4312 (
            .O(N__26714),
            .I(\current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ));
    InMux I__4311 (
            .O(N__26711),
            .I(N__26708));
    LocalMux I__4310 (
            .O(N__26708),
            .I(N__26705));
    Odrv4 I__4309 (
            .O(N__26705),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ));
    CascadeMux I__4308 (
            .O(N__26702),
            .I(N__26699));
    InMux I__4307 (
            .O(N__26699),
            .I(N__26696));
    LocalMux I__4306 (
            .O(N__26696),
            .I(N__26693));
    Span4Mux_v I__4305 (
            .O(N__26693),
            .I(N__26690));
    Odrv4 I__4304 (
            .O(N__26690),
            .I(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ));
    CascadeMux I__4303 (
            .O(N__26687),
            .I(N__26684));
    InMux I__4302 (
            .O(N__26684),
            .I(N__26681));
    LocalMux I__4301 (
            .O(N__26681),
            .I(N__26678));
    Span4Mux_v I__4300 (
            .O(N__26678),
            .I(N__26675));
    Odrv4 I__4299 (
            .O(N__26675),
            .I(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ));
    CascadeMux I__4298 (
            .O(N__26672),
            .I(N__26669));
    InMux I__4297 (
            .O(N__26669),
            .I(N__26666));
    LocalMux I__4296 (
            .O(N__26666),
            .I(N__26663));
    Odrv4 I__4295 (
            .O(N__26663),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ));
    InMux I__4294 (
            .O(N__26660),
            .I(N__26657));
    LocalMux I__4293 (
            .O(N__26657),
            .I(N__26654));
    Span4Mux_h I__4292 (
            .O(N__26654),
            .I(N__26651));
    Odrv4 I__4291 (
            .O(N__26651),
            .I(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ));
    CascadeMux I__4290 (
            .O(N__26648),
            .I(N__26644));
    InMux I__4289 (
            .O(N__26647),
            .I(N__26639));
    InMux I__4288 (
            .O(N__26644),
            .I(N__26636));
    InMux I__4287 (
            .O(N__26643),
            .I(N__26633));
    InMux I__4286 (
            .O(N__26642),
            .I(N__26630));
    LocalMux I__4285 (
            .O(N__26639),
            .I(N__26625));
    LocalMux I__4284 (
            .O(N__26636),
            .I(N__26625));
    LocalMux I__4283 (
            .O(N__26633),
            .I(N__26620));
    LocalMux I__4282 (
            .O(N__26630),
            .I(N__26620));
    Span4Mux_v I__4281 (
            .O(N__26625),
            .I(N__26617));
    Span4Mux_v I__4280 (
            .O(N__26620),
            .I(N__26614));
    Odrv4 I__4279 (
            .O(N__26617),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    Odrv4 I__4278 (
            .O(N__26614),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    CascadeMux I__4277 (
            .O(N__26609),
            .I(N__26606));
    InMux I__4276 (
            .O(N__26606),
            .I(N__26599));
    InMux I__4275 (
            .O(N__26605),
            .I(N__26599));
    InMux I__4274 (
            .O(N__26604),
            .I(N__26596));
    LocalMux I__4273 (
            .O(N__26599),
            .I(\current_shift_inst.un4_control_input1_27 ));
    LocalMux I__4272 (
            .O(N__26596),
            .I(\current_shift_inst.un4_control_input1_27 ));
    InMux I__4271 (
            .O(N__26591),
            .I(\current_shift_inst.un38_control_input_cry_28_s1 ));
    CascadeMux I__4270 (
            .O(N__26588),
            .I(N__26585));
    InMux I__4269 (
            .O(N__26585),
            .I(N__26582));
    LocalMux I__4268 (
            .O(N__26582),
            .I(N__26579));
    Span4Mux_h I__4267 (
            .O(N__26579),
            .I(N__26576));
    Odrv4 I__4266 (
            .O(N__26576),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ));
    InMux I__4265 (
            .O(N__26573),
            .I(\current_shift_inst.un38_control_input_cry_29_s1 ));
    InMux I__4264 (
            .O(N__26570),
            .I(\current_shift_inst.un38_control_input_cry_30_s1 ));
    CascadeMux I__4263 (
            .O(N__26567),
            .I(N__26563));
    CascadeMux I__4262 (
            .O(N__26566),
            .I(N__26560));
    InMux I__4261 (
            .O(N__26563),
            .I(N__26557));
    InMux I__4260 (
            .O(N__26560),
            .I(N__26554));
    LocalMux I__4259 (
            .O(N__26557),
            .I(N__26551));
    LocalMux I__4258 (
            .O(N__26554),
            .I(N__26546));
    Span4Mux_v I__4257 (
            .O(N__26551),
            .I(N__26543));
    InMux I__4256 (
            .O(N__26550),
            .I(N__26538));
    InMux I__4255 (
            .O(N__26549),
            .I(N__26538));
    Span4Mux_h I__4254 (
            .O(N__26546),
            .I(N__26531));
    Span4Mux_h I__4253 (
            .O(N__26543),
            .I(N__26531));
    LocalMux I__4252 (
            .O(N__26538),
            .I(N__26531));
    Odrv4 I__4251 (
            .O(N__26531),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    InMux I__4250 (
            .O(N__26528),
            .I(N__26523));
    InMux I__4249 (
            .O(N__26527),
            .I(N__26520));
    InMux I__4248 (
            .O(N__26526),
            .I(N__26517));
    LocalMux I__4247 (
            .O(N__26523),
            .I(N__26514));
    LocalMux I__4246 (
            .O(N__26520),
            .I(\current_shift_inst.un4_control_input1_9 ));
    LocalMux I__4245 (
            .O(N__26517),
            .I(\current_shift_inst.un4_control_input1_9 ));
    Odrv4 I__4244 (
            .O(N__26514),
            .I(\current_shift_inst.un4_control_input1_9 ));
    CascadeMux I__4243 (
            .O(N__26507),
            .I(N__26504));
    InMux I__4242 (
            .O(N__26504),
            .I(N__26501));
    LocalMux I__4241 (
            .O(N__26501),
            .I(N__26498));
    Odrv4 I__4240 (
            .O(N__26498),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ));
    InMux I__4239 (
            .O(N__26495),
            .I(N__26492));
    LocalMux I__4238 (
            .O(N__26492),
            .I(\current_shift_inst.un4_control_input_1_axb_11 ));
    InMux I__4237 (
            .O(N__26489),
            .I(N__26486));
    LocalMux I__4236 (
            .O(N__26486),
            .I(\current_shift_inst.un4_control_input_1_axb_14 ));
    CascadeMux I__4235 (
            .O(N__26483),
            .I(N__26480));
    InMux I__4234 (
            .O(N__26480),
            .I(N__26477));
    LocalMux I__4233 (
            .O(N__26477),
            .I(N__26474));
    Odrv4 I__4232 (
            .O(N__26474),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ));
    InMux I__4231 (
            .O(N__26471),
            .I(N__26468));
    LocalMux I__4230 (
            .O(N__26468),
            .I(N__26465));
    Odrv4 I__4229 (
            .O(N__26465),
            .I(\current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ));
    CascadeMux I__4228 (
            .O(N__26462),
            .I(N__26459));
    InMux I__4227 (
            .O(N__26459),
            .I(N__26456));
    LocalMux I__4226 (
            .O(N__26456),
            .I(N__26453));
    Odrv12 I__4225 (
            .O(N__26453),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ));
    InMux I__4224 (
            .O(N__26450),
            .I(N__26447));
    LocalMux I__4223 (
            .O(N__26447),
            .I(N__26444));
    Span4Mux_h I__4222 (
            .O(N__26444),
            .I(N__26441));
    Odrv4 I__4221 (
            .O(N__26441),
            .I(\current_shift_inst.un38_control_input_0_s1_21 ));
    InMux I__4220 (
            .O(N__26438),
            .I(\current_shift_inst.un38_control_input_cry_20_s1 ));
    InMux I__4219 (
            .O(N__26435),
            .I(N__26432));
    LocalMux I__4218 (
            .O(N__26432),
            .I(N__26429));
    Span4Mux_v I__4217 (
            .O(N__26429),
            .I(N__26426));
    Odrv4 I__4216 (
            .O(N__26426),
            .I(\current_shift_inst.un38_control_input_0_s1_22 ));
    InMux I__4215 (
            .O(N__26423),
            .I(\current_shift_inst.un38_control_input_cry_21_s1 ));
    InMux I__4214 (
            .O(N__26420),
            .I(N__26417));
    LocalMux I__4213 (
            .O(N__26417),
            .I(N__26414));
    Span4Mux_h I__4212 (
            .O(N__26414),
            .I(N__26411));
    Odrv4 I__4211 (
            .O(N__26411),
            .I(\current_shift_inst.un38_control_input_0_s1_23 ));
    InMux I__4210 (
            .O(N__26408),
            .I(\current_shift_inst.un38_control_input_cry_22_s1 ));
    InMux I__4209 (
            .O(N__26405),
            .I(N__26402));
    LocalMux I__4208 (
            .O(N__26402),
            .I(N__26399));
    Span4Mux_h I__4207 (
            .O(N__26399),
            .I(N__26396));
    Odrv4 I__4206 (
            .O(N__26396),
            .I(\current_shift_inst.un38_control_input_0_s1_24 ));
    InMux I__4205 (
            .O(N__26393),
            .I(bfn_11_18_0_));
    InMux I__4204 (
            .O(N__26390),
            .I(N__26387));
    LocalMux I__4203 (
            .O(N__26387),
            .I(N__26384));
    Span4Mux_h I__4202 (
            .O(N__26384),
            .I(N__26381));
    Odrv4 I__4201 (
            .O(N__26381),
            .I(\current_shift_inst.un38_control_input_0_s1_25 ));
    InMux I__4200 (
            .O(N__26378),
            .I(\current_shift_inst.un38_control_input_cry_24_s1 ));
    InMux I__4199 (
            .O(N__26375),
            .I(N__26372));
    LocalMux I__4198 (
            .O(N__26372),
            .I(N__26369));
    Span4Mux_h I__4197 (
            .O(N__26369),
            .I(N__26366));
    Odrv4 I__4196 (
            .O(N__26366),
            .I(\current_shift_inst.un38_control_input_0_s1_26 ));
    InMux I__4195 (
            .O(N__26363),
            .I(\current_shift_inst.un38_control_input_cry_25_s1 ));
    InMux I__4194 (
            .O(N__26360),
            .I(N__26357));
    LocalMux I__4193 (
            .O(N__26357),
            .I(N__26354));
    Span4Mux_h I__4192 (
            .O(N__26354),
            .I(N__26351));
    Odrv4 I__4191 (
            .O(N__26351),
            .I(\current_shift_inst.un38_control_input_0_s1_27 ));
    InMux I__4190 (
            .O(N__26348),
            .I(\current_shift_inst.un38_control_input_cry_26_s1 ));
    InMux I__4189 (
            .O(N__26345),
            .I(\current_shift_inst.un38_control_input_cry_27_s1 ));
    InMux I__4188 (
            .O(N__26342),
            .I(N__26339));
    LocalMux I__4187 (
            .O(N__26339),
            .I(\current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ));
    CascadeMux I__4186 (
            .O(N__26336),
            .I(N__26333));
    InMux I__4185 (
            .O(N__26333),
            .I(N__26330));
    LocalMux I__4184 (
            .O(N__26330),
            .I(\current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ));
    CascadeMux I__4183 (
            .O(N__26327),
            .I(N__26324));
    InMux I__4182 (
            .O(N__26324),
            .I(N__26321));
    LocalMux I__4181 (
            .O(N__26321),
            .I(N__26318));
    Span4Mux_v I__4180 (
            .O(N__26318),
            .I(N__26315));
    Odrv4 I__4179 (
            .O(N__26315),
            .I(\current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ));
    InMux I__4178 (
            .O(N__26312),
            .I(N__26309));
    LocalMux I__4177 (
            .O(N__26309),
            .I(N__26306));
    Odrv4 I__4176 (
            .O(N__26306),
            .I(\current_shift_inst.un38_control_input_0_s1_20 ));
    InMux I__4175 (
            .O(N__26303),
            .I(\current_shift_inst.un38_control_input_cry_19_s1 ));
    InMux I__4174 (
            .O(N__26300),
            .I(N__26297));
    LocalMux I__4173 (
            .O(N__26297),
            .I(\current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ));
    CascadeMux I__4172 (
            .O(N__26294),
            .I(N__26291));
    InMux I__4171 (
            .O(N__26291),
            .I(N__26288));
    LocalMux I__4170 (
            .O(N__26288),
            .I(\current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ));
    InMux I__4169 (
            .O(N__26285),
            .I(N__26282));
    LocalMux I__4168 (
            .O(N__26282),
            .I(\current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ));
    CascadeMux I__4167 (
            .O(N__26279),
            .I(N__26276));
    InMux I__4166 (
            .O(N__26276),
            .I(N__26273));
    LocalMux I__4165 (
            .O(N__26273),
            .I(\current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ));
    InMux I__4164 (
            .O(N__26270),
            .I(N__26267));
    LocalMux I__4163 (
            .O(N__26267),
            .I(\current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ));
    CascadeMux I__4162 (
            .O(N__26264),
            .I(N__26261));
    InMux I__4161 (
            .O(N__26261),
            .I(N__26258));
    LocalMux I__4160 (
            .O(N__26258),
            .I(\current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ));
    CascadeMux I__4159 (
            .O(N__26255),
            .I(N__26252));
    InMux I__4158 (
            .O(N__26252),
            .I(N__26249));
    LocalMux I__4157 (
            .O(N__26249),
            .I(\current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ));
    InMux I__4156 (
            .O(N__26246),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ));
    InMux I__4155 (
            .O(N__26243),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ));
    InMux I__4154 (
            .O(N__26240),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ));
    CascadeMux I__4153 (
            .O(N__26237),
            .I(N__26233));
    CascadeMux I__4152 (
            .O(N__26236),
            .I(N__26229));
    InMux I__4151 (
            .O(N__26233),
            .I(N__26222));
    InMux I__4150 (
            .O(N__26232),
            .I(N__26222));
    InMux I__4149 (
            .O(N__26229),
            .I(N__26222));
    LocalMux I__4148 (
            .O(N__26222),
            .I(N__26218));
    InMux I__4147 (
            .O(N__26221),
            .I(N__26215));
    Sp12to4 I__4146 (
            .O(N__26218),
            .I(N__26212));
    LocalMux I__4145 (
            .O(N__26215),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    Odrv12 I__4144 (
            .O(N__26212),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    InMux I__4143 (
            .O(N__26207),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ));
    IoInMux I__4142 (
            .O(N__26204),
            .I(N__26189));
    InMux I__4141 (
            .O(N__26203),
            .I(N__26186));
    InMux I__4140 (
            .O(N__26202),
            .I(N__26177));
    InMux I__4139 (
            .O(N__26201),
            .I(N__26177));
    InMux I__4138 (
            .O(N__26200),
            .I(N__26177));
    InMux I__4137 (
            .O(N__26199),
            .I(N__26177));
    InMux I__4136 (
            .O(N__26198),
            .I(N__26170));
    InMux I__4135 (
            .O(N__26197),
            .I(N__26170));
    InMux I__4134 (
            .O(N__26196),
            .I(N__26170));
    InMux I__4133 (
            .O(N__26195),
            .I(N__26161));
    InMux I__4132 (
            .O(N__26194),
            .I(N__26161));
    InMux I__4131 (
            .O(N__26193),
            .I(N__26161));
    InMux I__4130 (
            .O(N__26192),
            .I(N__26161));
    LocalMux I__4129 (
            .O(N__26189),
            .I(N__26139));
    LocalMux I__4128 (
            .O(N__26186),
            .I(N__26130));
    LocalMux I__4127 (
            .O(N__26177),
            .I(N__26130));
    LocalMux I__4126 (
            .O(N__26170),
            .I(N__26130));
    LocalMux I__4125 (
            .O(N__26161),
            .I(N__26130));
    InMux I__4124 (
            .O(N__26160),
            .I(N__26121));
    InMux I__4123 (
            .O(N__26159),
            .I(N__26121));
    InMux I__4122 (
            .O(N__26158),
            .I(N__26121));
    InMux I__4121 (
            .O(N__26157),
            .I(N__26121));
    InMux I__4120 (
            .O(N__26156),
            .I(N__26112));
    InMux I__4119 (
            .O(N__26155),
            .I(N__26112));
    InMux I__4118 (
            .O(N__26154),
            .I(N__26112));
    InMux I__4117 (
            .O(N__26153),
            .I(N__26112));
    InMux I__4116 (
            .O(N__26152),
            .I(N__26103));
    InMux I__4115 (
            .O(N__26151),
            .I(N__26103));
    InMux I__4114 (
            .O(N__26150),
            .I(N__26103));
    InMux I__4113 (
            .O(N__26149),
            .I(N__26103));
    InMux I__4112 (
            .O(N__26148),
            .I(N__26094));
    InMux I__4111 (
            .O(N__26147),
            .I(N__26094));
    InMux I__4110 (
            .O(N__26146),
            .I(N__26094));
    InMux I__4109 (
            .O(N__26145),
            .I(N__26094));
    InMux I__4108 (
            .O(N__26144),
            .I(N__26087));
    InMux I__4107 (
            .O(N__26143),
            .I(N__26087));
    InMux I__4106 (
            .O(N__26142),
            .I(N__26087));
    Span4Mux_s0_v I__4105 (
            .O(N__26139),
            .I(N__26084));
    Span4Mux_v I__4104 (
            .O(N__26130),
            .I(N__26081));
    LocalMux I__4103 (
            .O(N__26121),
            .I(N__26070));
    LocalMux I__4102 (
            .O(N__26112),
            .I(N__26070));
    LocalMux I__4101 (
            .O(N__26103),
            .I(N__26070));
    LocalMux I__4100 (
            .O(N__26094),
            .I(N__26070));
    LocalMux I__4099 (
            .O(N__26087),
            .I(N__26070));
    Sp12to4 I__4098 (
            .O(N__26084),
            .I(N__26067));
    Span4Mux_h I__4097 (
            .O(N__26081),
            .I(N__26062));
    Span4Mux_v I__4096 (
            .O(N__26070),
            .I(N__26062));
    Span12Mux_s5_h I__4095 (
            .O(N__26067),
            .I(N__26059));
    Span4Mux_h I__4094 (
            .O(N__26062),
            .I(N__26056));
    Span12Mux_v I__4093 (
            .O(N__26059),
            .I(N__26053));
    Odrv4 I__4092 (
            .O(N__26056),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv12 I__4091 (
            .O(N__26053),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    InMux I__4090 (
            .O(N__26048),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ));
    CascadeMux I__4089 (
            .O(N__26045),
            .I(N__26041));
    InMux I__4088 (
            .O(N__26044),
            .I(N__26033));
    InMux I__4087 (
            .O(N__26041),
            .I(N__26033));
    InMux I__4086 (
            .O(N__26040),
            .I(N__26033));
    LocalMux I__4085 (
            .O(N__26033),
            .I(N__26029));
    InMux I__4084 (
            .O(N__26032),
            .I(N__26026));
    Span4Mux_h I__4083 (
            .O(N__26029),
            .I(N__26023));
    LocalMux I__4082 (
            .O(N__26026),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    Odrv4 I__4081 (
            .O(N__26023),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    CascadeMux I__4080 (
            .O(N__26018),
            .I(N__26015));
    InMux I__4079 (
            .O(N__26015),
            .I(N__26012));
    LocalMux I__4078 (
            .O(N__26012),
            .I(N__26009));
    Odrv4 I__4077 (
            .O(N__26009),
            .I(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ));
    CascadeMux I__4076 (
            .O(N__26006),
            .I(N__26003));
    InMux I__4075 (
            .O(N__26003),
            .I(N__26000));
    LocalMux I__4074 (
            .O(N__26000),
            .I(\current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ));
    CascadeMux I__4073 (
            .O(N__25997),
            .I(N__25993));
    CascadeMux I__4072 (
            .O(N__25996),
            .I(N__25990));
    InMux I__4071 (
            .O(N__25993),
            .I(N__25987));
    InMux I__4070 (
            .O(N__25990),
            .I(N__25984));
    LocalMux I__4069 (
            .O(N__25987),
            .I(N__25978));
    LocalMux I__4068 (
            .O(N__25984),
            .I(N__25978));
    InMux I__4067 (
            .O(N__25983),
            .I(N__25975));
    Span4Mux_h I__4066 (
            .O(N__25978),
            .I(N__25972));
    LocalMux I__4065 (
            .O(N__25975),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv4 I__4064 (
            .O(N__25972),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__4063 (
            .O(N__25967),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ));
    InMux I__4062 (
            .O(N__25964),
            .I(N__25960));
    InMux I__4061 (
            .O(N__25963),
            .I(N__25957));
    LocalMux I__4060 (
            .O(N__25960),
            .I(N__25951));
    LocalMux I__4059 (
            .O(N__25957),
            .I(N__25951));
    InMux I__4058 (
            .O(N__25956),
            .I(N__25948));
    Span4Mux_h I__4057 (
            .O(N__25951),
            .I(N__25945));
    LocalMux I__4056 (
            .O(N__25948),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv4 I__4055 (
            .O(N__25945),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__4054 (
            .O(N__25940),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ));
    InMux I__4053 (
            .O(N__25937),
            .I(N__25931));
    InMux I__4052 (
            .O(N__25936),
            .I(N__25931));
    LocalMux I__4051 (
            .O(N__25931),
            .I(N__25927));
    InMux I__4050 (
            .O(N__25930),
            .I(N__25924));
    Span4Mux_h I__4049 (
            .O(N__25927),
            .I(N__25921));
    LocalMux I__4048 (
            .O(N__25924),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ));
    Odrv4 I__4047 (
            .O(N__25921),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ));
    InMux I__4046 (
            .O(N__25916),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ));
    CascadeMux I__4045 (
            .O(N__25913),
            .I(N__25909));
    InMux I__4044 (
            .O(N__25912),
            .I(N__25904));
    InMux I__4043 (
            .O(N__25909),
            .I(N__25904));
    LocalMux I__4042 (
            .O(N__25904),
            .I(N__25900));
    InMux I__4041 (
            .O(N__25903),
            .I(N__25897));
    Span4Mux_v I__4040 (
            .O(N__25900),
            .I(N__25894));
    LocalMux I__4039 (
            .O(N__25897),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ));
    Odrv4 I__4038 (
            .O(N__25894),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ));
    InMux I__4037 (
            .O(N__25889),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ));
    CascadeMux I__4036 (
            .O(N__25886),
            .I(N__25882));
    InMux I__4035 (
            .O(N__25885),
            .I(N__25877));
    InMux I__4034 (
            .O(N__25882),
            .I(N__25877));
    LocalMux I__4033 (
            .O(N__25877),
            .I(N__25873));
    InMux I__4032 (
            .O(N__25876),
            .I(N__25870));
    Span4Mux_h I__4031 (
            .O(N__25873),
            .I(N__25867));
    LocalMux I__4030 (
            .O(N__25870),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ));
    Odrv4 I__4029 (
            .O(N__25867),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ));
    InMux I__4028 (
            .O(N__25862),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ));
    InMux I__4027 (
            .O(N__25859),
            .I(N__25853));
    InMux I__4026 (
            .O(N__25858),
            .I(N__25853));
    LocalMux I__4025 (
            .O(N__25853),
            .I(N__25849));
    InMux I__4024 (
            .O(N__25852),
            .I(N__25846));
    Span4Mux_v I__4023 (
            .O(N__25849),
            .I(N__25843));
    LocalMux I__4022 (
            .O(N__25846),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ));
    Odrv4 I__4021 (
            .O(N__25843),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ));
    InMux I__4020 (
            .O(N__25838),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ));
    InMux I__4019 (
            .O(N__25835),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ));
    InMux I__4018 (
            .O(N__25832),
            .I(bfn_11_14_0_));
    InMux I__4017 (
            .O(N__25829),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ));
    InMux I__4016 (
            .O(N__25826),
            .I(N__25822));
    InMux I__4015 (
            .O(N__25825),
            .I(N__25819));
    LocalMux I__4014 (
            .O(N__25822),
            .I(N__25816));
    LocalMux I__4013 (
            .O(N__25819),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    Odrv4 I__4012 (
            .O(N__25816),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__4011 (
            .O(N__25811),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__4010 (
            .O(N__25808),
            .I(N__25804));
    InMux I__4009 (
            .O(N__25807),
            .I(N__25801));
    LocalMux I__4008 (
            .O(N__25804),
            .I(N__25798));
    LocalMux I__4007 (
            .O(N__25801),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    Odrv12 I__4006 (
            .O(N__25798),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__4005 (
            .O(N__25793),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__4004 (
            .O(N__25790),
            .I(N__25786));
    InMux I__4003 (
            .O(N__25789),
            .I(N__25783));
    LocalMux I__4002 (
            .O(N__25786),
            .I(N__25780));
    LocalMux I__4001 (
            .O(N__25783),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__4000 (
            .O(N__25780),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__3999 (
            .O(N__25775),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__3998 (
            .O(N__25772),
            .I(N__25768));
    InMux I__3997 (
            .O(N__25771),
            .I(N__25765));
    LocalMux I__3996 (
            .O(N__25768),
            .I(N__25762));
    LocalMux I__3995 (
            .O(N__25765),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    Odrv12 I__3994 (
            .O(N__25762),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__3993 (
            .O(N__25757),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__3992 (
            .O(N__25754),
            .I(N__25750));
    InMux I__3991 (
            .O(N__25753),
            .I(N__25747));
    LocalMux I__3990 (
            .O(N__25750),
            .I(N__25744));
    LocalMux I__3989 (
            .O(N__25747),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    Odrv12 I__3988 (
            .O(N__25744),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__3987 (
            .O(N__25739),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__3986 (
            .O(N__25736),
            .I(N__25732));
    InMux I__3985 (
            .O(N__25735),
            .I(N__25729));
    LocalMux I__3984 (
            .O(N__25732),
            .I(N__25726));
    LocalMux I__3983 (
            .O(N__25729),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv4 I__3982 (
            .O(N__25726),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__3981 (
            .O(N__25721),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ));
    InMux I__3980 (
            .O(N__25718),
            .I(N__25713));
    InMux I__3979 (
            .O(N__25717),
            .I(N__25708));
    InMux I__3978 (
            .O(N__25716),
            .I(N__25708));
    LocalMux I__3977 (
            .O(N__25713),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    LocalMux I__3976 (
            .O(N__25708),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__3975 (
            .O(N__25703),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ));
    InMux I__3974 (
            .O(N__25700),
            .I(N__25695));
    InMux I__3973 (
            .O(N__25699),
            .I(N__25690));
    InMux I__3972 (
            .O(N__25698),
            .I(N__25690));
    LocalMux I__3971 (
            .O(N__25695),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    LocalMux I__3970 (
            .O(N__25690),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__3969 (
            .O(N__25685),
            .I(bfn_11_13_0_));
    InMux I__3968 (
            .O(N__25682),
            .I(N__25678));
    InMux I__3967 (
            .O(N__25681),
            .I(N__25675));
    LocalMux I__3966 (
            .O(N__25678),
            .I(N__25672));
    LocalMux I__3965 (
            .O(N__25675),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    Odrv4 I__3964 (
            .O(N__25672),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__3963 (
            .O(N__25667),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ));
    CascadeMux I__3962 (
            .O(N__25664),
            .I(N__25661));
    InMux I__3961 (
            .O(N__25661),
            .I(N__25658));
    LocalMux I__3960 (
            .O(N__25658),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28 ));
    InMux I__3959 (
            .O(N__25655),
            .I(N__25651));
    InMux I__3958 (
            .O(N__25654),
            .I(N__25648));
    LocalMux I__3957 (
            .O(N__25651),
            .I(N__25645));
    LocalMux I__3956 (
            .O(N__25648),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    Odrv4 I__3955 (
            .O(N__25645),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__3954 (
            .O(N__25640),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__3953 (
            .O(N__25637),
            .I(N__25634));
    LocalMux I__3952 (
            .O(N__25634),
            .I(N__25630));
    InMux I__3951 (
            .O(N__25633),
            .I(N__25627));
    Span4Mux_h I__3950 (
            .O(N__25630),
            .I(N__25624));
    LocalMux I__3949 (
            .O(N__25627),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    Odrv4 I__3948 (
            .O(N__25624),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__3947 (
            .O(N__25619),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__3946 (
            .O(N__25616),
            .I(N__25612));
    InMux I__3945 (
            .O(N__25615),
            .I(N__25609));
    LocalMux I__3944 (
            .O(N__25612),
            .I(N__25606));
    LocalMux I__3943 (
            .O(N__25609),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    Odrv4 I__3942 (
            .O(N__25606),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__3941 (
            .O(N__25601),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__3940 (
            .O(N__25598),
            .I(N__25594));
    InMux I__3939 (
            .O(N__25597),
            .I(N__25591));
    LocalMux I__3938 (
            .O(N__25594),
            .I(N__25588));
    LocalMux I__3937 (
            .O(N__25591),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    Odrv12 I__3936 (
            .O(N__25588),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__3935 (
            .O(N__25583),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__3934 (
            .O(N__25580),
            .I(N__25577));
    LocalMux I__3933 (
            .O(N__25577),
            .I(N__25573));
    InMux I__3932 (
            .O(N__25576),
            .I(N__25570));
    Span4Mux_h I__3931 (
            .O(N__25573),
            .I(N__25567));
    LocalMux I__3930 (
            .O(N__25570),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    Odrv4 I__3929 (
            .O(N__25567),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__3928 (
            .O(N__25562),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__3927 (
            .O(N__25559),
            .I(N__25555));
    InMux I__3926 (
            .O(N__25558),
            .I(N__25552));
    LocalMux I__3925 (
            .O(N__25555),
            .I(N__25549));
    LocalMux I__3924 (
            .O(N__25552),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    Odrv4 I__3923 (
            .O(N__25549),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__3922 (
            .O(N__25544),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__3921 (
            .O(N__25541),
            .I(N__25537));
    InMux I__3920 (
            .O(N__25540),
            .I(N__25534));
    LocalMux I__3919 (
            .O(N__25537),
            .I(N__25531));
    LocalMux I__3918 (
            .O(N__25534),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    Odrv4 I__3917 (
            .O(N__25531),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__3916 (
            .O(N__25526),
            .I(bfn_11_12_0_));
    InMux I__3915 (
            .O(N__25523),
            .I(N__25520));
    LocalMux I__3914 (
            .O(N__25520),
            .I(N__25517));
    Span4Mux_v I__3913 (
            .O(N__25517),
            .I(N__25514));
    Odrv4 I__3912 (
            .O(N__25514),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ));
    CascadeMux I__3911 (
            .O(N__25511),
            .I(N__25508));
    InMux I__3910 (
            .O(N__25508),
            .I(N__25505));
    LocalMux I__3909 (
            .O(N__25505),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt24 ));
    InMux I__3908 (
            .O(N__25502),
            .I(N__25499));
    LocalMux I__3907 (
            .O(N__25499),
            .I(N__25496));
    Odrv12 I__3906 (
            .O(N__25496),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt26 ));
    CascadeMux I__3905 (
            .O(N__25493),
            .I(N__25490));
    InMux I__3904 (
            .O(N__25490),
            .I(N__25487));
    LocalMux I__3903 (
            .O(N__25487),
            .I(N__25484));
    Span4Mux_v I__3902 (
            .O(N__25484),
            .I(N__25481));
    Odrv4 I__3901 (
            .O(N__25481),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ));
    InMux I__3900 (
            .O(N__25478),
            .I(N__25475));
    LocalMux I__3899 (
            .O(N__25475),
            .I(N__25472));
    Odrv4 I__3898 (
            .O(N__25472),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ));
    CascadeMux I__3897 (
            .O(N__25469),
            .I(N__25466));
    InMux I__3896 (
            .O(N__25466),
            .I(N__25463));
    LocalMux I__3895 (
            .O(N__25463),
            .I(N__25460));
    Span4Mux_v I__3894 (
            .O(N__25460),
            .I(N__25456));
    InMux I__3893 (
            .O(N__25459),
            .I(N__25453));
    Odrv4 I__3892 (
            .O(N__25456),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt30 ));
    LocalMux I__3891 (
            .O(N__25453),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt30 ));
    InMux I__3890 (
            .O(N__25448),
            .I(N__25445));
    LocalMux I__3889 (
            .O(N__25445),
            .I(N__25442));
    Odrv12 I__3888 (
            .O(N__25442),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO ));
    InMux I__3887 (
            .O(N__25439),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ));
    InMux I__3886 (
            .O(N__25436),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30 ));
    InMux I__3885 (
            .O(N__25433),
            .I(N__25430));
    LocalMux I__3884 (
            .O(N__25430),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt28 ));
    InMux I__3883 (
            .O(N__25427),
            .I(N__25424));
    LocalMux I__3882 (
            .O(N__25424),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ));
    CascadeMux I__3881 (
            .O(N__25421),
            .I(N__25417));
    InMux I__3880 (
            .O(N__25420),
            .I(N__25413));
    InMux I__3879 (
            .O(N__25417),
            .I(N__25410));
    InMux I__3878 (
            .O(N__25416),
            .I(N__25407));
    LocalMux I__3877 (
            .O(N__25413),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__3876 (
            .O(N__25410),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__3875 (
            .O(N__25407),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__3874 (
            .O(N__25400),
            .I(N__25397));
    LocalMux I__3873 (
            .O(N__25397),
            .I(N__25394));
    Span4Mux_h I__3872 (
            .O(N__25394),
            .I(N__25391));
    Odrv4 I__3871 (
            .O(N__25391),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ));
    CascadeMux I__3870 (
            .O(N__25388),
            .I(N__25385));
    InMux I__3869 (
            .O(N__25385),
            .I(N__25382));
    LocalMux I__3868 (
            .O(N__25382),
            .I(N__25379));
    Odrv4 I__3867 (
            .O(N__25379),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    InMux I__3866 (
            .O(N__25376),
            .I(N__25373));
    LocalMux I__3865 (
            .O(N__25373),
            .I(N__25370));
    Span4Mux_h I__3864 (
            .O(N__25370),
            .I(N__25367));
    Odrv4 I__3863 (
            .O(N__25367),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ));
    CascadeMux I__3862 (
            .O(N__25364),
            .I(N__25361));
    InMux I__3861 (
            .O(N__25361),
            .I(N__25358));
    LocalMux I__3860 (
            .O(N__25358),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    CascadeMux I__3859 (
            .O(N__25355),
            .I(N__25352));
    InMux I__3858 (
            .O(N__25352),
            .I(N__25349));
    LocalMux I__3857 (
            .O(N__25349),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    CascadeMux I__3856 (
            .O(N__25346),
            .I(N__25343));
    InMux I__3855 (
            .O(N__25343),
            .I(N__25340));
    LocalMux I__3854 (
            .O(N__25340),
            .I(N__25337));
    Span4Mux_v I__3853 (
            .O(N__25337),
            .I(N__25334));
    Odrv4 I__3852 (
            .O(N__25334),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ));
    InMux I__3851 (
            .O(N__25331),
            .I(N__25328));
    LocalMux I__3850 (
            .O(N__25328),
            .I(N__25325));
    Odrv4 I__3849 (
            .O(N__25325),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    InMux I__3848 (
            .O(N__25322),
            .I(N__25319));
    LocalMux I__3847 (
            .O(N__25319),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ));
    CascadeMux I__3846 (
            .O(N__25316),
            .I(N__25313));
    InMux I__3845 (
            .O(N__25313),
            .I(N__25310));
    LocalMux I__3844 (
            .O(N__25310),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt18 ));
    InMux I__3843 (
            .O(N__25307),
            .I(N__25304));
    LocalMux I__3842 (
            .O(N__25304),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ));
    CascadeMux I__3841 (
            .O(N__25301),
            .I(N__25298));
    InMux I__3840 (
            .O(N__25298),
            .I(N__25295));
    LocalMux I__3839 (
            .O(N__25295),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    CascadeMux I__3838 (
            .O(N__25292),
            .I(N__25289));
    InMux I__3837 (
            .O(N__25289),
            .I(N__25286));
    LocalMux I__3836 (
            .O(N__25286),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ));
    InMux I__3835 (
            .O(N__25283),
            .I(N__25280));
    LocalMux I__3834 (
            .O(N__25280),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    InMux I__3833 (
            .O(N__25277),
            .I(N__25274));
    LocalMux I__3832 (
            .O(N__25274),
            .I(N__25271));
    Odrv4 I__3831 (
            .O(N__25271),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ));
    CascadeMux I__3830 (
            .O(N__25268),
            .I(N__25265));
    InMux I__3829 (
            .O(N__25265),
            .I(N__25262));
    LocalMux I__3828 (
            .O(N__25262),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    InMux I__3827 (
            .O(N__25259),
            .I(N__25256));
    LocalMux I__3826 (
            .O(N__25256),
            .I(N__25253));
    Odrv4 I__3825 (
            .O(N__25253),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ));
    CascadeMux I__3824 (
            .O(N__25250),
            .I(N__25247));
    InMux I__3823 (
            .O(N__25247),
            .I(N__25244));
    LocalMux I__3822 (
            .O(N__25244),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    CascadeMux I__3821 (
            .O(N__25241),
            .I(N__25238));
    InMux I__3820 (
            .O(N__25238),
            .I(N__25235));
    LocalMux I__3819 (
            .O(N__25235),
            .I(N__25232));
    Odrv4 I__3818 (
            .O(N__25232),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ));
    InMux I__3817 (
            .O(N__25229),
            .I(N__25226));
    LocalMux I__3816 (
            .O(N__25226),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    InMux I__3815 (
            .O(N__25223),
            .I(N__25220));
    LocalMux I__3814 (
            .O(N__25220),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ));
    CascadeMux I__3813 (
            .O(N__25217),
            .I(N__25214));
    InMux I__3812 (
            .O(N__25214),
            .I(N__25211));
    LocalMux I__3811 (
            .O(N__25211),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    InMux I__3810 (
            .O(N__25208),
            .I(N__25205));
    LocalMux I__3809 (
            .O(N__25205),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ));
    CascadeMux I__3808 (
            .O(N__25202),
            .I(N__25199));
    InMux I__3807 (
            .O(N__25199),
            .I(N__25196));
    LocalMux I__3806 (
            .O(N__25196),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    InMux I__3805 (
            .O(N__25193),
            .I(N__25190));
    LocalMux I__3804 (
            .O(N__25190),
            .I(N__25187));
    Odrv12 I__3803 (
            .O(N__25187),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ));
    CascadeMux I__3802 (
            .O(N__25184),
            .I(N__25181));
    InMux I__3801 (
            .O(N__25181),
            .I(N__25178));
    LocalMux I__3800 (
            .O(N__25178),
            .I(N__25175));
    Odrv4 I__3799 (
            .O(N__25175),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    InMux I__3798 (
            .O(N__25172),
            .I(N__25169));
    LocalMux I__3797 (
            .O(N__25169),
            .I(N__25166));
    Span4Mux_v I__3796 (
            .O(N__25166),
            .I(N__25161));
    InMux I__3795 (
            .O(N__25165),
            .I(N__25158));
    InMux I__3794 (
            .O(N__25164),
            .I(N__25155));
    Span4Mux_v I__3793 (
            .O(N__25161),
            .I(N__25149));
    LocalMux I__3792 (
            .O(N__25158),
            .I(N__25149));
    LocalMux I__3791 (
            .O(N__25155),
            .I(N__25146));
    InMux I__3790 (
            .O(N__25154),
            .I(N__25143));
    Span4Mux_h I__3789 (
            .O(N__25149),
            .I(N__25140));
    Span12Mux_h I__3788 (
            .O(N__25146),
            .I(N__25137));
    LocalMux I__3787 (
            .O(N__25143),
            .I(N__25134));
    Odrv4 I__3786 (
            .O(N__25140),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    Odrv12 I__3785 (
            .O(N__25137),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    Odrv12 I__3784 (
            .O(N__25134),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    InMux I__3783 (
            .O(N__25127),
            .I(N__25124));
    LocalMux I__3782 (
            .O(N__25124),
            .I(N__25119));
    InMux I__3781 (
            .O(N__25123),
            .I(N__25116));
    InMux I__3780 (
            .O(N__25122),
            .I(N__25113));
    Span4Mux_v I__3779 (
            .O(N__25119),
            .I(N__25108));
    LocalMux I__3778 (
            .O(N__25116),
            .I(N__25108));
    LocalMux I__3777 (
            .O(N__25113),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    Odrv4 I__3776 (
            .O(N__25108),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    CascadeMux I__3775 (
            .O(N__25103),
            .I(N__25098));
    InMux I__3774 (
            .O(N__25102),
            .I(N__25095));
    InMux I__3773 (
            .O(N__25101),
            .I(N__25092));
    InMux I__3772 (
            .O(N__25098),
            .I(N__25089));
    LocalMux I__3771 (
            .O(N__25095),
            .I(N__25084));
    LocalMux I__3770 (
            .O(N__25092),
            .I(N__25084));
    LocalMux I__3769 (
            .O(N__25089),
            .I(N__25081));
    Span4Mux_h I__3768 (
            .O(N__25084),
            .I(N__25077));
    Span4Mux_v I__3767 (
            .O(N__25081),
            .I(N__25074));
    InMux I__3766 (
            .O(N__25080),
            .I(N__25071));
    Span4Mux_v I__3765 (
            .O(N__25077),
            .I(N__25068));
    Span4Mux_h I__3764 (
            .O(N__25074),
            .I(N__25063));
    LocalMux I__3763 (
            .O(N__25071),
            .I(N__25063));
    Odrv4 I__3762 (
            .O(N__25068),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    Odrv4 I__3761 (
            .O(N__25063),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    InMux I__3760 (
            .O(N__25058),
            .I(N__25054));
    InMux I__3759 (
            .O(N__25057),
            .I(N__25050));
    LocalMux I__3758 (
            .O(N__25054),
            .I(N__25047));
    InMux I__3757 (
            .O(N__25053),
            .I(N__25044));
    LocalMux I__3756 (
            .O(N__25050),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    Odrv12 I__3755 (
            .O(N__25047),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    LocalMux I__3754 (
            .O(N__25044),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    InMux I__3753 (
            .O(N__25037),
            .I(N__25028));
    InMux I__3752 (
            .O(N__25036),
            .I(N__25028));
    InMux I__3751 (
            .O(N__25035),
            .I(N__25028));
    LocalMux I__3750 (
            .O(N__25028),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ));
    CascadeMux I__3749 (
            .O(N__25025),
            .I(N__25022));
    InMux I__3748 (
            .O(N__25022),
            .I(N__25013));
    InMux I__3747 (
            .O(N__25021),
            .I(N__25013));
    InMux I__3746 (
            .O(N__25020),
            .I(N__25013));
    LocalMux I__3745 (
            .O(N__25013),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ));
    CascadeMux I__3744 (
            .O(N__25010),
            .I(\phase_controller_inst1.stoper_hc.un4_running_df30_cascade_ ));
    InMux I__3743 (
            .O(N__25007),
            .I(N__25004));
    LocalMux I__3742 (
            .O(N__25004),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ));
    CascadeMux I__3741 (
            .O(N__25001),
            .I(N__24998));
    InMux I__3740 (
            .O(N__24998),
            .I(N__24995));
    LocalMux I__3739 (
            .O(N__24995),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    InMux I__3738 (
            .O(N__24992),
            .I(N__24989));
    LocalMux I__3737 (
            .O(N__24989),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ));
    CascadeMux I__3736 (
            .O(N__24986),
            .I(N__24983));
    InMux I__3735 (
            .O(N__24983),
            .I(N__24980));
    LocalMux I__3734 (
            .O(N__24980),
            .I(N__24977));
    Odrv4 I__3733 (
            .O(N__24977),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    InMux I__3732 (
            .O(N__24974),
            .I(N__24971));
    LocalMux I__3731 (
            .O(N__24971),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ));
    CascadeMux I__3730 (
            .O(N__24968),
            .I(N__24965));
    InMux I__3729 (
            .O(N__24965),
            .I(N__24962));
    LocalMux I__3728 (
            .O(N__24962),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    InMux I__3727 (
            .O(N__24959),
            .I(N__24956));
    LocalMux I__3726 (
            .O(N__24956),
            .I(\current_shift_inst.un4_control_input_1_axb_26 ));
    InMux I__3725 (
            .O(N__24953),
            .I(N__24947));
    InMux I__3724 (
            .O(N__24952),
            .I(N__24947));
    LocalMux I__3723 (
            .O(N__24947),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ));
    InMux I__3722 (
            .O(N__24944),
            .I(N__24941));
    LocalMux I__3721 (
            .O(N__24941),
            .I(N__24938));
    Span12Mux_s11_h I__3720 (
            .O(N__24938),
            .I(N__24934));
    InMux I__3719 (
            .O(N__24937),
            .I(N__24931));
    Odrv12 I__3718 (
            .O(N__24934),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    LocalMux I__3717 (
            .O(N__24931),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    CascadeMux I__3716 (
            .O(N__24926),
            .I(elapsed_time_ns_1_RNII43T9_0_6_cascade_));
    InMux I__3715 (
            .O(N__24923),
            .I(N__24917));
    InMux I__3714 (
            .O(N__24922),
            .I(N__24917));
    LocalMux I__3713 (
            .O(N__24917),
            .I(N__24913));
    InMux I__3712 (
            .O(N__24916),
            .I(N__24910));
    Span4Mux_v I__3711 (
            .O(N__24913),
            .I(N__24906));
    LocalMux I__3710 (
            .O(N__24910),
            .I(N__24903));
    InMux I__3709 (
            .O(N__24909),
            .I(N__24900));
    Span4Mux_v I__3708 (
            .O(N__24906),
            .I(N__24895));
    Span4Mux_v I__3707 (
            .O(N__24903),
            .I(N__24895));
    LocalMux I__3706 (
            .O(N__24900),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    Odrv4 I__3705 (
            .O(N__24895),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    InMux I__3704 (
            .O(N__24890),
            .I(N__24887));
    LocalMux I__3703 (
            .O(N__24887),
            .I(\current_shift_inst.un4_control_input_1_axb_25 ));
    InMux I__3702 (
            .O(N__24884),
            .I(bfn_10_21_0_));
    InMux I__3701 (
            .O(N__24881),
            .I(\current_shift_inst.un4_control_input_1_cry_25 ));
    InMux I__3700 (
            .O(N__24878),
            .I(\current_shift_inst.un4_control_input_1_cry_26 ));
    InMux I__3699 (
            .O(N__24875),
            .I(N__24872));
    LocalMux I__3698 (
            .O(N__24872),
            .I(\current_shift_inst.un4_control_input_1_axb_28 ));
    InMux I__3697 (
            .O(N__24869),
            .I(\current_shift_inst.un4_control_input_1_cry_27 ));
    InMux I__3696 (
            .O(N__24866),
            .I(N__24863));
    LocalMux I__3695 (
            .O(N__24863),
            .I(N__24860));
    Span4Mux_h I__3694 (
            .O(N__24860),
            .I(N__24857));
    Odrv4 I__3693 (
            .O(N__24857),
            .I(\current_shift_inst.un4_control_input_1_axb_29 ));
    InMux I__3692 (
            .O(N__24854),
            .I(\current_shift_inst.un4_control_input_1_cry_28 ));
    InMux I__3691 (
            .O(N__24851),
            .I(\current_shift_inst.un4_control_input1_31 ));
    CascadeMux I__3690 (
            .O(N__24848),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO_cascade_ ));
    InMux I__3689 (
            .O(N__24845),
            .I(N__24842));
    LocalMux I__3688 (
            .O(N__24842),
            .I(\current_shift_inst.un4_control_input_1_axb_18 ));
    InMux I__3687 (
            .O(N__24839),
            .I(N__24836));
    LocalMux I__3686 (
            .O(N__24836),
            .I(\current_shift_inst.un4_control_input_1_axb_27 ));
    InMux I__3685 (
            .O(N__24833),
            .I(N__24830));
    LocalMux I__3684 (
            .O(N__24830),
            .I(\current_shift_inst.un4_control_input_1_axb_17 ));
    InMux I__3683 (
            .O(N__24827),
            .I(bfn_10_20_0_));
    InMux I__3682 (
            .O(N__24824),
            .I(\current_shift_inst.un4_control_input_1_cry_17 ));
    CascadeMux I__3681 (
            .O(N__24821),
            .I(N__24818));
    InMux I__3680 (
            .O(N__24818),
            .I(N__24815));
    LocalMux I__3679 (
            .O(N__24815),
            .I(N__24812));
    Odrv4 I__3678 (
            .O(N__24812),
            .I(\current_shift_inst.un4_control_input_1_axb_19 ));
    InMux I__3677 (
            .O(N__24809),
            .I(\current_shift_inst.un4_control_input_1_cry_18 ));
    InMux I__3676 (
            .O(N__24806),
            .I(N__24803));
    LocalMux I__3675 (
            .O(N__24803),
            .I(\current_shift_inst.un4_control_input_1_axb_20 ));
    InMux I__3674 (
            .O(N__24800),
            .I(\current_shift_inst.un4_control_input_1_cry_19 ));
    InMux I__3673 (
            .O(N__24797),
            .I(N__24794));
    LocalMux I__3672 (
            .O(N__24794),
            .I(N__24791));
    Odrv4 I__3671 (
            .O(N__24791),
            .I(\current_shift_inst.un4_control_input_1_axb_21 ));
    InMux I__3670 (
            .O(N__24788),
            .I(N__24783));
    InMux I__3669 (
            .O(N__24787),
            .I(N__24780));
    InMux I__3668 (
            .O(N__24786),
            .I(N__24777));
    LocalMux I__3667 (
            .O(N__24783),
            .I(N__24774));
    LocalMux I__3666 (
            .O(N__24780),
            .I(N__24769));
    LocalMux I__3665 (
            .O(N__24777),
            .I(N__24769));
    Sp12to4 I__3664 (
            .O(N__24774),
            .I(N__24766));
    Span4Mux_v I__3663 (
            .O(N__24769),
            .I(N__24763));
    Odrv12 I__3662 (
            .O(N__24766),
            .I(\current_shift_inst.un4_control_input1_22 ));
    Odrv4 I__3661 (
            .O(N__24763),
            .I(\current_shift_inst.un4_control_input1_22 ));
    InMux I__3660 (
            .O(N__24758),
            .I(\current_shift_inst.un4_control_input_1_cry_20 ));
    InMux I__3659 (
            .O(N__24755),
            .I(N__24752));
    LocalMux I__3658 (
            .O(N__24752),
            .I(N__24749));
    Span4Mux_h I__3657 (
            .O(N__24749),
            .I(N__24746));
    Odrv4 I__3656 (
            .O(N__24746),
            .I(\current_shift_inst.un4_control_input_1_axb_22 ));
    InMux I__3655 (
            .O(N__24743),
            .I(\current_shift_inst.un4_control_input_1_cry_21 ));
    InMux I__3654 (
            .O(N__24740),
            .I(N__24737));
    LocalMux I__3653 (
            .O(N__24737),
            .I(N__24734));
    Odrv4 I__3652 (
            .O(N__24734),
            .I(\current_shift_inst.un4_control_input_1_axb_23 ));
    InMux I__3651 (
            .O(N__24731),
            .I(\current_shift_inst.un4_control_input_1_cry_22 ));
    InMux I__3650 (
            .O(N__24728),
            .I(N__24725));
    LocalMux I__3649 (
            .O(N__24725),
            .I(\current_shift_inst.un4_control_input_1_axb_24 ));
    InMux I__3648 (
            .O(N__24722),
            .I(\current_shift_inst.un4_control_input_1_cry_23 ));
    InMux I__3647 (
            .O(N__24719),
            .I(N__24716));
    LocalMux I__3646 (
            .O(N__24716),
            .I(N__24713));
    Odrv4 I__3645 (
            .O(N__24713),
            .I(\current_shift_inst.un4_control_input_1_axb_8 ));
    InMux I__3644 (
            .O(N__24710),
            .I(\current_shift_inst.un4_control_input_1_cry_7 ));
    InMux I__3643 (
            .O(N__24707),
            .I(N__24704));
    LocalMux I__3642 (
            .O(N__24704),
            .I(N__24701));
    Odrv4 I__3641 (
            .O(N__24701),
            .I(\current_shift_inst.un4_control_input_1_axb_9 ));
    InMux I__3640 (
            .O(N__24698),
            .I(N__24693));
    InMux I__3639 (
            .O(N__24697),
            .I(N__24690));
    InMux I__3638 (
            .O(N__24696),
            .I(N__24687));
    LocalMux I__3637 (
            .O(N__24693),
            .I(N__24684));
    LocalMux I__3636 (
            .O(N__24690),
            .I(N__24679));
    LocalMux I__3635 (
            .O(N__24687),
            .I(N__24679));
    Odrv12 I__3634 (
            .O(N__24684),
            .I(\current_shift_inst.un4_control_input1_10 ));
    Odrv12 I__3633 (
            .O(N__24679),
            .I(\current_shift_inst.un4_control_input1_10 ));
    InMux I__3632 (
            .O(N__24674),
            .I(bfn_10_19_0_));
    InMux I__3631 (
            .O(N__24671),
            .I(N__24668));
    LocalMux I__3630 (
            .O(N__24668),
            .I(N__24665));
    Odrv4 I__3629 (
            .O(N__24665),
            .I(\current_shift_inst.un4_control_input_1_axb_10 ));
    InMux I__3628 (
            .O(N__24662),
            .I(\current_shift_inst.un4_control_input_1_cry_9 ));
    InMux I__3627 (
            .O(N__24659),
            .I(\current_shift_inst.un4_control_input_1_cry_10 ));
    InMux I__3626 (
            .O(N__24656),
            .I(N__24653));
    LocalMux I__3625 (
            .O(N__24653),
            .I(N__24650));
    Odrv12 I__3624 (
            .O(N__24650),
            .I(\current_shift_inst.un4_control_input_1_axb_12 ));
    InMux I__3623 (
            .O(N__24647),
            .I(\current_shift_inst.un4_control_input_1_cry_11 ));
    InMux I__3622 (
            .O(N__24644),
            .I(N__24641));
    LocalMux I__3621 (
            .O(N__24641),
            .I(N__24638));
    Odrv4 I__3620 (
            .O(N__24638),
            .I(\current_shift_inst.un4_control_input_1_axb_13 ));
    InMux I__3619 (
            .O(N__24635),
            .I(\current_shift_inst.un4_control_input_1_cry_12 ));
    InMux I__3618 (
            .O(N__24632),
            .I(\current_shift_inst.un4_control_input_1_cry_13 ));
    InMux I__3617 (
            .O(N__24629),
            .I(N__24626));
    LocalMux I__3616 (
            .O(N__24626),
            .I(N__24623));
    Odrv12 I__3615 (
            .O(N__24623),
            .I(\current_shift_inst.un4_control_input_1_axb_15 ));
    InMux I__3614 (
            .O(N__24620),
            .I(N__24615));
    InMux I__3613 (
            .O(N__24619),
            .I(N__24610));
    InMux I__3612 (
            .O(N__24618),
            .I(N__24610));
    LocalMux I__3611 (
            .O(N__24615),
            .I(N__24605));
    LocalMux I__3610 (
            .O(N__24610),
            .I(N__24605));
    Odrv12 I__3609 (
            .O(N__24605),
            .I(\current_shift_inst.un4_control_input1_16 ));
    InMux I__3608 (
            .O(N__24602),
            .I(\current_shift_inst.un4_control_input_1_cry_14 ));
    InMux I__3607 (
            .O(N__24599),
            .I(N__24596));
    LocalMux I__3606 (
            .O(N__24596),
            .I(N__24593));
    Odrv12 I__3605 (
            .O(N__24593),
            .I(\current_shift_inst.un4_control_input_1_axb_16 ));
    InMux I__3604 (
            .O(N__24590),
            .I(\current_shift_inst.un4_control_input_1_cry_15 ));
    CascadeMux I__3603 (
            .O(N__24587),
            .I(N__24584));
    InMux I__3602 (
            .O(N__24584),
            .I(N__24581));
    LocalMux I__3601 (
            .O(N__24581),
            .I(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ));
    InMux I__3600 (
            .O(N__24578),
            .I(N__24575));
    LocalMux I__3599 (
            .O(N__24575),
            .I(N__24572));
    Odrv12 I__3598 (
            .O(N__24572),
            .I(\current_shift_inst.un4_control_input_1_axb_1 ));
    InMux I__3597 (
            .O(N__24569),
            .I(N__24560));
    InMux I__3596 (
            .O(N__24568),
            .I(N__24560));
    InMux I__3595 (
            .O(N__24567),
            .I(N__24560));
    LocalMux I__3594 (
            .O(N__24560),
            .I(N__24557));
    Odrv12 I__3593 (
            .O(N__24557),
            .I(\current_shift_inst.un4_control_input1_2 ));
    InMux I__3592 (
            .O(N__24554),
            .I(N__24551));
    LocalMux I__3591 (
            .O(N__24551),
            .I(N__24548));
    Span4Mux_h I__3590 (
            .O(N__24548),
            .I(N__24545));
    Odrv4 I__3589 (
            .O(N__24545),
            .I(\current_shift_inst.un4_control_input_1_axb_2 ));
    InMux I__3588 (
            .O(N__24542),
            .I(\current_shift_inst.un4_control_input_1_cry_1 ));
    InMux I__3587 (
            .O(N__24539),
            .I(N__24536));
    LocalMux I__3586 (
            .O(N__24536),
            .I(N__24533));
    Span4Mux_h I__3585 (
            .O(N__24533),
            .I(N__24530));
    Odrv4 I__3584 (
            .O(N__24530),
            .I(\current_shift_inst.un4_control_input_1_axb_3 ));
    InMux I__3583 (
            .O(N__24527),
            .I(\current_shift_inst.un4_control_input_1_cry_2 ));
    InMux I__3582 (
            .O(N__24524),
            .I(N__24521));
    LocalMux I__3581 (
            .O(N__24521),
            .I(N__24518));
    Span4Mux_v I__3580 (
            .O(N__24518),
            .I(N__24515));
    Odrv4 I__3579 (
            .O(N__24515),
            .I(\current_shift_inst.un4_control_input_1_axb_4 ));
    InMux I__3578 (
            .O(N__24512),
            .I(\current_shift_inst.un4_control_input_1_cry_3 ));
    InMux I__3577 (
            .O(N__24509),
            .I(N__24506));
    LocalMux I__3576 (
            .O(N__24506),
            .I(N__24503));
    Odrv12 I__3575 (
            .O(N__24503),
            .I(\current_shift_inst.un4_control_input_1_axb_5 ));
    CascadeMux I__3574 (
            .O(N__24500),
            .I(N__24496));
    CascadeMux I__3573 (
            .O(N__24499),
            .I(N__24493));
    InMux I__3572 (
            .O(N__24496),
            .I(N__24490));
    InMux I__3571 (
            .O(N__24493),
            .I(N__24487));
    LocalMux I__3570 (
            .O(N__24490),
            .I(N__24484));
    LocalMux I__3569 (
            .O(N__24487),
            .I(N__24478));
    Span4Mux_v I__3568 (
            .O(N__24484),
            .I(N__24478));
    InMux I__3567 (
            .O(N__24483),
            .I(N__24475));
    Odrv4 I__3566 (
            .O(N__24478),
            .I(\current_shift_inst.un4_control_input1_6 ));
    LocalMux I__3565 (
            .O(N__24475),
            .I(\current_shift_inst.un4_control_input1_6 ));
    InMux I__3564 (
            .O(N__24470),
            .I(\current_shift_inst.un4_control_input_1_cry_4 ));
    InMux I__3563 (
            .O(N__24467),
            .I(N__24464));
    LocalMux I__3562 (
            .O(N__24464),
            .I(N__24461));
    Span4Mux_h I__3561 (
            .O(N__24461),
            .I(N__24458));
    Odrv4 I__3560 (
            .O(N__24458),
            .I(\current_shift_inst.un4_control_input_1_axb_6 ));
    InMux I__3559 (
            .O(N__24455),
            .I(\current_shift_inst.un4_control_input_1_cry_5 ));
    InMux I__3558 (
            .O(N__24452),
            .I(N__24449));
    LocalMux I__3557 (
            .O(N__24449),
            .I(N__24446));
    Odrv12 I__3556 (
            .O(N__24446),
            .I(\current_shift_inst.un4_control_input_1_axb_7 ));
    InMux I__3555 (
            .O(N__24443),
            .I(\current_shift_inst.un4_control_input_1_cry_6 ));
    InMux I__3554 (
            .O(N__24440),
            .I(N__24437));
    LocalMux I__3553 (
            .O(N__24437),
            .I(N__24432));
    InMux I__3552 (
            .O(N__24436),
            .I(N__24427));
    InMux I__3551 (
            .O(N__24435),
            .I(N__24427));
    Span4Mux_v I__3550 (
            .O(N__24432),
            .I(N__24422));
    LocalMux I__3549 (
            .O(N__24427),
            .I(N__24422));
    Span4Mux_h I__3548 (
            .O(N__24422),
            .I(N__24418));
    InMux I__3547 (
            .O(N__24421),
            .I(N__24415));
    Span4Mux_v I__3546 (
            .O(N__24418),
            .I(N__24412));
    LocalMux I__3545 (
            .O(N__24415),
            .I(N__24409));
    Odrv4 I__3544 (
            .O(N__24412),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    Odrv4 I__3543 (
            .O(N__24409),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    CascadeMux I__3542 (
            .O(N__24404),
            .I(N__24401));
    InMux I__3541 (
            .O(N__24401),
            .I(N__24398));
    LocalMux I__3540 (
            .O(N__24398),
            .I(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ));
    InMux I__3539 (
            .O(N__24395),
            .I(N__24391));
    InMux I__3538 (
            .O(N__24394),
            .I(N__24388));
    LocalMux I__3537 (
            .O(N__24391),
            .I(N__24382));
    LocalMux I__3536 (
            .O(N__24388),
            .I(N__24382));
    InMux I__3535 (
            .O(N__24387),
            .I(N__24379));
    Span4Mux_v I__3534 (
            .O(N__24382),
            .I(N__24375));
    LocalMux I__3533 (
            .O(N__24379),
            .I(N__24372));
    InMux I__3532 (
            .O(N__24378),
            .I(N__24369));
    Span4Mux_h I__3531 (
            .O(N__24375),
            .I(N__24366));
    Span4Mux_h I__3530 (
            .O(N__24372),
            .I(N__24361));
    LocalMux I__3529 (
            .O(N__24369),
            .I(N__24361));
    Odrv4 I__3528 (
            .O(N__24366),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    Odrv4 I__3527 (
            .O(N__24361),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    CascadeMux I__3526 (
            .O(N__24356),
            .I(N__24353));
    InMux I__3525 (
            .O(N__24353),
            .I(N__24350));
    LocalMux I__3524 (
            .O(N__24350),
            .I(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ));
    CascadeMux I__3523 (
            .O(N__24347),
            .I(N__24344));
    InMux I__3522 (
            .O(N__24344),
            .I(N__24341));
    LocalMux I__3521 (
            .O(N__24341),
            .I(N__24338));
    Odrv4 I__3520 (
            .O(N__24338),
            .I(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ));
    CascadeMux I__3519 (
            .O(N__24335),
            .I(N__24332));
    InMux I__3518 (
            .O(N__24332),
            .I(N__24329));
    LocalMux I__3517 (
            .O(N__24329),
            .I(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ));
    InMux I__3516 (
            .O(N__24326),
            .I(N__24323));
    LocalMux I__3515 (
            .O(N__24323),
            .I(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ));
    InMux I__3514 (
            .O(N__24320),
            .I(N__24317));
    LocalMux I__3513 (
            .O(N__24317),
            .I(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ));
    InMux I__3512 (
            .O(N__24314),
            .I(N__24311));
    LocalMux I__3511 (
            .O(N__24311),
            .I(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ));
    CascadeMux I__3510 (
            .O(N__24308),
            .I(N__24305));
    InMux I__3509 (
            .O(N__24305),
            .I(N__24302));
    LocalMux I__3508 (
            .O(N__24302),
            .I(N__24299));
    Span4Mux_v I__3507 (
            .O(N__24299),
            .I(N__24296));
    Odrv4 I__3506 (
            .O(N__24296),
            .I(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ));
    InMux I__3505 (
            .O(N__24293),
            .I(N__24290));
    LocalMux I__3504 (
            .O(N__24290),
            .I(\current_shift_inst.control_input_axb_0 ));
    CascadeMux I__3503 (
            .O(N__24287),
            .I(\current_shift_inst.control_input_axb_0_cascade_ ));
    CascadeMux I__3502 (
            .O(N__24284),
            .I(N__24279));
    InMux I__3501 (
            .O(N__24283),
            .I(N__24276));
    InMux I__3500 (
            .O(N__24282),
            .I(N__24273));
    InMux I__3499 (
            .O(N__24279),
            .I(N__24270));
    LocalMux I__3498 (
            .O(N__24276),
            .I(\current_shift_inst.N_1288_i ));
    LocalMux I__3497 (
            .O(N__24273),
            .I(\current_shift_inst.N_1288_i ));
    LocalMux I__3496 (
            .O(N__24270),
            .I(\current_shift_inst.N_1288_i ));
    CascadeMux I__3495 (
            .O(N__24263),
            .I(N__24259));
    InMux I__3494 (
            .O(N__24262),
            .I(N__24256));
    InMux I__3493 (
            .O(N__24259),
            .I(N__24253));
    LocalMux I__3492 (
            .O(N__24256),
            .I(N__24250));
    LocalMux I__3491 (
            .O(N__24253),
            .I(N__24246));
    Span4Mux_v I__3490 (
            .O(N__24250),
            .I(N__24243));
    InMux I__3489 (
            .O(N__24249),
            .I(N__24240));
    Span4Mux_h I__3488 (
            .O(N__24246),
            .I(N__24237));
    Sp12to4 I__3487 (
            .O(N__24243),
            .I(N__24232));
    LocalMux I__3486 (
            .O(N__24240),
            .I(N__24232));
    Span4Mux_v I__3485 (
            .O(N__24237),
            .I(N__24228));
    Span12Mux_h I__3484 (
            .O(N__24232),
            .I(N__24225));
    InMux I__3483 (
            .O(N__24231),
            .I(N__24222));
    Odrv4 I__3482 (
            .O(N__24228),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    Odrv12 I__3481 (
            .O(N__24225),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    LocalMux I__3480 (
            .O(N__24222),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    CascadeMux I__3479 (
            .O(N__24215),
            .I(N__24212));
    InMux I__3478 (
            .O(N__24212),
            .I(N__24209));
    LocalMux I__3477 (
            .O(N__24209),
            .I(N__24206));
    Span4Mux_v I__3476 (
            .O(N__24206),
            .I(N__24203));
    Span4Mux_h I__3475 (
            .O(N__24203),
            .I(N__24200));
    Odrv4 I__3474 (
            .O(N__24200),
            .I(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ));
    InMux I__3473 (
            .O(N__24197),
            .I(N__24194));
    LocalMux I__3472 (
            .O(N__24194),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt26 ));
    CascadeMux I__3471 (
            .O(N__24191),
            .I(N__24188));
    InMux I__3470 (
            .O(N__24188),
            .I(N__24178));
    InMux I__3469 (
            .O(N__24187),
            .I(N__24178));
    InMux I__3468 (
            .O(N__24186),
            .I(N__24178));
    InMux I__3467 (
            .O(N__24185),
            .I(N__24175));
    LocalMux I__3466 (
            .O(N__24178),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    LocalMux I__3465 (
            .O(N__24175),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    InMux I__3464 (
            .O(N__24170),
            .I(N__24167));
    LocalMux I__3463 (
            .O(N__24167),
            .I(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ));
    CascadeMux I__3462 (
            .O(N__24164),
            .I(N__24161));
    InMux I__3461 (
            .O(N__24161),
            .I(N__24158));
    LocalMux I__3460 (
            .O(N__24158),
            .I(N__24155));
    Odrv4 I__3459 (
            .O(N__24155),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt16 ));
    InMux I__3458 (
            .O(N__24152),
            .I(N__24149));
    LocalMux I__3457 (
            .O(N__24149),
            .I(N__24144));
    InMux I__3456 (
            .O(N__24148),
            .I(N__24139));
    InMux I__3455 (
            .O(N__24147),
            .I(N__24139));
    Span4Mux_v I__3454 (
            .O(N__24144),
            .I(N__24136));
    LocalMux I__3453 (
            .O(N__24139),
            .I(N__24132));
    Span4Mux_v I__3452 (
            .O(N__24136),
            .I(N__24129));
    InMux I__3451 (
            .O(N__24135),
            .I(N__24126));
    Span4Mux_v I__3450 (
            .O(N__24132),
            .I(N__24123));
    Span4Mux_v I__3449 (
            .O(N__24129),
            .I(N__24118));
    LocalMux I__3448 (
            .O(N__24126),
            .I(N__24118));
    Odrv4 I__3447 (
            .O(N__24123),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    Odrv4 I__3446 (
            .O(N__24118),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    InMux I__3445 (
            .O(N__24113),
            .I(N__24110));
    LocalMux I__3444 (
            .O(N__24110),
            .I(N__24107));
    Span4Mux_v I__3443 (
            .O(N__24107),
            .I(N__24104));
    Span4Mux_v I__3442 (
            .O(N__24104),
            .I(N__24101));
    Odrv4 I__3441 (
            .O(N__24101),
            .I(il_min_comp1_D1));
    InMux I__3440 (
            .O(N__24098),
            .I(N__24092));
    InMux I__3439 (
            .O(N__24097),
            .I(N__24092));
    LocalMux I__3438 (
            .O(N__24092),
            .I(N__24089));
    Odrv4 I__3437 (
            .O(N__24089),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ));
    CascadeMux I__3436 (
            .O(N__24086),
            .I(N__24082));
    CascadeMux I__3435 (
            .O(N__24085),
            .I(N__24079));
    InMux I__3434 (
            .O(N__24082),
            .I(N__24074));
    InMux I__3433 (
            .O(N__24079),
            .I(N__24074));
    LocalMux I__3432 (
            .O(N__24074),
            .I(N__24071));
    Odrv4 I__3431 (
            .O(N__24071),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ));
    InMux I__3430 (
            .O(N__24068),
            .I(N__24065));
    LocalMux I__3429 (
            .O(N__24065),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ));
    InMux I__3428 (
            .O(N__24062),
            .I(N__24059));
    LocalMux I__3427 (
            .O(N__24059),
            .I(N__24054));
    InMux I__3426 (
            .O(N__24058),
            .I(N__24051));
    InMux I__3425 (
            .O(N__24057),
            .I(N__24048));
    Span4Mux_v I__3424 (
            .O(N__24054),
            .I(N__24043));
    LocalMux I__3423 (
            .O(N__24051),
            .I(N__24043));
    LocalMux I__3422 (
            .O(N__24048),
            .I(N__24037));
    Span4Mux_h I__3421 (
            .O(N__24043),
            .I(N__24037));
    InMux I__3420 (
            .O(N__24042),
            .I(N__24034));
    Span4Mux_v I__3419 (
            .O(N__24037),
            .I(N__24029));
    LocalMux I__3418 (
            .O(N__24034),
            .I(N__24029));
    Span4Mux_v I__3417 (
            .O(N__24029),
            .I(N__24026));
    Odrv4 I__3416 (
            .O(N__24026),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    InMux I__3415 (
            .O(N__24023),
            .I(N__24018));
    InMux I__3414 (
            .O(N__24022),
            .I(N__24015));
    InMux I__3413 (
            .O(N__24021),
            .I(N__24012));
    LocalMux I__3412 (
            .O(N__24018),
            .I(N__24009));
    LocalMux I__3411 (
            .O(N__24015),
            .I(N__24006));
    LocalMux I__3410 (
            .O(N__24012),
            .I(N__24000));
    Span4Mux_h I__3409 (
            .O(N__24009),
            .I(N__24000));
    Span4Mux_v I__3408 (
            .O(N__24006),
            .I(N__23997));
    InMux I__3407 (
            .O(N__24005),
            .I(N__23994));
    Span4Mux_v I__3406 (
            .O(N__24000),
            .I(N__23991));
    Span4Mux_v I__3405 (
            .O(N__23997),
            .I(N__23986));
    LocalMux I__3404 (
            .O(N__23994),
            .I(N__23986));
    Odrv4 I__3403 (
            .O(N__23991),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    Odrv4 I__3402 (
            .O(N__23986),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    InMux I__3401 (
            .O(N__23981),
            .I(N__23978));
    LocalMux I__3400 (
            .O(N__23978),
            .I(N__23975));
    Span4Mux_h I__3399 (
            .O(N__23975),
            .I(N__23972));
    Span4Mux_v I__3398 (
            .O(N__23972),
            .I(N__23969));
    Odrv4 I__3397 (
            .O(N__23969),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ));
    InMux I__3396 (
            .O(N__23966),
            .I(N__23963));
    LocalMux I__3395 (
            .O(N__23963),
            .I(N__23960));
    Span4Mux_v I__3394 (
            .O(N__23960),
            .I(N__23957));
    Span4Mux_v I__3393 (
            .O(N__23957),
            .I(N__23952));
    InMux I__3392 (
            .O(N__23956),
            .I(N__23949));
    InMux I__3391 (
            .O(N__23955),
            .I(N__23946));
    Odrv4 I__3390 (
            .O(N__23952),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    LocalMux I__3389 (
            .O(N__23949),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    LocalMux I__3388 (
            .O(N__23946),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    InMux I__3387 (
            .O(N__23939),
            .I(N__23934));
    InMux I__3386 (
            .O(N__23938),
            .I(N__23930));
    InMux I__3385 (
            .O(N__23937),
            .I(N__23927));
    LocalMux I__3384 (
            .O(N__23934),
            .I(N__23924));
    InMux I__3383 (
            .O(N__23933),
            .I(N__23921));
    LocalMux I__3382 (
            .O(N__23930),
            .I(N__23918));
    LocalMux I__3381 (
            .O(N__23927),
            .I(N__23915));
    Span4Mux_h I__3380 (
            .O(N__23924),
            .I(N__23912));
    LocalMux I__3379 (
            .O(N__23921),
            .I(N__23909));
    Span4Mux_v I__3378 (
            .O(N__23918),
            .I(N__23904));
    Span4Mux_h I__3377 (
            .O(N__23915),
            .I(N__23904));
    Span4Mux_v I__3376 (
            .O(N__23912),
            .I(N__23899));
    Span4Mux_h I__3375 (
            .O(N__23909),
            .I(N__23899));
    Span4Mux_v I__3374 (
            .O(N__23904),
            .I(N__23896));
    Odrv4 I__3373 (
            .O(N__23899),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    Odrv4 I__3372 (
            .O(N__23896),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    InMux I__3371 (
            .O(N__23891),
            .I(N__23888));
    LocalMux I__3370 (
            .O(N__23888),
            .I(N__23885));
    Span4Mux_v I__3369 (
            .O(N__23885),
            .I(N__23880));
    InMux I__3368 (
            .O(N__23884),
            .I(N__23877));
    InMux I__3367 (
            .O(N__23883),
            .I(N__23874));
    Sp12to4 I__3366 (
            .O(N__23880),
            .I(N__23869));
    LocalMux I__3365 (
            .O(N__23877),
            .I(N__23869));
    LocalMux I__3364 (
            .O(N__23874),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    Odrv12 I__3363 (
            .O(N__23869),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    InMux I__3362 (
            .O(N__23864),
            .I(N__23860));
    InMux I__3361 (
            .O(N__23863),
            .I(N__23857));
    LocalMux I__3360 (
            .O(N__23860),
            .I(N__23853));
    LocalMux I__3359 (
            .O(N__23857),
            .I(N__23849));
    InMux I__3358 (
            .O(N__23856),
            .I(N__23846));
    Span4Mux_v I__3357 (
            .O(N__23853),
            .I(N__23843));
    InMux I__3356 (
            .O(N__23852),
            .I(N__23840));
    Odrv4 I__3355 (
            .O(N__23849),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    LocalMux I__3354 (
            .O(N__23846),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    Odrv4 I__3353 (
            .O(N__23843),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    LocalMux I__3352 (
            .O(N__23840),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    InMux I__3351 (
            .O(N__23831),
            .I(N__23828));
    LocalMux I__3350 (
            .O(N__23828),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ));
    CascadeMux I__3349 (
            .O(N__23825),
            .I(\phase_controller_inst2.stoper_hc.un4_running_df30_cascade_ ));
    InMux I__3348 (
            .O(N__23822),
            .I(N__23819));
    LocalMux I__3347 (
            .O(N__23819),
            .I(N__23816));
    Odrv4 I__3346 (
            .O(N__23816),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO ));
    CascadeMux I__3345 (
            .O(N__23813),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ));
    CascadeMux I__3344 (
            .O(N__23810),
            .I(N__23807));
    InMux I__3343 (
            .O(N__23807),
            .I(N__23804));
    LocalMux I__3342 (
            .O(N__23804),
            .I(N__23801));
    Span4Mux_v I__3341 (
            .O(N__23801),
            .I(N__23797));
    InMux I__3340 (
            .O(N__23800),
            .I(N__23794));
    Odrv4 I__3339 (
            .O(N__23797),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt30 ));
    LocalMux I__3338 (
            .O(N__23794),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt30 ));
    InMux I__3337 (
            .O(N__23789),
            .I(N__23780));
    InMux I__3336 (
            .O(N__23788),
            .I(N__23780));
    InMux I__3335 (
            .O(N__23787),
            .I(N__23780));
    LocalMux I__3334 (
            .O(N__23780),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ));
    InMux I__3333 (
            .O(N__23777),
            .I(N__23768));
    InMux I__3332 (
            .O(N__23776),
            .I(N__23768));
    InMux I__3331 (
            .O(N__23775),
            .I(N__23768));
    LocalMux I__3330 (
            .O(N__23768),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ));
    InMux I__3329 (
            .O(N__23765),
            .I(N__23762));
    LocalMux I__3328 (
            .O(N__23762),
            .I(N__23759));
    Odrv4 I__3327 (
            .O(N__23759),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ));
    CascadeMux I__3326 (
            .O(N__23756),
            .I(N__23753));
    InMux I__3325 (
            .O(N__23753),
            .I(N__23749));
    InMux I__3324 (
            .O(N__23752),
            .I(N__23746));
    LocalMux I__3323 (
            .O(N__23749),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ));
    LocalMux I__3322 (
            .O(N__23746),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ));
    InMux I__3321 (
            .O(N__23741),
            .I(N__23738));
    LocalMux I__3320 (
            .O(N__23738),
            .I(N__23733));
    InMux I__3319 (
            .O(N__23737),
            .I(N__23730));
    InMux I__3318 (
            .O(N__23736),
            .I(N__23727));
    Span4Mux_v I__3317 (
            .O(N__23733),
            .I(N__23724));
    LocalMux I__3316 (
            .O(N__23730),
            .I(N__23721));
    LocalMux I__3315 (
            .O(N__23727),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    Odrv4 I__3314 (
            .O(N__23724),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    Odrv12 I__3313 (
            .O(N__23721),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    InMux I__3312 (
            .O(N__23714),
            .I(N__23710));
    InMux I__3311 (
            .O(N__23713),
            .I(N__23707));
    LocalMux I__3310 (
            .O(N__23710),
            .I(N__23704));
    LocalMux I__3309 (
            .O(N__23707),
            .I(N__23700));
    Span4Mux_h I__3308 (
            .O(N__23704),
            .I(N__23696));
    InMux I__3307 (
            .O(N__23703),
            .I(N__23693));
    Span4Mux_h I__3306 (
            .O(N__23700),
            .I(N__23690));
    InMux I__3305 (
            .O(N__23699),
            .I(N__23687));
    Odrv4 I__3304 (
            .O(N__23696),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    LocalMux I__3303 (
            .O(N__23693),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    Odrv4 I__3302 (
            .O(N__23690),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    LocalMux I__3301 (
            .O(N__23687),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    InMux I__3300 (
            .O(N__23678),
            .I(N__23674));
    InMux I__3299 (
            .O(N__23677),
            .I(N__23671));
    LocalMux I__3298 (
            .O(N__23674),
            .I(N__23667));
    LocalMux I__3297 (
            .O(N__23671),
            .I(N__23664));
    InMux I__3296 (
            .O(N__23670),
            .I(N__23661));
    Span4Mux_v I__3295 (
            .O(N__23667),
            .I(N__23656));
    Span4Mux_h I__3294 (
            .O(N__23664),
            .I(N__23656));
    LocalMux I__3293 (
            .O(N__23661),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    Odrv4 I__3292 (
            .O(N__23656),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    InMux I__3291 (
            .O(N__23651),
            .I(N__23647));
    InMux I__3290 (
            .O(N__23650),
            .I(N__23644));
    LocalMux I__3289 (
            .O(N__23647),
            .I(N__23640));
    LocalMux I__3288 (
            .O(N__23644),
            .I(N__23637));
    InMux I__3287 (
            .O(N__23643),
            .I(N__23633));
    Span4Mux_h I__3286 (
            .O(N__23640),
            .I(N__23628));
    Span4Mux_h I__3285 (
            .O(N__23637),
            .I(N__23628));
    InMux I__3284 (
            .O(N__23636),
            .I(N__23625));
    LocalMux I__3283 (
            .O(N__23633),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    Odrv4 I__3282 (
            .O(N__23628),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    LocalMux I__3281 (
            .O(N__23625),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    InMux I__3280 (
            .O(N__23618),
            .I(N__23615));
    LocalMux I__3279 (
            .O(N__23615),
            .I(N__23612));
    Span4Mux_h I__3278 (
            .O(N__23612),
            .I(N__23607));
    InMux I__3277 (
            .O(N__23611),
            .I(N__23604));
    InMux I__3276 (
            .O(N__23610),
            .I(N__23601));
    Span4Mux_h I__3275 (
            .O(N__23607),
            .I(N__23598));
    LocalMux I__3274 (
            .O(N__23604),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    LocalMux I__3273 (
            .O(N__23601),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    Odrv4 I__3272 (
            .O(N__23598),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    InMux I__3271 (
            .O(N__23591),
            .I(N__23586));
    InMux I__3270 (
            .O(N__23590),
            .I(N__23583));
    InMux I__3269 (
            .O(N__23589),
            .I(N__23580));
    LocalMux I__3268 (
            .O(N__23586),
            .I(N__23576));
    LocalMux I__3267 (
            .O(N__23583),
            .I(N__23571));
    LocalMux I__3266 (
            .O(N__23580),
            .I(N__23571));
    InMux I__3265 (
            .O(N__23579),
            .I(N__23568));
    Span4Mux_v I__3264 (
            .O(N__23576),
            .I(N__23565));
    Span4Mux_v I__3263 (
            .O(N__23571),
            .I(N__23562));
    LocalMux I__3262 (
            .O(N__23568),
            .I(N__23559));
    Span4Mux_v I__3261 (
            .O(N__23565),
            .I(N__23556));
    Span4Mux_h I__3260 (
            .O(N__23562),
            .I(N__23551));
    Span4Mux_v I__3259 (
            .O(N__23559),
            .I(N__23551));
    Odrv4 I__3258 (
            .O(N__23556),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    Odrv4 I__3257 (
            .O(N__23551),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    CascadeMux I__3256 (
            .O(N__23546),
            .I(N__23543));
    InMux I__3255 (
            .O(N__23543),
            .I(N__23537));
    InMux I__3254 (
            .O(N__23542),
            .I(N__23537));
    LocalMux I__3253 (
            .O(N__23537),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ));
    InMux I__3252 (
            .O(N__23534),
            .I(N__23529));
    InMux I__3251 (
            .O(N__23533),
            .I(N__23526));
    InMux I__3250 (
            .O(N__23532),
            .I(N__23523));
    LocalMux I__3249 (
            .O(N__23529),
            .I(N__23520));
    LocalMux I__3248 (
            .O(N__23526),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    LocalMux I__3247 (
            .O(N__23523),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    Odrv4 I__3246 (
            .O(N__23520),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    InMux I__3245 (
            .O(N__23513),
            .I(N__23507));
    InMux I__3244 (
            .O(N__23512),
            .I(N__23504));
    InMux I__3243 (
            .O(N__23511),
            .I(N__23499));
    InMux I__3242 (
            .O(N__23510),
            .I(N__23499));
    LocalMux I__3241 (
            .O(N__23507),
            .I(N__23496));
    LocalMux I__3240 (
            .O(N__23504),
            .I(N__23493));
    LocalMux I__3239 (
            .O(N__23499),
            .I(N__23490));
    Span4Mux_v I__3238 (
            .O(N__23496),
            .I(N__23487));
    Span4Mux_v I__3237 (
            .O(N__23493),
            .I(N__23484));
    Span4Mux_h I__3236 (
            .O(N__23490),
            .I(N__23481));
    Odrv4 I__3235 (
            .O(N__23487),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    Odrv4 I__3234 (
            .O(N__23484),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    Odrv4 I__3233 (
            .O(N__23481),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    InMux I__3232 (
            .O(N__23474),
            .I(N__23471));
    LocalMux I__3231 (
            .O(N__23471),
            .I(N__23468));
    Odrv4 I__3230 (
            .O(N__23468),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ));
    InMux I__3229 (
            .O(N__23465),
            .I(N__23460));
    InMux I__3228 (
            .O(N__23464),
            .I(N__23457));
    InMux I__3227 (
            .O(N__23463),
            .I(N__23454));
    LocalMux I__3226 (
            .O(N__23460),
            .I(N__23449));
    LocalMux I__3225 (
            .O(N__23457),
            .I(N__23449));
    LocalMux I__3224 (
            .O(N__23454),
            .I(N__23446));
    Odrv4 I__3223 (
            .O(N__23449),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    Odrv4 I__3222 (
            .O(N__23446),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    InMux I__3221 (
            .O(N__23441),
            .I(N__23436));
    InMux I__3220 (
            .O(N__23440),
            .I(N__23433));
    CascadeMux I__3219 (
            .O(N__23439),
            .I(N__23429));
    LocalMux I__3218 (
            .O(N__23436),
            .I(N__23426));
    LocalMux I__3217 (
            .O(N__23433),
            .I(N__23423));
    InMux I__3216 (
            .O(N__23432),
            .I(N__23420));
    InMux I__3215 (
            .O(N__23429),
            .I(N__23417));
    Span4Mux_h I__3214 (
            .O(N__23426),
            .I(N__23412));
    Span4Mux_h I__3213 (
            .O(N__23423),
            .I(N__23412));
    LocalMux I__3212 (
            .O(N__23420),
            .I(N__23409));
    LocalMux I__3211 (
            .O(N__23417),
            .I(N__23406));
    Span4Mux_v I__3210 (
            .O(N__23412),
            .I(N__23403));
    Span4Mux_v I__3209 (
            .O(N__23409),
            .I(N__23400));
    Span4Mux_h I__3208 (
            .O(N__23406),
            .I(N__23397));
    Span4Mux_v I__3207 (
            .O(N__23403),
            .I(N__23392));
    Span4Mux_v I__3206 (
            .O(N__23400),
            .I(N__23392));
    Span4Mux_v I__3205 (
            .O(N__23397),
            .I(N__23389));
    Odrv4 I__3204 (
            .O(N__23392),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    Odrv4 I__3203 (
            .O(N__23389),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    InMux I__3202 (
            .O(N__23384),
            .I(N__23381));
    LocalMux I__3201 (
            .O(N__23381),
            .I(N__23376));
    InMux I__3200 (
            .O(N__23380),
            .I(N__23373));
    InMux I__3199 (
            .O(N__23379),
            .I(N__23370));
    Span4Mux_v I__3198 (
            .O(N__23376),
            .I(N__23365));
    LocalMux I__3197 (
            .O(N__23373),
            .I(N__23365));
    LocalMux I__3196 (
            .O(N__23370),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    Odrv4 I__3195 (
            .O(N__23365),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    InMux I__3194 (
            .O(N__23360),
            .I(N__23354));
    InMux I__3193 (
            .O(N__23359),
            .I(N__23354));
    LocalMux I__3192 (
            .O(N__23354),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    CascadeMux I__3191 (
            .O(N__23351),
            .I(N__23347));
    InMux I__3190 (
            .O(N__23350),
            .I(N__23342));
    InMux I__3189 (
            .O(N__23347),
            .I(N__23342));
    LocalMux I__3188 (
            .O(N__23342),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    InMux I__3187 (
            .O(N__23339),
            .I(N__23336));
    LocalMux I__3186 (
            .O(N__23336),
            .I(N__23332));
    InMux I__3185 (
            .O(N__23335),
            .I(N__23329));
    Odrv4 I__3184 (
            .O(N__23332),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ));
    LocalMux I__3183 (
            .O(N__23329),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ));
    InMux I__3182 (
            .O(N__23324),
            .I(N__23321));
    LocalMux I__3181 (
            .O(N__23321),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ));
    CascadeMux I__3180 (
            .O(N__23318),
            .I(N__23315));
    InMux I__3179 (
            .O(N__23315),
            .I(N__23312));
    LocalMux I__3178 (
            .O(N__23312),
            .I(N__23309));
    Span4Mux_h I__3177 (
            .O(N__23309),
            .I(N__23306));
    Odrv4 I__3176 (
            .O(N__23306),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ));
    InMux I__3175 (
            .O(N__23303),
            .I(N__23300));
    LocalMux I__3174 (
            .O(N__23300),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ));
    CascadeMux I__3173 (
            .O(N__23297),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ));
    InMux I__3172 (
            .O(N__23294),
            .I(N__23289));
    InMux I__3171 (
            .O(N__23293),
            .I(N__23286));
    InMux I__3170 (
            .O(N__23292),
            .I(N__23283));
    LocalMux I__3169 (
            .O(N__23289),
            .I(N__23277));
    LocalMux I__3168 (
            .O(N__23286),
            .I(N__23277));
    LocalMux I__3167 (
            .O(N__23283),
            .I(N__23274));
    InMux I__3166 (
            .O(N__23282),
            .I(N__23271));
    Span4Mux_s3_v I__3165 (
            .O(N__23277),
            .I(N__23268));
    Span4Mux_s3_v I__3164 (
            .O(N__23274),
            .I(N__23265));
    LocalMux I__3163 (
            .O(N__23271),
            .I(N__23262));
    Span4Mux_v I__3162 (
            .O(N__23268),
            .I(N__23259));
    Span4Mux_v I__3161 (
            .O(N__23265),
            .I(N__23254));
    Span4Mux_h I__3160 (
            .O(N__23262),
            .I(N__23254));
    Odrv4 I__3159 (
            .O(N__23259),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    Odrv4 I__3158 (
            .O(N__23254),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    InMux I__3157 (
            .O(N__23249),
            .I(N__23246));
    LocalMux I__3156 (
            .O(N__23246),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ));
    InMux I__3155 (
            .O(N__23243),
            .I(N__23240));
    LocalMux I__3154 (
            .O(N__23240),
            .I(N__23236));
    InMux I__3153 (
            .O(N__23239),
            .I(N__23231));
    Span4Mux_h I__3152 (
            .O(N__23236),
            .I(N__23228));
    InMux I__3151 (
            .O(N__23235),
            .I(N__23223));
    InMux I__3150 (
            .O(N__23234),
            .I(N__23223));
    LocalMux I__3149 (
            .O(N__23231),
            .I(N__23220));
    Odrv4 I__3148 (
            .O(N__23228),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    LocalMux I__3147 (
            .O(N__23223),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    Odrv4 I__3146 (
            .O(N__23220),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    InMux I__3145 (
            .O(N__23213),
            .I(N__23209));
    InMux I__3144 (
            .O(N__23212),
            .I(N__23206));
    LocalMux I__3143 (
            .O(N__23209),
            .I(elapsed_time_ns_1_RNIK63T9_0_8));
    LocalMux I__3142 (
            .O(N__23206),
            .I(elapsed_time_ns_1_RNIK63T9_0_8));
    CascadeMux I__3141 (
            .O(N__23201),
            .I(N__23198));
    InMux I__3140 (
            .O(N__23198),
            .I(N__23194));
    InMux I__3139 (
            .O(N__23197),
            .I(N__23191));
    LocalMux I__3138 (
            .O(N__23194),
            .I(N__23188));
    LocalMux I__3137 (
            .O(N__23191),
            .I(N__23185));
    Odrv4 I__3136 (
            .O(N__23188),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ));
    Odrv12 I__3135 (
            .O(N__23185),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ));
    InMux I__3134 (
            .O(N__23180),
            .I(N__23175));
    InMux I__3133 (
            .O(N__23179),
            .I(N__23172));
    InMux I__3132 (
            .O(N__23178),
            .I(N__23169));
    LocalMux I__3131 (
            .O(N__23175),
            .I(N__23166));
    LocalMux I__3130 (
            .O(N__23172),
            .I(N__23163));
    LocalMux I__3129 (
            .O(N__23169),
            .I(N__23159));
    Span4Mux_v I__3128 (
            .O(N__23166),
            .I(N__23154));
    Span4Mux_v I__3127 (
            .O(N__23163),
            .I(N__23154));
    InMux I__3126 (
            .O(N__23162),
            .I(N__23151));
    Span4Mux_v I__3125 (
            .O(N__23159),
            .I(N__23148));
    Span4Mux_v I__3124 (
            .O(N__23154),
            .I(N__23145));
    LocalMux I__3123 (
            .O(N__23151),
            .I(N__23142));
    Odrv4 I__3122 (
            .O(N__23148),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    Odrv4 I__3121 (
            .O(N__23145),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    Odrv4 I__3120 (
            .O(N__23142),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    InMux I__3119 (
            .O(N__23135),
            .I(N__23130));
    InMux I__3118 (
            .O(N__23134),
            .I(N__23127));
    InMux I__3117 (
            .O(N__23133),
            .I(N__23124));
    LocalMux I__3116 (
            .O(N__23130),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    LocalMux I__3115 (
            .O(N__23127),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    LocalMux I__3114 (
            .O(N__23124),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    InMux I__3113 (
            .O(N__23117),
            .I(N__23112));
    InMux I__3112 (
            .O(N__23116),
            .I(N__23109));
    InMux I__3111 (
            .O(N__23115),
            .I(N__23106));
    LocalMux I__3110 (
            .O(N__23112),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    LocalMux I__3109 (
            .O(N__23109),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    LocalMux I__3108 (
            .O(N__23106),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    InMux I__3107 (
            .O(N__23099),
            .I(N__23094));
    CascadeMux I__3106 (
            .O(N__23098),
            .I(N__23090));
    InMux I__3105 (
            .O(N__23097),
            .I(N__23087));
    LocalMux I__3104 (
            .O(N__23094),
            .I(N__23084));
    InMux I__3103 (
            .O(N__23093),
            .I(N__23081));
    InMux I__3102 (
            .O(N__23090),
            .I(N__23078));
    LocalMux I__3101 (
            .O(N__23087),
            .I(N__23069));
    Span4Mux_h I__3100 (
            .O(N__23084),
            .I(N__23069));
    LocalMux I__3099 (
            .O(N__23081),
            .I(N__23069));
    LocalMux I__3098 (
            .O(N__23078),
            .I(N__23069));
    Odrv4 I__3097 (
            .O(N__23069),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    InMux I__3096 (
            .O(N__23066),
            .I(N__23061));
    InMux I__3095 (
            .O(N__23065),
            .I(N__23058));
    InMux I__3094 (
            .O(N__23064),
            .I(N__23055));
    LocalMux I__3093 (
            .O(N__23061),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    LocalMux I__3092 (
            .O(N__23058),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    LocalMux I__3091 (
            .O(N__23055),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    CascadeMux I__3090 (
            .O(N__23048),
            .I(N__23045));
    InMux I__3089 (
            .O(N__23045),
            .I(N__23042));
    LocalMux I__3088 (
            .O(N__23042),
            .I(N__23036));
    InMux I__3087 (
            .O(N__23041),
            .I(N__23033));
    InMux I__3086 (
            .O(N__23040),
            .I(N__23028));
    InMux I__3085 (
            .O(N__23039),
            .I(N__23028));
    Odrv4 I__3084 (
            .O(N__23036),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    LocalMux I__3083 (
            .O(N__23033),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    LocalMux I__3082 (
            .O(N__23028),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    InMux I__3081 (
            .O(N__23021),
            .I(N__23016));
    InMux I__3080 (
            .O(N__23020),
            .I(N__23013));
    InMux I__3079 (
            .O(N__23019),
            .I(N__23010));
    LocalMux I__3078 (
            .O(N__23016),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    LocalMux I__3077 (
            .O(N__23013),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    LocalMux I__3076 (
            .O(N__23010),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    InMux I__3075 (
            .O(N__23003),
            .I(N__23000));
    LocalMux I__3074 (
            .O(N__23000),
            .I(N__22994));
    InMux I__3073 (
            .O(N__22999),
            .I(N__22991));
    InMux I__3072 (
            .O(N__22998),
            .I(N__22986));
    InMux I__3071 (
            .O(N__22997),
            .I(N__22986));
    Span4Mux_h I__3070 (
            .O(N__22994),
            .I(N__22979));
    LocalMux I__3069 (
            .O(N__22991),
            .I(N__22979));
    LocalMux I__3068 (
            .O(N__22986),
            .I(N__22979));
    Odrv4 I__3067 (
            .O(N__22979),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    InMux I__3066 (
            .O(N__22976),
            .I(N__22973));
    LocalMux I__3065 (
            .O(N__22973),
            .I(N__22968));
    InMux I__3064 (
            .O(N__22972),
            .I(N__22965));
    InMux I__3063 (
            .O(N__22971),
            .I(N__22962));
    Span4Mux_h I__3062 (
            .O(N__22968),
            .I(N__22957));
    LocalMux I__3061 (
            .O(N__22965),
            .I(N__22957));
    LocalMux I__3060 (
            .O(N__22962),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    Odrv4 I__3059 (
            .O(N__22957),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    InMux I__3058 (
            .O(N__22952),
            .I(N__22949));
    LocalMux I__3057 (
            .O(N__22949),
            .I(N__22945));
    InMux I__3056 (
            .O(N__22948),
            .I(N__22941));
    Span4Mux_h I__3055 (
            .O(N__22945),
            .I(N__22938));
    InMux I__3054 (
            .O(N__22944),
            .I(N__22935));
    LocalMux I__3053 (
            .O(N__22941),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    Odrv4 I__3052 (
            .O(N__22938),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    LocalMux I__3051 (
            .O(N__22935),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    InMux I__3050 (
            .O(N__22928),
            .I(N__22925));
    LocalMux I__3049 (
            .O(N__22925),
            .I(N__22922));
    Span4Mux_h I__3048 (
            .O(N__22922),
            .I(N__22918));
    InMux I__3047 (
            .O(N__22921),
            .I(N__22915));
    Sp12to4 I__3046 (
            .O(N__22918),
            .I(N__22912));
    LocalMux I__3045 (
            .O(N__22915),
            .I(N__22909));
    Span12Mux_v I__3044 (
            .O(N__22912),
            .I(N__22904));
    Span12Mux_v I__3043 (
            .O(N__22909),
            .I(N__22904));
    Odrv12 I__3042 (
            .O(N__22904),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    InMux I__3041 (
            .O(N__22901),
            .I(N__22897));
    InMux I__3040 (
            .O(N__22900),
            .I(N__22894));
    LocalMux I__3039 (
            .O(N__22897),
            .I(N__22891));
    LocalMux I__3038 (
            .O(N__22894),
            .I(N__22888));
    Span4Mux_h I__3037 (
            .O(N__22891),
            .I(N__22885));
    Span4Mux_v I__3036 (
            .O(N__22888),
            .I(N__22882));
    Sp12to4 I__3035 (
            .O(N__22885),
            .I(N__22879));
    Span4Mux_h I__3034 (
            .O(N__22882),
            .I(N__22876));
    Odrv12 I__3033 (
            .O(N__22879),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    Odrv4 I__3032 (
            .O(N__22876),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    InMux I__3031 (
            .O(N__22871),
            .I(N__22868));
    LocalMux I__3030 (
            .O(N__22868),
            .I(N__22864));
    InMux I__3029 (
            .O(N__22867),
            .I(N__22861));
    Span4Mux_h I__3028 (
            .O(N__22864),
            .I(N__22858));
    LocalMux I__3027 (
            .O(N__22861),
            .I(N__22855));
    Sp12to4 I__3026 (
            .O(N__22858),
            .I(N__22850));
    Span12Mux_s7_h I__3025 (
            .O(N__22855),
            .I(N__22850));
    Odrv12 I__3024 (
            .O(N__22850),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    InMux I__3023 (
            .O(N__22847),
            .I(N__22843));
    InMux I__3022 (
            .O(N__22846),
            .I(N__22840));
    LocalMux I__3021 (
            .O(N__22843),
            .I(N__22837));
    LocalMux I__3020 (
            .O(N__22840),
            .I(N__22834));
    Sp12to4 I__3019 (
            .O(N__22837),
            .I(N__22831));
    Span4Mux_s3_h I__3018 (
            .O(N__22834),
            .I(N__22828));
    Span12Mux_v I__3017 (
            .O(N__22831),
            .I(N__22825));
    Span4Mux_h I__3016 (
            .O(N__22828),
            .I(N__22822));
    Odrv12 I__3015 (
            .O(N__22825),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    Odrv4 I__3014 (
            .O(N__22822),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    CascadeMux I__3013 (
            .O(N__22817),
            .I(N__22814));
    InMux I__3012 (
            .O(N__22814),
            .I(N__22811));
    LocalMux I__3011 (
            .O(N__22811),
            .I(N__22808));
    Odrv12 I__3010 (
            .O(N__22808),
            .I(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ));
    InMux I__3009 (
            .O(N__22805),
            .I(N__22801));
    InMux I__3008 (
            .O(N__22804),
            .I(N__22798));
    LocalMux I__3007 (
            .O(N__22801),
            .I(N__22795));
    LocalMux I__3006 (
            .O(N__22798),
            .I(N__22792));
    Span4Mux_h I__3005 (
            .O(N__22795),
            .I(N__22789));
    Span4Mux_s3_h I__3004 (
            .O(N__22792),
            .I(N__22786));
    Sp12to4 I__3003 (
            .O(N__22789),
            .I(N__22783));
    Span4Mux_h I__3002 (
            .O(N__22786),
            .I(N__22780));
    Odrv12 I__3001 (
            .O(N__22783),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    Odrv4 I__3000 (
            .O(N__22780),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    CascadeMux I__2999 (
            .O(N__22775),
            .I(N__22772));
    InMux I__2998 (
            .O(N__22772),
            .I(N__22769));
    LocalMux I__2997 (
            .O(N__22769),
            .I(N__22766));
    Odrv4 I__2996 (
            .O(N__22766),
            .I(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ));
    CascadeMux I__2995 (
            .O(N__22763),
            .I(N__22760));
    InMux I__2994 (
            .O(N__22760),
            .I(N__22757));
    LocalMux I__2993 (
            .O(N__22757),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ));
    InMux I__2992 (
            .O(N__22754),
            .I(N__22751));
    LocalMux I__2991 (
            .O(N__22751),
            .I(N__22748));
    Odrv4 I__2990 (
            .O(N__22748),
            .I(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ));
    InMux I__2989 (
            .O(N__22745),
            .I(N__22742));
    LocalMux I__2988 (
            .O(N__22742),
            .I(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ));
    InMux I__2987 (
            .O(N__22739),
            .I(N__22736));
    LocalMux I__2986 (
            .O(N__22736),
            .I(N__22733));
    Odrv12 I__2985 (
            .O(N__22733),
            .I(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ));
    InMux I__2984 (
            .O(N__22730),
            .I(N__22727));
    LocalMux I__2983 (
            .O(N__22727),
            .I(N__22724));
    Odrv4 I__2982 (
            .O(N__22724),
            .I(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ));
    CascadeMux I__2981 (
            .O(N__22721),
            .I(N__22718));
    InMux I__2980 (
            .O(N__22718),
            .I(N__22715));
    LocalMux I__2979 (
            .O(N__22715),
            .I(N__22712));
    Odrv4 I__2978 (
            .O(N__22712),
            .I(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ));
    CascadeMux I__2977 (
            .O(N__22709),
            .I(N__22706));
    InMux I__2976 (
            .O(N__22706),
            .I(N__22703));
    LocalMux I__2975 (
            .O(N__22703),
            .I(N__22700));
    Odrv4 I__2974 (
            .O(N__22700),
            .I(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ));
    InMux I__2973 (
            .O(N__22697),
            .I(\current_shift_inst.un10_control_input_cry_30 ));
    InMux I__2972 (
            .O(N__22694),
            .I(N__22691));
    LocalMux I__2971 (
            .O(N__22691),
            .I(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ));
    CascadeMux I__2970 (
            .O(N__22688),
            .I(N__22685));
    InMux I__2969 (
            .O(N__22685),
            .I(N__22682));
    LocalMux I__2968 (
            .O(N__22682),
            .I(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ));
    InMux I__2967 (
            .O(N__22679),
            .I(N__22676));
    LocalMux I__2966 (
            .O(N__22676),
            .I(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ));
    InMux I__2965 (
            .O(N__22673),
            .I(N__22670));
    LocalMux I__2964 (
            .O(N__22670),
            .I(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ));
    InMux I__2963 (
            .O(N__22667),
            .I(N__22664));
    LocalMux I__2962 (
            .O(N__22664),
            .I(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ));
    CascadeMux I__2961 (
            .O(N__22661),
            .I(N__22658));
    InMux I__2960 (
            .O(N__22658),
            .I(N__22655));
    LocalMux I__2959 (
            .O(N__22655),
            .I(N__22652));
    Odrv4 I__2958 (
            .O(N__22652),
            .I(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ));
    InMux I__2957 (
            .O(N__22649),
            .I(N__22646));
    LocalMux I__2956 (
            .O(N__22646),
            .I(\current_shift_inst.control_input_axb_3 ));
    CascadeMux I__2955 (
            .O(N__22643),
            .I(N__22640));
    InMux I__2954 (
            .O(N__22640),
            .I(N__22637));
    LocalMux I__2953 (
            .O(N__22637),
            .I(N__22633));
    InMux I__2952 (
            .O(N__22636),
            .I(N__22630));
    Span4Mux_h I__2951 (
            .O(N__22633),
            .I(N__22627));
    LocalMux I__2950 (
            .O(N__22630),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    Odrv4 I__2949 (
            .O(N__22627),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    InMux I__2948 (
            .O(N__22622),
            .I(N__22619));
    LocalMux I__2947 (
            .O(N__22619),
            .I(\current_shift_inst.control_input_axb_7 ));
    InMux I__2946 (
            .O(N__22616),
            .I(N__22613));
    LocalMux I__2945 (
            .O(N__22613),
            .I(N__22610));
    Span4Mux_h I__2944 (
            .O(N__22610),
            .I(N__22607));
    Odrv4 I__2943 (
            .O(N__22607),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ));
    InMux I__2942 (
            .O(N__22604),
            .I(\current_shift_inst.control_input_cry_6 ));
    InMux I__2941 (
            .O(N__22601),
            .I(N__22598));
    LocalMux I__2940 (
            .O(N__22598),
            .I(N__22595));
    Span4Mux_v I__2939 (
            .O(N__22595),
            .I(N__22592));
    Odrv4 I__2938 (
            .O(N__22592),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ));
    InMux I__2937 (
            .O(N__22589),
            .I(bfn_9_15_0_));
    InMux I__2936 (
            .O(N__22586),
            .I(N__22583));
    LocalMux I__2935 (
            .O(N__22583),
            .I(N__22580));
    Span4Mux_v I__2934 (
            .O(N__22580),
            .I(N__22577));
    Odrv4 I__2933 (
            .O(N__22577),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ));
    InMux I__2932 (
            .O(N__22574),
            .I(\current_shift_inst.control_input_cry_8 ));
    InMux I__2931 (
            .O(N__22571),
            .I(N__22568));
    LocalMux I__2930 (
            .O(N__22568),
            .I(N__22565));
    Span4Mux_h I__2929 (
            .O(N__22565),
            .I(N__22562));
    Odrv4 I__2928 (
            .O(N__22562),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ));
    InMux I__2927 (
            .O(N__22559),
            .I(\current_shift_inst.control_input_cry_9 ));
    InMux I__2926 (
            .O(N__22556),
            .I(N__22553));
    LocalMux I__2925 (
            .O(N__22553),
            .I(N__22550));
    Span4Mux_h I__2924 (
            .O(N__22550),
            .I(N__22547));
    Odrv4 I__2923 (
            .O(N__22547),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ));
    InMux I__2922 (
            .O(N__22544),
            .I(\current_shift_inst.control_input_cry_10 ));
    InMux I__2921 (
            .O(N__22541),
            .I(N__22538));
    LocalMux I__2920 (
            .O(N__22538),
            .I(\current_shift_inst.control_input_axb_12 ));
    InMux I__2919 (
            .O(N__22535),
            .I(N__22532));
    LocalMux I__2918 (
            .O(N__22532),
            .I(N__22529));
    Span4Mux_h I__2917 (
            .O(N__22529),
            .I(N__22526));
    Odrv4 I__2916 (
            .O(N__22526),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ));
    InMux I__2915 (
            .O(N__22523),
            .I(\current_shift_inst.control_input_cry_11 ));
    InMux I__2914 (
            .O(N__22520),
            .I(\current_shift_inst.control_input_cry_12 ));
    InMux I__2913 (
            .O(N__22517),
            .I(N__22514));
    LocalMux I__2912 (
            .O(N__22514),
            .I(N__22511));
    Span4Mux_h I__2911 (
            .O(N__22511),
            .I(N__22507));
    InMux I__2910 (
            .O(N__22510),
            .I(N__22504));
    Odrv4 I__2909 (
            .O(N__22507),
            .I(\current_shift_inst.control_input_31 ));
    LocalMux I__2908 (
            .O(N__22504),
            .I(\current_shift_inst.control_input_31 ));
    InMux I__2907 (
            .O(N__22499),
            .I(N__22496));
    LocalMux I__2906 (
            .O(N__22496),
            .I(\current_shift_inst.control_input_axb_1 ));
    InMux I__2905 (
            .O(N__22493),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ));
    InMux I__2904 (
            .O(N__22490),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30 ));
    InMux I__2903 (
            .O(N__22487),
            .I(N__22484));
    LocalMux I__2902 (
            .O(N__22484),
            .I(N__22481));
    Span4Mux_v I__2901 (
            .O(N__22481),
            .I(N__22478));
    Odrv4 I__2900 (
            .O(N__22478),
            .I(\current_shift_inst.control_input_18 ));
    InMux I__2899 (
            .O(N__22475),
            .I(N__22472));
    LocalMux I__2898 (
            .O(N__22472),
            .I(N__22469));
    Span4Mux_v I__2897 (
            .O(N__22469),
            .I(N__22466));
    Odrv4 I__2896 (
            .O(N__22466),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ));
    InMux I__2895 (
            .O(N__22463),
            .I(\current_shift_inst.control_input_cry_0 ));
    InMux I__2894 (
            .O(N__22460),
            .I(N__22457));
    LocalMux I__2893 (
            .O(N__22457),
            .I(\current_shift_inst.control_input_axb_2 ));
    InMux I__2892 (
            .O(N__22454),
            .I(N__22451));
    LocalMux I__2891 (
            .O(N__22451),
            .I(N__22448));
    Span4Mux_h I__2890 (
            .O(N__22448),
            .I(N__22445));
    Odrv4 I__2889 (
            .O(N__22445),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ));
    InMux I__2888 (
            .O(N__22442),
            .I(\current_shift_inst.control_input_cry_1 ));
    InMux I__2887 (
            .O(N__22439),
            .I(N__22436));
    LocalMux I__2886 (
            .O(N__22436),
            .I(N__22433));
    Span4Mux_h I__2885 (
            .O(N__22433),
            .I(N__22430));
    Odrv4 I__2884 (
            .O(N__22430),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ));
    InMux I__2883 (
            .O(N__22427),
            .I(\current_shift_inst.control_input_cry_2 ));
    InMux I__2882 (
            .O(N__22424),
            .I(N__22421));
    LocalMux I__2881 (
            .O(N__22421),
            .I(\current_shift_inst.control_input_axb_4 ));
    InMux I__2880 (
            .O(N__22418),
            .I(N__22415));
    LocalMux I__2879 (
            .O(N__22415),
            .I(N__22412));
    Span4Mux_h I__2878 (
            .O(N__22412),
            .I(N__22409));
    Odrv4 I__2877 (
            .O(N__22409),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ));
    InMux I__2876 (
            .O(N__22406),
            .I(\current_shift_inst.control_input_cry_3 ));
    InMux I__2875 (
            .O(N__22403),
            .I(N__22400));
    LocalMux I__2874 (
            .O(N__22400),
            .I(\current_shift_inst.control_input_axb_5 ));
    InMux I__2873 (
            .O(N__22397),
            .I(N__22394));
    LocalMux I__2872 (
            .O(N__22394),
            .I(N__22391));
    Span4Mux_h I__2871 (
            .O(N__22391),
            .I(N__22388));
    Odrv4 I__2870 (
            .O(N__22388),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ));
    InMux I__2869 (
            .O(N__22385),
            .I(\current_shift_inst.control_input_cry_4 ));
    InMux I__2868 (
            .O(N__22382),
            .I(N__22379));
    LocalMux I__2867 (
            .O(N__22379),
            .I(\current_shift_inst.control_input_axb_6 ));
    InMux I__2866 (
            .O(N__22376),
            .I(N__22373));
    LocalMux I__2865 (
            .O(N__22373),
            .I(N__22370));
    Span4Mux_h I__2864 (
            .O(N__22370),
            .I(N__22367));
    Odrv4 I__2863 (
            .O(N__22367),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ));
    InMux I__2862 (
            .O(N__22364),
            .I(\current_shift_inst.control_input_cry_5 ));
    InMux I__2861 (
            .O(N__22361),
            .I(N__22358));
    LocalMux I__2860 (
            .O(N__22358),
            .I(N__22355));
    Span12Mux_v I__2859 (
            .O(N__22355),
            .I(N__22352));
    Odrv12 I__2858 (
            .O(N__22352),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ));
    CascadeMux I__2857 (
            .O(N__22349),
            .I(N__22346));
    InMux I__2856 (
            .O(N__22346),
            .I(N__22343));
    LocalMux I__2855 (
            .O(N__22343),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ));
    InMux I__2854 (
            .O(N__22340),
            .I(N__22337));
    LocalMux I__2853 (
            .O(N__22337),
            .I(N__22334));
    Odrv12 I__2852 (
            .O(N__22334),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt18 ));
    CascadeMux I__2851 (
            .O(N__22331),
            .I(N__22328));
    InMux I__2850 (
            .O(N__22328),
            .I(N__22325));
    LocalMux I__2849 (
            .O(N__22325),
            .I(N__22322));
    Span4Mux_h I__2848 (
            .O(N__22322),
            .I(N__22319));
    Span4Mux_v I__2847 (
            .O(N__22319),
            .I(N__22316));
    Odrv4 I__2846 (
            .O(N__22316),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ));
    InMux I__2845 (
            .O(N__22313),
            .I(N__22310));
    LocalMux I__2844 (
            .O(N__22310),
            .I(N__22307));
    Odrv12 I__2843 (
            .O(N__22307),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ));
    CascadeMux I__2842 (
            .O(N__22304),
            .I(N__22301));
    InMux I__2841 (
            .O(N__22301),
            .I(N__22298));
    LocalMux I__2840 (
            .O(N__22298),
            .I(N__22295));
    Span4Mux_v I__2839 (
            .O(N__22295),
            .I(N__22292));
    Odrv4 I__2838 (
            .O(N__22292),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt20 ));
    InMux I__2837 (
            .O(N__22289),
            .I(N__22286));
    LocalMux I__2836 (
            .O(N__22286),
            .I(N__22283));
    Span4Mux_h I__2835 (
            .O(N__22283),
            .I(N__22280));
    Odrv4 I__2834 (
            .O(N__22280),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt22 ));
    CascadeMux I__2833 (
            .O(N__22277),
            .I(N__22274));
    InMux I__2832 (
            .O(N__22274),
            .I(N__22271));
    LocalMux I__2831 (
            .O(N__22271),
            .I(N__22268));
    Span4Mux_h I__2830 (
            .O(N__22268),
            .I(N__22265));
    Odrv4 I__2829 (
            .O(N__22265),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ));
    InMux I__2828 (
            .O(N__22262),
            .I(N__22259));
    LocalMux I__2827 (
            .O(N__22259),
            .I(N__22256));
    Odrv12 I__2826 (
            .O(N__22256),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ));
    CascadeMux I__2825 (
            .O(N__22253),
            .I(N__22250));
    InMux I__2824 (
            .O(N__22250),
            .I(N__22247));
    LocalMux I__2823 (
            .O(N__22247),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ));
    InMux I__2822 (
            .O(N__22244),
            .I(N__22241));
    LocalMux I__2821 (
            .O(N__22241),
            .I(N__22238));
    Odrv4 I__2820 (
            .O(N__22238),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ));
    CascadeMux I__2819 (
            .O(N__22235),
            .I(N__22232));
    InMux I__2818 (
            .O(N__22232),
            .I(N__22229));
    LocalMux I__2817 (
            .O(N__22229),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ));
    CascadeMux I__2816 (
            .O(N__22226),
            .I(N__22223));
    InMux I__2815 (
            .O(N__22223),
            .I(N__22220));
    LocalMux I__2814 (
            .O(N__22220),
            .I(N__22217));
    Odrv4 I__2813 (
            .O(N__22217),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ));
    InMux I__2812 (
            .O(N__22214),
            .I(N__22211));
    LocalMux I__2811 (
            .O(N__22211),
            .I(N__22208));
    Span4Mux_h I__2810 (
            .O(N__22208),
            .I(N__22205));
    Odrv4 I__2809 (
            .O(N__22205),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ));
    InMux I__2808 (
            .O(N__22202),
            .I(N__22199));
    LocalMux I__2807 (
            .O(N__22199),
            .I(N__22196));
    Odrv4 I__2806 (
            .O(N__22196),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ));
    CascadeMux I__2805 (
            .O(N__22193),
            .I(N__22190));
    InMux I__2804 (
            .O(N__22190),
            .I(N__22187));
    LocalMux I__2803 (
            .O(N__22187),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ));
    InMux I__2802 (
            .O(N__22184),
            .I(N__22181));
    LocalMux I__2801 (
            .O(N__22181),
            .I(N__22178));
    Odrv12 I__2800 (
            .O(N__22178),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ));
    CascadeMux I__2799 (
            .O(N__22175),
            .I(N__22172));
    InMux I__2798 (
            .O(N__22172),
            .I(N__22169));
    LocalMux I__2797 (
            .O(N__22169),
            .I(N__22166));
    Odrv4 I__2796 (
            .O(N__22166),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ));
    InMux I__2795 (
            .O(N__22163),
            .I(N__22160));
    LocalMux I__2794 (
            .O(N__22160),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ));
    CascadeMux I__2793 (
            .O(N__22157),
            .I(N__22154));
    InMux I__2792 (
            .O(N__22154),
            .I(N__22151));
    LocalMux I__2791 (
            .O(N__22151),
            .I(N__22148));
    Odrv4 I__2790 (
            .O(N__22148),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ));
    InMux I__2789 (
            .O(N__22145),
            .I(N__22142));
    LocalMux I__2788 (
            .O(N__22142),
            .I(N__22139));
    Span4Mux_v I__2787 (
            .O(N__22139),
            .I(N__22136));
    Odrv4 I__2786 (
            .O(N__22136),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ));
    CascadeMux I__2785 (
            .O(N__22133),
            .I(N__22130));
    InMux I__2784 (
            .O(N__22130),
            .I(N__22127));
    LocalMux I__2783 (
            .O(N__22127),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ));
    CascadeMux I__2782 (
            .O(N__22124),
            .I(elapsed_time_ns_1_RNIK63T9_0_8_cascade_));
    CascadeMux I__2781 (
            .O(N__22121),
            .I(N__22118));
    InMux I__2780 (
            .O(N__22118),
            .I(N__22115));
    LocalMux I__2779 (
            .O(N__22115),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ));
    InMux I__2778 (
            .O(N__22112),
            .I(N__22109));
    LocalMux I__2777 (
            .O(N__22109),
            .I(N__22106));
    Odrv4 I__2776 (
            .O(N__22106),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ));
    CascadeMux I__2775 (
            .O(N__22103),
            .I(N__22100));
    InMux I__2774 (
            .O(N__22100),
            .I(N__22097));
    LocalMux I__2773 (
            .O(N__22097),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ));
    CascadeMux I__2772 (
            .O(N__22094),
            .I(N__22091));
    InMux I__2771 (
            .O(N__22091),
            .I(N__22088));
    LocalMux I__2770 (
            .O(N__22088),
            .I(N__22085));
    Odrv4 I__2769 (
            .O(N__22085),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ));
    InMux I__2768 (
            .O(N__22082),
            .I(N__22079));
    LocalMux I__2767 (
            .O(N__22079),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ));
    InMux I__2766 (
            .O(N__22076),
            .I(N__22073));
    LocalMux I__2765 (
            .O(N__22073),
            .I(N__22070));
    Odrv4 I__2764 (
            .O(N__22070),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ));
    CascadeMux I__2763 (
            .O(N__22067),
            .I(N__22064));
    InMux I__2762 (
            .O(N__22064),
            .I(N__22061));
    LocalMux I__2761 (
            .O(N__22061),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ));
    InMux I__2760 (
            .O(N__22058),
            .I(N__22055));
    LocalMux I__2759 (
            .O(N__22055),
            .I(N__22052));
    Span4Mux_v I__2758 (
            .O(N__22052),
            .I(N__22049));
    Odrv4 I__2757 (
            .O(N__22049),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ));
    CascadeMux I__2756 (
            .O(N__22046),
            .I(N__22043));
    InMux I__2755 (
            .O(N__22043),
            .I(N__22040));
    LocalMux I__2754 (
            .O(N__22040),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ));
    InMux I__2753 (
            .O(N__22037),
            .I(N__22034));
    LocalMux I__2752 (
            .O(N__22034),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ));
    CascadeMux I__2751 (
            .O(N__22031),
            .I(N__22028));
    InMux I__2750 (
            .O(N__22028),
            .I(N__22025));
    LocalMux I__2749 (
            .O(N__22025),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ));
    InMux I__2748 (
            .O(N__22022),
            .I(N__22018));
    InMux I__2747 (
            .O(N__22021),
            .I(N__22015));
    LocalMux I__2746 (
            .O(N__22018),
            .I(N__22012));
    LocalMux I__2745 (
            .O(N__22015),
            .I(N__22009));
    Odrv4 I__2744 (
            .O(N__22012),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ));
    Odrv4 I__2743 (
            .O(N__22009),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ));
    InMux I__2742 (
            .O(N__22004),
            .I(N__22001));
    LocalMux I__2741 (
            .O(N__22001),
            .I(N__21997));
    InMux I__2740 (
            .O(N__22000),
            .I(N__21994));
    Span4Mux_h I__2739 (
            .O(N__21997),
            .I(N__21991));
    LocalMux I__2738 (
            .O(N__21994),
            .I(N__21988));
    Odrv4 I__2737 (
            .O(N__21991),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ));
    Odrv4 I__2736 (
            .O(N__21988),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ));
    InMux I__2735 (
            .O(N__21983),
            .I(N__21977));
    InMux I__2734 (
            .O(N__21982),
            .I(N__21977));
    LocalMux I__2733 (
            .O(N__21977),
            .I(N__21974));
    Span4Mux_v I__2732 (
            .O(N__21974),
            .I(N__21971));
    Odrv4 I__2731 (
            .O(N__21971),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ));
    InMux I__2730 (
            .O(N__21968),
            .I(N__21965));
    LocalMux I__2729 (
            .O(N__21965),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ));
    CascadeMux I__2728 (
            .O(N__21962),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21_cascade_ ));
    CascadeMux I__2727 (
            .O(N__21959),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ));
    InMux I__2726 (
            .O(N__21956),
            .I(N__21952));
    InMux I__2725 (
            .O(N__21955),
            .I(N__21948));
    LocalMux I__2724 (
            .O(N__21952),
            .I(N__21945));
    InMux I__2723 (
            .O(N__21951),
            .I(N__21942));
    LocalMux I__2722 (
            .O(N__21948),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    Odrv12 I__2721 (
            .O(N__21945),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__2720 (
            .O(N__21942),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    CascadeMux I__2719 (
            .O(N__21935),
            .I(N__21932));
    InMux I__2718 (
            .O(N__21932),
            .I(N__21929));
    LocalMux I__2717 (
            .O(N__21929),
            .I(N__21924));
    InMux I__2716 (
            .O(N__21928),
            .I(N__21921));
    InMux I__2715 (
            .O(N__21927),
            .I(N__21918));
    Span4Mux_v I__2714 (
            .O(N__21924),
            .I(N__21915));
    LocalMux I__2713 (
            .O(N__21921),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__2712 (
            .O(N__21918),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    Odrv4 I__2711 (
            .O(N__21915),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    InMux I__2710 (
            .O(N__21908),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    InMux I__2709 (
            .O(N__21905),
            .I(N__21901));
    InMux I__2708 (
            .O(N__21904),
            .I(N__21898));
    LocalMux I__2707 (
            .O(N__21901),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    LocalMux I__2706 (
            .O(N__21898),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    IoInMux I__2705 (
            .O(N__21893),
            .I(N__21890));
    LocalMux I__2704 (
            .O(N__21890),
            .I(N__21887));
    Odrv4 I__2703 (
            .O(N__21887),
            .I(s4_phy_c));
    IoInMux I__2702 (
            .O(N__21884),
            .I(N__21881));
    LocalMux I__2701 (
            .O(N__21881),
            .I(GB_BUFFER_clock_output_0_THRU_CO));
    InMux I__2700 (
            .O(N__21878),
            .I(N__21875));
    LocalMux I__2699 (
            .O(N__21875),
            .I(N__21872));
    Odrv4 I__2698 (
            .O(N__21872),
            .I(il_min_comp1_c));
    InMux I__2697 (
            .O(N__21869),
            .I(N__21864));
    InMux I__2696 (
            .O(N__21868),
            .I(N__21861));
    InMux I__2695 (
            .O(N__21867),
            .I(N__21858));
    LocalMux I__2694 (
            .O(N__21864),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    LocalMux I__2693 (
            .O(N__21861),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    LocalMux I__2692 (
            .O(N__21858),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    InMux I__2691 (
            .O(N__21851),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    CascadeMux I__2690 (
            .O(N__21848),
            .I(N__21844));
    InMux I__2689 (
            .O(N__21847),
            .I(N__21840));
    InMux I__2688 (
            .O(N__21844),
            .I(N__21837));
    InMux I__2687 (
            .O(N__21843),
            .I(N__21834));
    LocalMux I__2686 (
            .O(N__21840),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    LocalMux I__2685 (
            .O(N__21837),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    LocalMux I__2684 (
            .O(N__21834),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    InMux I__2683 (
            .O(N__21827),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    CascadeMux I__2682 (
            .O(N__21824),
            .I(N__21820));
    InMux I__2681 (
            .O(N__21823),
            .I(N__21816));
    InMux I__2680 (
            .O(N__21820),
            .I(N__21813));
    InMux I__2679 (
            .O(N__21819),
            .I(N__21810));
    LocalMux I__2678 (
            .O(N__21816),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    LocalMux I__2677 (
            .O(N__21813),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    LocalMux I__2676 (
            .O(N__21810),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    InMux I__2675 (
            .O(N__21803),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    CascadeMux I__2674 (
            .O(N__21800),
            .I(N__21796));
    InMux I__2673 (
            .O(N__21799),
            .I(N__21792));
    InMux I__2672 (
            .O(N__21796),
            .I(N__21789));
    InMux I__2671 (
            .O(N__21795),
            .I(N__21786));
    LocalMux I__2670 (
            .O(N__21792),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    LocalMux I__2669 (
            .O(N__21789),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    LocalMux I__2668 (
            .O(N__21786),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__2667 (
            .O(N__21779),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    CascadeMux I__2666 (
            .O(N__21776),
            .I(N__21772));
    InMux I__2665 (
            .O(N__21775),
            .I(N__21768));
    InMux I__2664 (
            .O(N__21772),
            .I(N__21765));
    InMux I__2663 (
            .O(N__21771),
            .I(N__21762));
    LocalMux I__2662 (
            .O(N__21768),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    LocalMux I__2661 (
            .O(N__21765),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    LocalMux I__2660 (
            .O(N__21762),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    InMux I__2659 (
            .O(N__21755),
            .I(bfn_8_22_0_));
    CascadeMux I__2658 (
            .O(N__21752),
            .I(N__21748));
    InMux I__2657 (
            .O(N__21751),
            .I(N__21744));
    InMux I__2656 (
            .O(N__21748),
            .I(N__21741));
    InMux I__2655 (
            .O(N__21747),
            .I(N__21738));
    LocalMux I__2654 (
            .O(N__21744),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    LocalMux I__2653 (
            .O(N__21741),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    LocalMux I__2652 (
            .O(N__21738),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    InMux I__2651 (
            .O(N__21731),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    CascadeMux I__2650 (
            .O(N__21728),
            .I(N__21724));
    InMux I__2649 (
            .O(N__21727),
            .I(N__21720));
    InMux I__2648 (
            .O(N__21724),
            .I(N__21717));
    InMux I__2647 (
            .O(N__21723),
            .I(N__21714));
    LocalMux I__2646 (
            .O(N__21720),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    LocalMux I__2645 (
            .O(N__21717),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    LocalMux I__2644 (
            .O(N__21714),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__2643 (
            .O(N__21707),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    CascadeMux I__2642 (
            .O(N__21704),
            .I(N__21700));
    InMux I__2641 (
            .O(N__21703),
            .I(N__21696));
    InMux I__2640 (
            .O(N__21700),
            .I(N__21693));
    InMux I__2639 (
            .O(N__21699),
            .I(N__21690));
    LocalMux I__2638 (
            .O(N__21696),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    LocalMux I__2637 (
            .O(N__21693),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    LocalMux I__2636 (
            .O(N__21690),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    InMux I__2635 (
            .O(N__21683),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    InMux I__2634 (
            .O(N__21680),
            .I(N__21676));
    InMux I__2633 (
            .O(N__21679),
            .I(N__21673));
    LocalMux I__2632 (
            .O(N__21676),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    LocalMux I__2631 (
            .O(N__21673),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    InMux I__2630 (
            .O(N__21668),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    CascadeMux I__2629 (
            .O(N__21665),
            .I(N__21661));
    InMux I__2628 (
            .O(N__21664),
            .I(N__21657));
    InMux I__2627 (
            .O(N__21661),
            .I(N__21654));
    InMux I__2626 (
            .O(N__21660),
            .I(N__21651));
    LocalMux I__2625 (
            .O(N__21657),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    LocalMux I__2624 (
            .O(N__21654),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    LocalMux I__2623 (
            .O(N__21651),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    InMux I__2622 (
            .O(N__21644),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    CascadeMux I__2621 (
            .O(N__21641),
            .I(N__21637));
    InMux I__2620 (
            .O(N__21640),
            .I(N__21633));
    InMux I__2619 (
            .O(N__21637),
            .I(N__21630));
    InMux I__2618 (
            .O(N__21636),
            .I(N__21627));
    LocalMux I__2617 (
            .O(N__21633),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    LocalMux I__2616 (
            .O(N__21630),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    LocalMux I__2615 (
            .O(N__21627),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    InMux I__2614 (
            .O(N__21620),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    CascadeMux I__2613 (
            .O(N__21617),
            .I(N__21613));
    InMux I__2612 (
            .O(N__21616),
            .I(N__21609));
    InMux I__2611 (
            .O(N__21613),
            .I(N__21606));
    InMux I__2610 (
            .O(N__21612),
            .I(N__21603));
    LocalMux I__2609 (
            .O(N__21609),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    LocalMux I__2608 (
            .O(N__21606),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    LocalMux I__2607 (
            .O(N__21603),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    InMux I__2606 (
            .O(N__21596),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    CascadeMux I__2605 (
            .O(N__21593),
            .I(N__21589));
    InMux I__2604 (
            .O(N__21592),
            .I(N__21585));
    InMux I__2603 (
            .O(N__21589),
            .I(N__21582));
    InMux I__2602 (
            .O(N__21588),
            .I(N__21579));
    LocalMux I__2601 (
            .O(N__21585),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    LocalMux I__2600 (
            .O(N__21582),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    LocalMux I__2599 (
            .O(N__21579),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__2598 (
            .O(N__21572),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    CascadeMux I__2597 (
            .O(N__21569),
            .I(N__21565));
    InMux I__2596 (
            .O(N__21568),
            .I(N__21561));
    InMux I__2595 (
            .O(N__21565),
            .I(N__21558));
    InMux I__2594 (
            .O(N__21564),
            .I(N__21555));
    LocalMux I__2593 (
            .O(N__21561),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    LocalMux I__2592 (
            .O(N__21558),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    LocalMux I__2591 (
            .O(N__21555),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    InMux I__2590 (
            .O(N__21548),
            .I(bfn_8_21_0_));
    CascadeMux I__2589 (
            .O(N__21545),
            .I(N__21541));
    InMux I__2588 (
            .O(N__21544),
            .I(N__21537));
    InMux I__2587 (
            .O(N__21541),
            .I(N__21534));
    InMux I__2586 (
            .O(N__21540),
            .I(N__21531));
    LocalMux I__2585 (
            .O(N__21537),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    LocalMux I__2584 (
            .O(N__21534),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    LocalMux I__2583 (
            .O(N__21531),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    InMux I__2582 (
            .O(N__21524),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    CascadeMux I__2581 (
            .O(N__21521),
            .I(N__21517));
    InMux I__2580 (
            .O(N__21520),
            .I(N__21513));
    InMux I__2579 (
            .O(N__21517),
            .I(N__21510));
    InMux I__2578 (
            .O(N__21516),
            .I(N__21507));
    LocalMux I__2577 (
            .O(N__21513),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    LocalMux I__2576 (
            .O(N__21510),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    LocalMux I__2575 (
            .O(N__21507),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    InMux I__2574 (
            .O(N__21500),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    CascadeMux I__2573 (
            .O(N__21497),
            .I(N__21493));
    InMux I__2572 (
            .O(N__21496),
            .I(N__21489));
    InMux I__2571 (
            .O(N__21493),
            .I(N__21486));
    InMux I__2570 (
            .O(N__21492),
            .I(N__21483));
    LocalMux I__2569 (
            .O(N__21489),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    LocalMux I__2568 (
            .O(N__21486),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    LocalMux I__2567 (
            .O(N__21483),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    InMux I__2566 (
            .O(N__21476),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    CascadeMux I__2565 (
            .O(N__21473),
            .I(N__21469));
    InMux I__2564 (
            .O(N__21472),
            .I(N__21465));
    InMux I__2563 (
            .O(N__21469),
            .I(N__21462));
    InMux I__2562 (
            .O(N__21468),
            .I(N__21459));
    LocalMux I__2561 (
            .O(N__21465),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    LocalMux I__2560 (
            .O(N__21462),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    LocalMux I__2559 (
            .O(N__21459),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    CascadeMux I__2558 (
            .O(N__21452),
            .I(N__21448));
    InMux I__2557 (
            .O(N__21451),
            .I(N__21444));
    InMux I__2556 (
            .O(N__21448),
            .I(N__21441));
    InMux I__2555 (
            .O(N__21447),
            .I(N__21438));
    LocalMux I__2554 (
            .O(N__21444),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    LocalMux I__2553 (
            .O(N__21441),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    LocalMux I__2552 (
            .O(N__21438),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    InMux I__2551 (
            .O(N__21431),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    CascadeMux I__2550 (
            .O(N__21428),
            .I(N__21424));
    InMux I__2549 (
            .O(N__21427),
            .I(N__21420));
    InMux I__2548 (
            .O(N__21424),
            .I(N__21417));
    InMux I__2547 (
            .O(N__21423),
            .I(N__21414));
    LocalMux I__2546 (
            .O(N__21420),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    LocalMux I__2545 (
            .O(N__21417),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    LocalMux I__2544 (
            .O(N__21414),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    InMux I__2543 (
            .O(N__21407),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    CascadeMux I__2542 (
            .O(N__21404),
            .I(N__21400));
    InMux I__2541 (
            .O(N__21403),
            .I(N__21396));
    InMux I__2540 (
            .O(N__21400),
            .I(N__21393));
    InMux I__2539 (
            .O(N__21399),
            .I(N__21390));
    LocalMux I__2538 (
            .O(N__21396),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    LocalMux I__2537 (
            .O(N__21393),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    LocalMux I__2536 (
            .O(N__21390),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    InMux I__2535 (
            .O(N__21383),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    CascadeMux I__2534 (
            .O(N__21380),
            .I(N__21376));
    InMux I__2533 (
            .O(N__21379),
            .I(N__21372));
    InMux I__2532 (
            .O(N__21376),
            .I(N__21369));
    InMux I__2531 (
            .O(N__21375),
            .I(N__21366));
    LocalMux I__2530 (
            .O(N__21372),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    LocalMux I__2529 (
            .O(N__21369),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    LocalMux I__2528 (
            .O(N__21366),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    InMux I__2527 (
            .O(N__21359),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    CascadeMux I__2526 (
            .O(N__21356),
            .I(N__21352));
    InMux I__2525 (
            .O(N__21355),
            .I(N__21348));
    InMux I__2524 (
            .O(N__21352),
            .I(N__21345));
    InMux I__2523 (
            .O(N__21351),
            .I(N__21342));
    LocalMux I__2522 (
            .O(N__21348),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    LocalMux I__2521 (
            .O(N__21345),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    LocalMux I__2520 (
            .O(N__21342),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    InMux I__2519 (
            .O(N__21335),
            .I(bfn_8_20_0_));
    CascadeMux I__2518 (
            .O(N__21332),
            .I(N__21328));
    InMux I__2517 (
            .O(N__21331),
            .I(N__21324));
    InMux I__2516 (
            .O(N__21328),
            .I(N__21321));
    InMux I__2515 (
            .O(N__21327),
            .I(N__21318));
    LocalMux I__2514 (
            .O(N__21324),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    LocalMux I__2513 (
            .O(N__21321),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    LocalMux I__2512 (
            .O(N__21318),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    InMux I__2511 (
            .O(N__21311),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    CascadeMux I__2510 (
            .O(N__21308),
            .I(N__21304));
    InMux I__2509 (
            .O(N__21307),
            .I(N__21300));
    InMux I__2508 (
            .O(N__21304),
            .I(N__21297));
    InMux I__2507 (
            .O(N__21303),
            .I(N__21294));
    LocalMux I__2506 (
            .O(N__21300),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    LocalMux I__2505 (
            .O(N__21297),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    LocalMux I__2504 (
            .O(N__21294),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    InMux I__2503 (
            .O(N__21287),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    CascadeMux I__2502 (
            .O(N__21284),
            .I(N__21280));
    InMux I__2501 (
            .O(N__21283),
            .I(N__21276));
    InMux I__2500 (
            .O(N__21280),
            .I(N__21273));
    InMux I__2499 (
            .O(N__21279),
            .I(N__21270));
    LocalMux I__2498 (
            .O(N__21276),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    LocalMux I__2497 (
            .O(N__21273),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    LocalMux I__2496 (
            .O(N__21270),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__2495 (
            .O(N__21263),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    InMux I__2494 (
            .O(N__21260),
            .I(N__21257));
    LocalMux I__2493 (
            .O(N__21257),
            .I(N__21252));
    InMux I__2492 (
            .O(N__21256),
            .I(N__21249));
    InMux I__2491 (
            .O(N__21255),
            .I(N__21246));
    Odrv4 I__2490 (
            .O(N__21252),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    LocalMux I__2489 (
            .O(N__21249),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    LocalMux I__2488 (
            .O(N__21246),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    InMux I__2487 (
            .O(N__21239),
            .I(bfn_8_19_0_));
    InMux I__2486 (
            .O(N__21236),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    CascadeMux I__2485 (
            .O(N__21233),
            .I(N__21228));
    CascadeMux I__2484 (
            .O(N__21232),
            .I(N__21225));
    InMux I__2483 (
            .O(N__21231),
            .I(N__21222));
    InMux I__2482 (
            .O(N__21228),
            .I(N__21217));
    InMux I__2481 (
            .O(N__21225),
            .I(N__21217));
    LocalMux I__2480 (
            .O(N__21222),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    LocalMux I__2479 (
            .O(N__21217),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    InMux I__2478 (
            .O(N__21212),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    CascadeMux I__2477 (
            .O(N__21209),
            .I(N__21204));
    CascadeMux I__2476 (
            .O(N__21208),
            .I(N__21201));
    InMux I__2475 (
            .O(N__21207),
            .I(N__21198));
    InMux I__2474 (
            .O(N__21204),
            .I(N__21193));
    InMux I__2473 (
            .O(N__21201),
            .I(N__21193));
    LocalMux I__2472 (
            .O(N__21198),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    LocalMux I__2471 (
            .O(N__21193),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    InMux I__2470 (
            .O(N__21188),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    InMux I__2469 (
            .O(N__21185),
            .I(N__21182));
    LocalMux I__2468 (
            .O(N__21182),
            .I(\current_shift_inst.elapsed_time_ns_s1_fast_31 ));
    CascadeMux I__2467 (
            .O(N__21179),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ));
    CascadeMux I__2466 (
            .O(N__21176),
            .I(N__21173));
    InMux I__2465 (
            .O(N__21173),
            .I(N__21169));
    InMux I__2464 (
            .O(N__21172),
            .I(N__21166));
    LocalMux I__2463 (
            .O(N__21169),
            .I(N__21160));
    LocalMux I__2462 (
            .O(N__21166),
            .I(N__21160));
    InMux I__2461 (
            .O(N__21165),
            .I(N__21157));
    Span4Mux_v I__2460 (
            .O(N__21160),
            .I(N__21154));
    LocalMux I__2459 (
            .O(N__21157),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__2458 (
            .O(N__21154),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__2457 (
            .O(N__21149),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__2456 (
            .O(N__21146),
            .I(N__21142));
    InMux I__2455 (
            .O(N__21145),
            .I(N__21139));
    LocalMux I__2454 (
            .O(N__21142),
            .I(N__21136));
    LocalMux I__2453 (
            .O(N__21139),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    Odrv12 I__2452 (
            .O(N__21136),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    CascadeMux I__2451 (
            .O(N__21131),
            .I(N__21128));
    InMux I__2450 (
            .O(N__21128),
            .I(N__21123));
    InMux I__2449 (
            .O(N__21127),
            .I(N__21120));
    InMux I__2448 (
            .O(N__21126),
            .I(N__21117));
    LocalMux I__2447 (
            .O(N__21123),
            .I(N__21112));
    LocalMux I__2446 (
            .O(N__21120),
            .I(N__21112));
    LocalMux I__2445 (
            .O(N__21117),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    Odrv12 I__2444 (
            .O(N__21112),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    InMux I__2443 (
            .O(N__21107),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__2442 (
            .O(N__21104),
            .I(N__21100));
    InMux I__2441 (
            .O(N__21103),
            .I(N__21097));
    LocalMux I__2440 (
            .O(N__21100),
            .I(N__21094));
    LocalMux I__2439 (
            .O(N__21097),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    Odrv12 I__2438 (
            .O(N__21094),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    CascadeMux I__2437 (
            .O(N__21089),
            .I(N__21086));
    InMux I__2436 (
            .O(N__21086),
            .I(N__21081));
    InMux I__2435 (
            .O(N__21085),
            .I(N__21078));
    InMux I__2434 (
            .O(N__21084),
            .I(N__21075));
    LocalMux I__2433 (
            .O(N__21081),
            .I(N__21070));
    LocalMux I__2432 (
            .O(N__21078),
            .I(N__21070));
    LocalMux I__2431 (
            .O(N__21075),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    Odrv12 I__2430 (
            .O(N__21070),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__2429 (
            .O(N__21065),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__2428 (
            .O(N__21062),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__2427 (
            .O(N__21059),
            .I(N__21056));
    LocalMux I__2426 (
            .O(N__21056),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ));
    CascadeMux I__2425 (
            .O(N__21053),
            .I(N__21050));
    InMux I__2424 (
            .O(N__21050),
            .I(N__21046));
    InMux I__2423 (
            .O(N__21049),
            .I(N__21043));
    LocalMux I__2422 (
            .O(N__21046),
            .I(N__21037));
    LocalMux I__2421 (
            .O(N__21043),
            .I(N__21037));
    InMux I__2420 (
            .O(N__21042),
            .I(N__21034));
    Span4Mux_v I__2419 (
            .O(N__21037),
            .I(N__21031));
    LocalMux I__2418 (
            .O(N__21034),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__2417 (
            .O(N__21031),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__2416 (
            .O(N__21026),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__2415 (
            .O(N__21023),
            .I(N__21020));
    InMux I__2414 (
            .O(N__21020),
            .I(N__21015));
    InMux I__2413 (
            .O(N__21019),
            .I(N__21012));
    InMux I__2412 (
            .O(N__21018),
            .I(N__21009));
    LocalMux I__2411 (
            .O(N__21015),
            .I(N__21004));
    LocalMux I__2410 (
            .O(N__21012),
            .I(N__21004));
    LocalMux I__2409 (
            .O(N__21009),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    Odrv12 I__2408 (
            .O(N__21004),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__2407 (
            .O(N__20999),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__2406 (
            .O(N__20996),
            .I(N__20989));
    InMux I__2405 (
            .O(N__20995),
            .I(N__20989));
    InMux I__2404 (
            .O(N__20994),
            .I(N__20986));
    LocalMux I__2403 (
            .O(N__20989),
            .I(N__20983));
    LocalMux I__2402 (
            .O(N__20986),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    Odrv12 I__2401 (
            .O(N__20983),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__2400 (
            .O(N__20978),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__2399 (
            .O(N__20975),
            .I(N__20968));
    InMux I__2398 (
            .O(N__20974),
            .I(N__20968));
    InMux I__2397 (
            .O(N__20973),
            .I(N__20965));
    LocalMux I__2396 (
            .O(N__20968),
            .I(N__20962));
    LocalMux I__2395 (
            .O(N__20965),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    Odrv12 I__2394 (
            .O(N__20962),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__2393 (
            .O(N__20957),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__2392 (
            .O(N__20954),
            .I(N__20950));
    InMux I__2391 (
            .O(N__20953),
            .I(N__20946));
    InMux I__2390 (
            .O(N__20950),
            .I(N__20943));
    InMux I__2389 (
            .O(N__20949),
            .I(N__20940));
    LocalMux I__2388 (
            .O(N__20946),
            .I(N__20935));
    LocalMux I__2387 (
            .O(N__20943),
            .I(N__20935));
    LocalMux I__2386 (
            .O(N__20940),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    Odrv12 I__2385 (
            .O(N__20935),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__2384 (
            .O(N__20930),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__2383 (
            .O(N__20927),
            .I(N__20923));
    CascadeMux I__2382 (
            .O(N__20926),
            .I(N__20920));
    InMux I__2381 (
            .O(N__20923),
            .I(N__20915));
    InMux I__2380 (
            .O(N__20920),
            .I(N__20915));
    LocalMux I__2379 (
            .O(N__20915),
            .I(N__20911));
    InMux I__2378 (
            .O(N__20914),
            .I(N__20908));
    Span4Mux_v I__2377 (
            .O(N__20911),
            .I(N__20905));
    LocalMux I__2376 (
            .O(N__20908),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    Odrv4 I__2375 (
            .O(N__20905),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__2374 (
            .O(N__20900),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__2373 (
            .O(N__20897),
            .I(N__20893));
    CascadeMux I__2372 (
            .O(N__20896),
            .I(N__20890));
    InMux I__2371 (
            .O(N__20893),
            .I(N__20884));
    InMux I__2370 (
            .O(N__20890),
            .I(N__20884));
    InMux I__2369 (
            .O(N__20889),
            .I(N__20881));
    LocalMux I__2368 (
            .O(N__20884),
            .I(N__20878));
    LocalMux I__2367 (
            .O(N__20881),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    Odrv12 I__2366 (
            .O(N__20878),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__2365 (
            .O(N__20873),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__2364 (
            .O(N__20870),
            .I(N__20867));
    InMux I__2363 (
            .O(N__20867),
            .I(N__20863));
    InMux I__2362 (
            .O(N__20866),
            .I(N__20860));
    LocalMux I__2361 (
            .O(N__20863),
            .I(N__20854));
    LocalMux I__2360 (
            .O(N__20860),
            .I(N__20854));
    InMux I__2359 (
            .O(N__20859),
            .I(N__20851));
    Span4Mux_v I__2358 (
            .O(N__20854),
            .I(N__20848));
    LocalMux I__2357 (
            .O(N__20851),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv4 I__2356 (
            .O(N__20848),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__2355 (
            .O(N__20843),
            .I(bfn_8_14_0_));
    CascadeMux I__2354 (
            .O(N__20840),
            .I(N__20837));
    InMux I__2353 (
            .O(N__20837),
            .I(N__20833));
    CascadeMux I__2352 (
            .O(N__20836),
            .I(N__20830));
    LocalMux I__2351 (
            .O(N__20833),
            .I(N__20826));
    InMux I__2350 (
            .O(N__20830),
            .I(N__20823));
    InMux I__2349 (
            .O(N__20829),
            .I(N__20820));
    Sp12to4 I__2348 (
            .O(N__20826),
            .I(N__20815));
    LocalMux I__2347 (
            .O(N__20823),
            .I(N__20815));
    LocalMux I__2346 (
            .O(N__20820),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv12 I__2345 (
            .O(N__20815),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__2344 (
            .O(N__20810),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__2343 (
            .O(N__20807),
            .I(N__20801));
    InMux I__2342 (
            .O(N__20806),
            .I(N__20801));
    LocalMux I__2341 (
            .O(N__20801),
            .I(N__20797));
    InMux I__2340 (
            .O(N__20800),
            .I(N__20794));
    Span4Mux_v I__2339 (
            .O(N__20797),
            .I(N__20791));
    LocalMux I__2338 (
            .O(N__20794),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    Odrv4 I__2337 (
            .O(N__20791),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__2336 (
            .O(N__20786),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__2335 (
            .O(N__20783),
            .I(N__20776));
    InMux I__2334 (
            .O(N__20782),
            .I(N__20776));
    InMux I__2333 (
            .O(N__20781),
            .I(N__20773));
    LocalMux I__2332 (
            .O(N__20776),
            .I(N__20770));
    LocalMux I__2331 (
            .O(N__20773),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    Odrv12 I__2330 (
            .O(N__20770),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__2329 (
            .O(N__20765),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__2328 (
            .O(N__20762),
            .I(N__20758));
    CascadeMux I__2327 (
            .O(N__20761),
            .I(N__20755));
    InMux I__2326 (
            .O(N__20758),
            .I(N__20749));
    InMux I__2325 (
            .O(N__20755),
            .I(N__20749));
    InMux I__2324 (
            .O(N__20754),
            .I(N__20746));
    LocalMux I__2323 (
            .O(N__20749),
            .I(N__20743));
    LocalMux I__2322 (
            .O(N__20746),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    Odrv12 I__2321 (
            .O(N__20743),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__2320 (
            .O(N__20738),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__2319 (
            .O(N__20735),
            .I(N__20731));
    CascadeMux I__2318 (
            .O(N__20734),
            .I(N__20728));
    InMux I__2317 (
            .O(N__20731),
            .I(N__20722));
    InMux I__2316 (
            .O(N__20728),
            .I(N__20722));
    InMux I__2315 (
            .O(N__20727),
            .I(N__20719));
    LocalMux I__2314 (
            .O(N__20722),
            .I(N__20716));
    LocalMux I__2313 (
            .O(N__20719),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    Odrv12 I__2312 (
            .O(N__20716),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__2311 (
            .O(N__20711),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__2310 (
            .O(N__20708),
            .I(N__20705));
    InMux I__2309 (
            .O(N__20705),
            .I(N__20701));
    InMux I__2308 (
            .O(N__20704),
            .I(N__20698));
    LocalMux I__2307 (
            .O(N__20701),
            .I(N__20692));
    LocalMux I__2306 (
            .O(N__20698),
            .I(N__20692));
    InMux I__2305 (
            .O(N__20697),
            .I(N__20689));
    Span4Mux_v I__2304 (
            .O(N__20692),
            .I(N__20686));
    LocalMux I__2303 (
            .O(N__20689),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    Odrv4 I__2302 (
            .O(N__20686),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__2301 (
            .O(N__20681),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__2300 (
            .O(N__20678),
            .I(N__20675));
    InMux I__2299 (
            .O(N__20675),
            .I(N__20671));
    InMux I__2298 (
            .O(N__20674),
            .I(N__20668));
    LocalMux I__2297 (
            .O(N__20671),
            .I(N__20662));
    LocalMux I__2296 (
            .O(N__20668),
            .I(N__20662));
    InMux I__2295 (
            .O(N__20667),
            .I(N__20659));
    Span4Mux_v I__2294 (
            .O(N__20662),
            .I(N__20656));
    LocalMux I__2293 (
            .O(N__20659),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    Odrv4 I__2292 (
            .O(N__20656),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__2291 (
            .O(N__20651),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__2290 (
            .O(N__20648),
            .I(N__20645));
    InMux I__2289 (
            .O(N__20645),
            .I(N__20640));
    InMux I__2288 (
            .O(N__20644),
            .I(N__20637));
    InMux I__2287 (
            .O(N__20643),
            .I(N__20634));
    LocalMux I__2286 (
            .O(N__20640),
            .I(N__20629));
    LocalMux I__2285 (
            .O(N__20637),
            .I(N__20629));
    LocalMux I__2284 (
            .O(N__20634),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv12 I__2283 (
            .O(N__20629),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__2282 (
            .O(N__20624),
            .I(bfn_8_13_0_));
    InMux I__2281 (
            .O(N__20621),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__2280 (
            .O(N__20618),
            .I(N__20614));
    InMux I__2279 (
            .O(N__20617),
            .I(N__20611));
    InMux I__2278 (
            .O(N__20614),
            .I(N__20608));
    LocalMux I__2277 (
            .O(N__20611),
            .I(N__20602));
    LocalMux I__2276 (
            .O(N__20608),
            .I(N__20602));
    InMux I__2275 (
            .O(N__20607),
            .I(N__20599));
    Span4Mux_v I__2274 (
            .O(N__20602),
            .I(N__20596));
    LocalMux I__2273 (
            .O(N__20599),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    Odrv4 I__2272 (
            .O(N__20596),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__2271 (
            .O(N__20591),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__2270 (
            .O(N__20588),
            .I(N__20582));
    InMux I__2269 (
            .O(N__20587),
            .I(N__20582));
    LocalMux I__2268 (
            .O(N__20582),
            .I(N__20578));
    InMux I__2267 (
            .O(N__20581),
            .I(N__20575));
    Span4Mux_v I__2266 (
            .O(N__20578),
            .I(N__20572));
    LocalMux I__2265 (
            .O(N__20575),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    Odrv4 I__2264 (
            .O(N__20572),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__2263 (
            .O(N__20567),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__2262 (
            .O(N__20564),
            .I(N__20560));
    CascadeMux I__2261 (
            .O(N__20563),
            .I(N__20557));
    InMux I__2260 (
            .O(N__20560),
            .I(N__20551));
    InMux I__2259 (
            .O(N__20557),
            .I(N__20551));
    InMux I__2258 (
            .O(N__20556),
            .I(N__20548));
    LocalMux I__2257 (
            .O(N__20551),
            .I(N__20545));
    LocalMux I__2256 (
            .O(N__20548),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    Odrv12 I__2255 (
            .O(N__20545),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__2254 (
            .O(N__20540),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__2253 (
            .O(N__20537),
            .I(N__20533));
    CascadeMux I__2252 (
            .O(N__20536),
            .I(N__20530));
    InMux I__2251 (
            .O(N__20533),
            .I(N__20524));
    InMux I__2250 (
            .O(N__20530),
            .I(N__20524));
    InMux I__2249 (
            .O(N__20529),
            .I(N__20521));
    LocalMux I__2248 (
            .O(N__20524),
            .I(N__20518));
    LocalMux I__2247 (
            .O(N__20521),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    Odrv12 I__2246 (
            .O(N__20518),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__2245 (
            .O(N__20513),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__2244 (
            .O(N__20510),
            .I(N__20504));
    InMux I__2243 (
            .O(N__20509),
            .I(N__20504));
    LocalMux I__2242 (
            .O(N__20504),
            .I(N__20500));
    InMux I__2241 (
            .O(N__20503),
            .I(N__20497));
    Span4Mux_v I__2240 (
            .O(N__20500),
            .I(N__20494));
    LocalMux I__2239 (
            .O(N__20497),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    Odrv4 I__2238 (
            .O(N__20494),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__2237 (
            .O(N__20489),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__2236 (
            .O(N__20486),
            .I(N__20480));
    InMux I__2235 (
            .O(N__20485),
            .I(N__20480));
    LocalMux I__2234 (
            .O(N__20480),
            .I(N__20476));
    InMux I__2233 (
            .O(N__20479),
            .I(N__20473));
    Span4Mux_v I__2232 (
            .O(N__20476),
            .I(N__20470));
    LocalMux I__2231 (
            .O(N__20473),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    Odrv4 I__2230 (
            .O(N__20470),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__2229 (
            .O(N__20465),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__2228 (
            .O(N__20462),
            .I(N__20458));
    CascadeMux I__2227 (
            .O(N__20461),
            .I(N__20455));
    InMux I__2226 (
            .O(N__20458),
            .I(N__20452));
    InMux I__2225 (
            .O(N__20455),
            .I(N__20449));
    LocalMux I__2224 (
            .O(N__20452),
            .I(N__20443));
    LocalMux I__2223 (
            .O(N__20449),
            .I(N__20443));
    InMux I__2222 (
            .O(N__20448),
            .I(N__20440));
    Span4Mux_v I__2221 (
            .O(N__20443),
            .I(N__20437));
    LocalMux I__2220 (
            .O(N__20440),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv4 I__2219 (
            .O(N__20437),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__2218 (
            .O(N__20432),
            .I(N__20427));
    InMux I__2217 (
            .O(N__20431),
            .I(N__20424));
    InMux I__2216 (
            .O(N__20430),
            .I(N__20421));
    LocalMux I__2215 (
            .O(N__20427),
            .I(N__20418));
    LocalMux I__2214 (
            .O(N__20424),
            .I(N__20415));
    LocalMux I__2213 (
            .O(N__20421),
            .I(N__20411));
    Span4Mux_v I__2212 (
            .O(N__20418),
            .I(N__20406));
    Span4Mux_h I__2211 (
            .O(N__20415),
            .I(N__20406));
    InMux I__2210 (
            .O(N__20414),
            .I(N__20403));
    Odrv12 I__2209 (
            .O(N__20411),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    Odrv4 I__2208 (
            .O(N__20406),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    LocalMux I__2207 (
            .O(N__20403),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    InMux I__2206 (
            .O(N__20396),
            .I(bfn_8_12_0_));
    InMux I__2205 (
            .O(N__20393),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    InMux I__2204 (
            .O(N__20390),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    InMux I__2203 (
            .O(N__20387),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    InMux I__2202 (
            .O(N__20384),
            .I(bfn_8_10_0_));
    InMux I__2201 (
            .O(N__20381),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    InMux I__2200 (
            .O(N__20378),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    InMux I__2199 (
            .O(N__20375),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    InMux I__2198 (
            .O(N__20372),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__2197 (
            .O(N__20369),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    InMux I__2196 (
            .O(N__20366),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    InMux I__2195 (
            .O(N__20363),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    InMux I__2194 (
            .O(N__20360),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    InMux I__2193 (
            .O(N__20357),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    InMux I__2192 (
            .O(N__20354),
            .I(bfn_8_9_0_));
    InMux I__2191 (
            .O(N__20351),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    InMux I__2190 (
            .O(N__20348),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    InMux I__2189 (
            .O(N__20345),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    InMux I__2188 (
            .O(N__20342),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    InMux I__2187 (
            .O(N__20339),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    InMux I__2186 (
            .O(N__20336),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    InMux I__2185 (
            .O(N__20333),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    InMux I__2184 (
            .O(N__20330),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    InMux I__2183 (
            .O(N__20327),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    InMux I__2182 (
            .O(N__20324),
            .I(bfn_8_8_0_));
    InMux I__2181 (
            .O(N__20321),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    InMux I__2180 (
            .O(N__20318),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    InMux I__2179 (
            .O(N__20315),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    InMux I__2178 (
            .O(N__20312),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    InMux I__2177 (
            .O(N__20309),
            .I(N__20305));
    InMux I__2176 (
            .O(N__20308),
            .I(N__20302));
    LocalMux I__2175 (
            .O(N__20305),
            .I(N__20299));
    LocalMux I__2174 (
            .O(N__20302),
            .I(N__20296));
    Span4Mux_v I__2173 (
            .O(N__20299),
            .I(N__20293));
    Span12Mux_v I__2172 (
            .O(N__20296),
            .I(N__20290));
    Span4Mux_h I__2171 (
            .O(N__20293),
            .I(N__20287));
    Odrv12 I__2170 (
            .O(N__20290),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv4 I__2169 (
            .O(N__20287),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    InMux I__2168 (
            .O(N__20282),
            .I(N__20279));
    LocalMux I__2167 (
            .O(N__20279),
            .I(N__20276));
    Odrv12 I__2166 (
            .O(N__20276),
            .I(il_max_comp1_c));
    InMux I__2165 (
            .O(N__20273),
            .I(bfn_8_7_0_));
    InMux I__2164 (
            .O(N__20270),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    InMux I__2163 (
            .O(N__20267),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    InMux I__2162 (
            .O(N__20264),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    InMux I__2161 (
            .O(N__20261),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    InMux I__2160 (
            .O(N__20258),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    InMux I__2159 (
            .O(N__20255),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    InMux I__2158 (
            .O(N__20252),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    InMux I__2157 (
            .O(N__20249),
            .I(bfn_7_23_0_));
    InMux I__2156 (
            .O(N__20246),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    InMux I__2155 (
            .O(N__20243),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    InMux I__2154 (
            .O(N__20240),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    InMux I__2153 (
            .O(N__20237),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    InMux I__2152 (
            .O(N__20234),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    InMux I__2151 (
            .O(N__20231),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    InMux I__2150 (
            .O(N__20228),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    InMux I__2149 (
            .O(N__20225),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    InMux I__2148 (
            .O(N__20222),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    InMux I__2147 (
            .O(N__20219),
            .I(bfn_7_22_0_));
    InMux I__2146 (
            .O(N__20216),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    InMux I__2145 (
            .O(N__20213),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    InMux I__2144 (
            .O(N__20210),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    InMux I__2143 (
            .O(N__20207),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    InMux I__2142 (
            .O(N__20204),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    InMux I__2141 (
            .O(N__20201),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    InMux I__2140 (
            .O(N__20198),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    InMux I__2139 (
            .O(N__20195),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    InMux I__2138 (
            .O(N__20192),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    InMux I__2137 (
            .O(N__20189),
            .I(bfn_7_21_0_));
    InMux I__2136 (
            .O(N__20186),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    InMux I__2135 (
            .O(N__20183),
            .I(bfn_7_14_0_));
    InMux I__2134 (
            .O(N__20180),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ));
    InMux I__2133 (
            .O(N__20177),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ));
    InMux I__2132 (
            .O(N__20174),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ));
    InMux I__2131 (
            .O(N__20171),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ));
    InMux I__2130 (
            .O(N__20168),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ));
    InMux I__2129 (
            .O(N__20165),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ));
    InMux I__2128 (
            .O(N__20162),
            .I(N__20159));
    LocalMux I__2127 (
            .O(N__20159),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ));
    InMux I__2126 (
            .O(N__20156),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ));
    InMux I__2125 (
            .O(N__20153),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ));
    InMux I__2124 (
            .O(N__20150),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ));
    InMux I__2123 (
            .O(N__20147),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ));
    InMux I__2122 (
            .O(N__20144),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ));
    InMux I__2121 (
            .O(N__20141),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ));
    InMux I__2120 (
            .O(N__20138),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ));
    CascadeMux I__2119 (
            .O(N__20135),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3_cascade_ ));
    InMux I__2118 (
            .O(N__20132),
            .I(N__20129));
    LocalMux I__2117 (
            .O(N__20129),
            .I(N__20126));
    Odrv4 I__2116 (
            .O(N__20126),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17 ));
    CascadeMux I__2115 (
            .O(N__20123),
            .I(N__20119));
    InMux I__2114 (
            .O(N__20122),
            .I(N__20114));
    InMux I__2113 (
            .O(N__20119),
            .I(N__20114));
    LocalMux I__2112 (
            .O(N__20114),
            .I(N__20111));
    Odrv4 I__2111 (
            .O(N__20111),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ));
    InMux I__2110 (
            .O(N__20108),
            .I(N__20102));
    InMux I__2109 (
            .O(N__20107),
            .I(N__20102));
    LocalMux I__2108 (
            .O(N__20102),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ));
    InMux I__2107 (
            .O(N__20099),
            .I(N__20096));
    LocalMux I__2106 (
            .O(N__20096),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ));
    InMux I__2105 (
            .O(N__20093),
            .I(N__20090));
    LocalMux I__2104 (
            .O(N__20090),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ));
    InMux I__2103 (
            .O(N__20087),
            .I(N__20084));
    LocalMux I__2102 (
            .O(N__20084),
            .I(N__20081));
    Glb2LocalMux I__2101 (
            .O(N__20081),
            .I(N__20078));
    GlobalMux I__2100 (
            .O(N__20078),
            .I(clk_12mhz));
    IoInMux I__2099 (
            .O(N__20075),
            .I(N__20072));
    LocalMux I__2098 (
            .O(N__20072),
            .I(N__20069));
    IoSpan4Mux I__2097 (
            .O(N__20069),
            .I(N__20066));
    Span4Mux_s0_v I__2096 (
            .O(N__20066),
            .I(N__20063));
    Odrv4 I__2095 (
            .O(N__20063),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__2094 (
            .O(N__20060),
            .I(N__20057));
    LocalMux I__2093 (
            .O(N__20057),
            .I(N__20052));
    InMux I__2092 (
            .O(N__20056),
            .I(N__20049));
    InMux I__2091 (
            .O(N__20055),
            .I(N__20046));
    Span4Mux_h I__2090 (
            .O(N__20052),
            .I(N__20043));
    LocalMux I__2089 (
            .O(N__20049),
            .I(N__20040));
    LocalMux I__2088 (
            .O(N__20046),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    Odrv4 I__2087 (
            .O(N__20043),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    Odrv4 I__2086 (
            .O(N__20040),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    CascadeMux I__2085 (
            .O(N__20033),
            .I(N__20030));
    InMux I__2084 (
            .O(N__20030),
            .I(N__20027));
    LocalMux I__2083 (
            .O(N__20027),
            .I(N__20024));
    Odrv4 I__2082 (
            .O(N__20024),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    CascadeMux I__2081 (
            .O(N__20021),
            .I(N__20018));
    InMux I__2080 (
            .O(N__20018),
            .I(N__20015));
    LocalMux I__2079 (
            .O(N__20015),
            .I(N__20012));
    Odrv4 I__2078 (
            .O(N__20012),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    InMux I__2077 (
            .O(N__20009),
            .I(N__20005));
    InMux I__2076 (
            .O(N__20008),
            .I(N__20002));
    LocalMux I__2075 (
            .O(N__20005),
            .I(N__19992));
    LocalMux I__2074 (
            .O(N__20002),
            .I(N__19992));
    InMux I__2073 (
            .O(N__20001),
            .I(N__19987));
    InMux I__2072 (
            .O(N__20000),
            .I(N__19987));
    InMux I__2071 (
            .O(N__19999),
            .I(N__19984));
    InMux I__2070 (
            .O(N__19998),
            .I(N__19973));
    InMux I__2069 (
            .O(N__19997),
            .I(N__19970));
    Span4Mux_v I__2068 (
            .O(N__19992),
            .I(N__19953));
    LocalMux I__2067 (
            .O(N__19987),
            .I(N__19953));
    LocalMux I__2066 (
            .O(N__19984),
            .I(N__19950));
    InMux I__2065 (
            .O(N__19983),
            .I(N__19947));
    InMux I__2064 (
            .O(N__19982),
            .I(N__19940));
    InMux I__2063 (
            .O(N__19981),
            .I(N__19940));
    InMux I__2062 (
            .O(N__19980),
            .I(N__19940));
    InMux I__2061 (
            .O(N__19979),
            .I(N__19931));
    InMux I__2060 (
            .O(N__19978),
            .I(N__19931));
    InMux I__2059 (
            .O(N__19977),
            .I(N__19931));
    InMux I__2058 (
            .O(N__19976),
            .I(N__19931));
    LocalMux I__2057 (
            .O(N__19973),
            .I(N__19928));
    LocalMux I__2056 (
            .O(N__19970),
            .I(N__19922));
    InMux I__2055 (
            .O(N__19969),
            .I(N__19907));
    InMux I__2054 (
            .O(N__19968),
            .I(N__19907));
    InMux I__2053 (
            .O(N__19967),
            .I(N__19907));
    InMux I__2052 (
            .O(N__19966),
            .I(N__19907));
    InMux I__2051 (
            .O(N__19965),
            .I(N__19907));
    InMux I__2050 (
            .O(N__19964),
            .I(N__19907));
    InMux I__2049 (
            .O(N__19963),
            .I(N__19907));
    InMux I__2048 (
            .O(N__19962),
            .I(N__19896));
    InMux I__2047 (
            .O(N__19961),
            .I(N__19896));
    InMux I__2046 (
            .O(N__19960),
            .I(N__19896));
    InMux I__2045 (
            .O(N__19959),
            .I(N__19896));
    InMux I__2044 (
            .O(N__19958),
            .I(N__19896));
    Span4Mux_v I__2043 (
            .O(N__19953),
            .I(N__19892));
    Span4Mux_v I__2042 (
            .O(N__19950),
            .I(N__19887));
    LocalMux I__2041 (
            .O(N__19947),
            .I(N__19887));
    LocalMux I__2040 (
            .O(N__19940),
            .I(N__19882));
    LocalMux I__2039 (
            .O(N__19931),
            .I(N__19882));
    Span4Mux_h I__2038 (
            .O(N__19928),
            .I(N__19879));
    InMux I__2037 (
            .O(N__19927),
            .I(N__19872));
    InMux I__2036 (
            .O(N__19926),
            .I(N__19872));
    InMux I__2035 (
            .O(N__19925),
            .I(N__19872));
    Span4Mux_h I__2034 (
            .O(N__19922),
            .I(N__19865));
    LocalMux I__2033 (
            .O(N__19907),
            .I(N__19865));
    LocalMux I__2032 (
            .O(N__19896),
            .I(N__19865));
    InMux I__2031 (
            .O(N__19895),
            .I(N__19862));
    Odrv4 I__2030 (
            .O(N__19892),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv4 I__2029 (
            .O(N__19887),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv12 I__2028 (
            .O(N__19882),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv4 I__2027 (
            .O(N__19879),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    LocalMux I__2026 (
            .O(N__19872),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv4 I__2025 (
            .O(N__19865),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    LocalMux I__2024 (
            .O(N__19862),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    CascadeMux I__2023 (
            .O(N__19847),
            .I(N__19844));
    InMux I__2022 (
            .O(N__19844),
            .I(N__19841));
    LocalMux I__2021 (
            .O(N__19841),
            .I(N__19838));
    Span4Mux_h I__2020 (
            .O(N__19838),
            .I(N__19835));
    Odrv4 I__2019 (
            .O(N__19835),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    CascadeMux I__2018 (
            .O(N__19832),
            .I(N__19825));
    InMux I__2017 (
            .O(N__19831),
            .I(N__19811));
    InMux I__2016 (
            .O(N__19830),
            .I(N__19808));
    CascadeMux I__2015 (
            .O(N__19829),
            .I(N__19799));
    InMux I__2014 (
            .O(N__19828),
            .I(N__19796));
    InMux I__2013 (
            .O(N__19825),
            .I(N__19789));
    InMux I__2012 (
            .O(N__19824),
            .I(N__19789));
    InMux I__2011 (
            .O(N__19823),
            .I(N__19789));
    CascadeMux I__2010 (
            .O(N__19822),
            .I(N__19785));
    CascadeMux I__2009 (
            .O(N__19821),
            .I(N__19782));
    CascadeMux I__2008 (
            .O(N__19820),
            .I(N__19779));
    CascadeMux I__2007 (
            .O(N__19819),
            .I(N__19773));
    CascadeMux I__2006 (
            .O(N__19818),
            .I(N__19770));
    CascadeMux I__2005 (
            .O(N__19817),
            .I(N__19767));
    CascadeMux I__2004 (
            .O(N__19816),
            .I(N__19764));
    InMux I__2003 (
            .O(N__19815),
            .I(N__19761));
    InMux I__2002 (
            .O(N__19814),
            .I(N__19758));
    LocalMux I__2001 (
            .O(N__19811),
            .I(N__19755));
    LocalMux I__2000 (
            .O(N__19808),
            .I(N__19752));
    CascadeMux I__1999 (
            .O(N__19807),
            .I(N__19749));
    CascadeMux I__1998 (
            .O(N__19806),
            .I(N__19744));
    InMux I__1997 (
            .O(N__19805),
            .I(N__19741));
    CascadeMux I__1996 (
            .O(N__19804),
            .I(N__19735));
    CascadeMux I__1995 (
            .O(N__19803),
            .I(N__19732));
    InMux I__1994 (
            .O(N__19802),
            .I(N__19729));
    InMux I__1993 (
            .O(N__19799),
            .I(N__19726));
    LocalMux I__1992 (
            .O(N__19796),
            .I(N__19721));
    LocalMux I__1991 (
            .O(N__19789),
            .I(N__19721));
    InMux I__1990 (
            .O(N__19788),
            .I(N__19712));
    InMux I__1989 (
            .O(N__19785),
            .I(N__19712));
    InMux I__1988 (
            .O(N__19782),
            .I(N__19712));
    InMux I__1987 (
            .O(N__19779),
            .I(N__19712));
    InMux I__1986 (
            .O(N__19778),
            .I(N__19697));
    InMux I__1985 (
            .O(N__19777),
            .I(N__19697));
    InMux I__1984 (
            .O(N__19776),
            .I(N__19697));
    InMux I__1983 (
            .O(N__19773),
            .I(N__19697));
    InMux I__1982 (
            .O(N__19770),
            .I(N__19697));
    InMux I__1981 (
            .O(N__19767),
            .I(N__19697));
    InMux I__1980 (
            .O(N__19764),
            .I(N__19697));
    LocalMux I__1979 (
            .O(N__19761),
            .I(N__19694));
    LocalMux I__1978 (
            .O(N__19758),
            .I(N__19687));
    Span4Mux_h I__1977 (
            .O(N__19755),
            .I(N__19687));
    Span4Mux_s3_h I__1976 (
            .O(N__19752),
            .I(N__19687));
    InMux I__1975 (
            .O(N__19749),
            .I(N__19684));
    InMux I__1974 (
            .O(N__19748),
            .I(N__19677));
    InMux I__1973 (
            .O(N__19747),
            .I(N__19677));
    InMux I__1972 (
            .O(N__19744),
            .I(N__19677));
    LocalMux I__1971 (
            .O(N__19741),
            .I(N__19674));
    InMux I__1970 (
            .O(N__19740),
            .I(N__19663));
    InMux I__1969 (
            .O(N__19739),
            .I(N__19663));
    InMux I__1968 (
            .O(N__19738),
            .I(N__19663));
    InMux I__1967 (
            .O(N__19735),
            .I(N__19663));
    InMux I__1966 (
            .O(N__19732),
            .I(N__19663));
    LocalMux I__1965 (
            .O(N__19729),
            .I(N__19658));
    LocalMux I__1964 (
            .O(N__19726),
            .I(N__19658));
    Span4Mux_h I__1963 (
            .O(N__19721),
            .I(N__19649));
    LocalMux I__1962 (
            .O(N__19712),
            .I(N__19649));
    LocalMux I__1961 (
            .O(N__19697),
            .I(N__19649));
    Span4Mux_h I__1960 (
            .O(N__19694),
            .I(N__19649));
    Span4Mux_v I__1959 (
            .O(N__19687),
            .I(N__19646));
    LocalMux I__1958 (
            .O(N__19684),
            .I(N__19635));
    LocalMux I__1957 (
            .O(N__19677),
            .I(N__19635));
    Span4Mux_h I__1956 (
            .O(N__19674),
            .I(N__19635));
    LocalMux I__1955 (
            .O(N__19663),
            .I(N__19635));
    Span4Mux_h I__1954 (
            .O(N__19658),
            .I(N__19635));
    Span4Mux_v I__1953 (
            .O(N__19649),
            .I(N__19632));
    Span4Mux_v I__1952 (
            .O(N__19646),
            .I(N__19629));
    Span4Mux_v I__1951 (
            .O(N__19635),
            .I(N__19626));
    Span4Mux_v I__1950 (
            .O(N__19632),
            .I(N__19623));
    Odrv4 I__1949 (
            .O(N__19629),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv4 I__1948 (
            .O(N__19626),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv4 I__1947 (
            .O(N__19623),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    CascadeMux I__1946 (
            .O(N__19616),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_ ));
    InMux I__1945 (
            .O(N__19613),
            .I(N__19610));
    LocalMux I__1944 (
            .O(N__19610),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3 ));
    CascadeMux I__1943 (
            .O(N__19607),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_ ));
    InMux I__1942 (
            .O(N__19604),
            .I(N__19601));
    LocalMux I__1941 (
            .O(N__19601),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17 ));
    InMux I__1940 (
            .O(N__19598),
            .I(N__19595));
    LocalMux I__1939 (
            .O(N__19595),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ));
    CascadeMux I__1938 (
            .O(N__19592),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_ ));
    InMux I__1937 (
            .O(N__19589),
            .I(N__19586));
    LocalMux I__1936 (
            .O(N__19586),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_2 ));
    CascadeMux I__1935 (
            .O(N__19583),
            .I(\current_shift_inst.PI_CTRL.N_77_cascade_ ));
    InMux I__1934 (
            .O(N__19580),
            .I(N__19577));
    LocalMux I__1933 (
            .O(N__19577),
            .I(\current_shift_inst.PI_CTRL.N_43 ));
    InMux I__1932 (
            .O(N__19574),
            .I(N__19571));
    LocalMux I__1931 (
            .O(N__19571),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ));
    CascadeMux I__1930 (
            .O(N__19568),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_ ));
    InMux I__1929 (
            .O(N__19565),
            .I(N__19562));
    LocalMux I__1928 (
            .O(N__19562),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ));
    CascadeMux I__1927 (
            .O(N__19559),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_ ));
    CascadeMux I__1926 (
            .O(N__19556),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ));
    CascadeMux I__1925 (
            .O(N__19553),
            .I(\current_shift_inst.PI_CTRL.N_44_cascade_ ));
    InMux I__1924 (
            .O(N__19550),
            .I(N__19547));
    LocalMux I__1923 (
            .O(N__19547),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ));
    InMux I__1922 (
            .O(N__19544),
            .I(N__19541));
    LocalMux I__1921 (
            .O(N__19541),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ));
    CascadeMux I__1920 (
            .O(N__19538),
            .I(N__19535));
    InMux I__1919 (
            .O(N__19535),
            .I(N__19532));
    LocalMux I__1918 (
            .O(N__19532),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    InMux I__1917 (
            .O(N__19529),
            .I(N__19526));
    LocalMux I__1916 (
            .O(N__19526),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    CascadeMux I__1915 (
            .O(N__19523),
            .I(N__19520));
    InMux I__1914 (
            .O(N__19520),
            .I(N__19517));
    LocalMux I__1913 (
            .O(N__19517),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    CascadeMux I__1912 (
            .O(N__19514),
            .I(N__19511));
    InMux I__1911 (
            .O(N__19511),
            .I(N__19508));
    LocalMux I__1910 (
            .O(N__19508),
            .I(N__19505));
    Odrv4 I__1909 (
            .O(N__19505),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    CascadeMux I__1908 (
            .O(N__19502),
            .I(N__19499));
    InMux I__1907 (
            .O(N__19499),
            .I(N__19496));
    LocalMux I__1906 (
            .O(N__19496),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    InMux I__1905 (
            .O(N__19493),
            .I(N__19490));
    LocalMux I__1904 (
            .O(N__19490),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ));
    InMux I__1903 (
            .O(N__19487),
            .I(N__19484));
    LocalMux I__1902 (
            .O(N__19484),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    CascadeMux I__1901 (
            .O(N__19481),
            .I(N__19478));
    InMux I__1900 (
            .O(N__19478),
            .I(N__19475));
    LocalMux I__1899 (
            .O(N__19475),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    InMux I__1898 (
            .O(N__19472),
            .I(N__19469));
    LocalMux I__1897 (
            .O(N__19469),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    InMux I__1896 (
            .O(N__19466),
            .I(N__19463));
    LocalMux I__1895 (
            .O(N__19463),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    InMux I__1894 (
            .O(N__19460),
            .I(N__19457));
    LocalMux I__1893 (
            .O(N__19457),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    InMux I__1892 (
            .O(N__19454),
            .I(N__19451));
    LocalMux I__1891 (
            .O(N__19451),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    InMux I__1890 (
            .O(N__19448),
            .I(N__19445));
    LocalMux I__1889 (
            .O(N__19445),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    CascadeMux I__1888 (
            .O(N__19442),
            .I(N__19439));
    InMux I__1887 (
            .O(N__19439),
            .I(N__19436));
    LocalMux I__1886 (
            .O(N__19436),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    InMux I__1885 (
            .O(N__19433),
            .I(N__19430));
    LocalMux I__1884 (
            .O(N__19430),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    CascadeMux I__1883 (
            .O(N__19427),
            .I(N__19424));
    InMux I__1882 (
            .O(N__19424),
            .I(N__19421));
    LocalMux I__1881 (
            .O(N__19421),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    InMux I__1880 (
            .O(N__19418),
            .I(N__19415));
    LocalMux I__1879 (
            .O(N__19415),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    InMux I__1878 (
            .O(N__19412),
            .I(N__19409));
    LocalMux I__1877 (
            .O(N__19409),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    InMux I__1876 (
            .O(N__19406),
            .I(N__19403));
    LocalMux I__1875 (
            .O(N__19403),
            .I(N__19400));
    Span4Mux_v I__1874 (
            .O(N__19400),
            .I(N__19397));
    Span4Mux_v I__1873 (
            .O(N__19397),
            .I(N__19394));
    Odrv4 I__1872 (
            .O(N__19394),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ));
    CascadeMux I__1871 (
            .O(N__19391),
            .I(N__19388));
    InMux I__1870 (
            .O(N__19388),
            .I(N__19385));
    LocalMux I__1869 (
            .O(N__19385),
            .I(N__19382));
    Span4Mux_v I__1868 (
            .O(N__19382),
            .I(N__19379));
    Odrv4 I__1867 (
            .O(N__19379),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ));
    InMux I__1866 (
            .O(N__19376),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ));
    InMux I__1865 (
            .O(N__19373),
            .I(N__19370));
    LocalMux I__1864 (
            .O(N__19370),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    CascadeMux I__1863 (
            .O(N__19367),
            .I(N__19364));
    InMux I__1862 (
            .O(N__19364),
            .I(N__19361));
    LocalMux I__1861 (
            .O(N__19361),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    CascadeMux I__1860 (
            .O(N__19358),
            .I(N__19355));
    InMux I__1859 (
            .O(N__19355),
            .I(N__19352));
    LocalMux I__1858 (
            .O(N__19352),
            .I(N__19349));
    Odrv4 I__1857 (
            .O(N__19349),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    InMux I__1856 (
            .O(N__19346),
            .I(N__19343));
    LocalMux I__1855 (
            .O(N__19343),
            .I(N__19340));
    Odrv4 I__1854 (
            .O(N__19340),
            .I(N_38_i_i));
    InMux I__1853 (
            .O(N__19337),
            .I(N__19334));
    LocalMux I__1852 (
            .O(N__19334),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ));
    InMux I__1851 (
            .O(N__19331),
            .I(N__19328));
    LocalMux I__1850 (
            .O(N__19328),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ));
    CascadeMux I__1849 (
            .O(N__19325),
            .I(N__19322));
    InMux I__1848 (
            .O(N__19322),
            .I(N__19319));
    LocalMux I__1847 (
            .O(N__19319),
            .I(N__19316));
    Span4Mux_v I__1846 (
            .O(N__19316),
            .I(N__19313));
    Odrv4 I__1845 (
            .O(N__19313),
            .I(\current_shift_inst.PI_CTRL.integrator_1_23 ));
    InMux I__1844 (
            .O(N__19310),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ));
    InMux I__1843 (
            .O(N__19307),
            .I(N__19304));
    LocalMux I__1842 (
            .O(N__19304),
            .I(N__19301));
    Span4Mux_v I__1841 (
            .O(N__19301),
            .I(N__19298));
    Odrv4 I__1840 (
            .O(N__19298),
            .I(\current_shift_inst.PI_CTRL.integrator_1_24 ));
    InMux I__1839 (
            .O(N__19295),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ));
    CascadeMux I__1838 (
            .O(N__19292),
            .I(N__19289));
    InMux I__1837 (
            .O(N__19289),
            .I(N__19286));
    LocalMux I__1836 (
            .O(N__19286),
            .I(N__19283));
    Span4Mux_h I__1835 (
            .O(N__19283),
            .I(N__19280));
    Span4Mux_v I__1834 (
            .O(N__19280),
            .I(N__19277));
    Odrv4 I__1833 (
            .O(N__19277),
            .I(\current_shift_inst.PI_CTRL.integrator_1_25 ));
    InMux I__1832 (
            .O(N__19274),
            .I(bfn_3_16_0_));
    CascadeMux I__1831 (
            .O(N__19271),
            .I(N__19268));
    InMux I__1830 (
            .O(N__19268),
            .I(N__19265));
    LocalMux I__1829 (
            .O(N__19265),
            .I(N__19262));
    Span4Mux_v I__1828 (
            .O(N__19262),
            .I(N__19259));
    Odrv4 I__1827 (
            .O(N__19259),
            .I(\current_shift_inst.PI_CTRL.integrator_1_26 ));
    InMux I__1826 (
            .O(N__19256),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ));
    CascadeMux I__1825 (
            .O(N__19253),
            .I(N__19250));
    InMux I__1824 (
            .O(N__19250),
            .I(N__19247));
    LocalMux I__1823 (
            .O(N__19247),
            .I(N__19244));
    Span4Mux_h I__1822 (
            .O(N__19244),
            .I(N__19241));
    Span4Mux_v I__1821 (
            .O(N__19241),
            .I(N__19238));
    Odrv4 I__1820 (
            .O(N__19238),
            .I(\current_shift_inst.PI_CTRL.integrator_1_27 ));
    CascadeMux I__1819 (
            .O(N__19235),
            .I(N__19232));
    InMux I__1818 (
            .O(N__19232),
            .I(N__19229));
    LocalMux I__1817 (
            .O(N__19229),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    InMux I__1816 (
            .O(N__19226),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ));
    CascadeMux I__1815 (
            .O(N__19223),
            .I(N__19220));
    InMux I__1814 (
            .O(N__19220),
            .I(N__19217));
    LocalMux I__1813 (
            .O(N__19217),
            .I(N__19214));
    Span4Mux_h I__1812 (
            .O(N__19214),
            .I(N__19211));
    Span4Mux_v I__1811 (
            .O(N__19211),
            .I(N__19208));
    Odrv4 I__1810 (
            .O(N__19208),
            .I(\current_shift_inst.PI_CTRL.integrator_1_28 ));
    InMux I__1809 (
            .O(N__19205),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ));
    CascadeMux I__1808 (
            .O(N__19202),
            .I(N__19199));
    InMux I__1807 (
            .O(N__19199),
            .I(N__19196));
    LocalMux I__1806 (
            .O(N__19196),
            .I(N__19193));
    Span4Mux_v I__1805 (
            .O(N__19193),
            .I(N__19190));
    Odrv4 I__1804 (
            .O(N__19190),
            .I(\current_shift_inst.PI_CTRL.integrator_1_29 ));
    InMux I__1803 (
            .O(N__19187),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ));
    InMux I__1802 (
            .O(N__19184),
            .I(N__19181));
    LocalMux I__1801 (
            .O(N__19181),
            .I(N__19178));
    Span4Mux_v I__1800 (
            .O(N__19178),
            .I(N__19175));
    Odrv4 I__1799 (
            .O(N__19175),
            .I(\current_shift_inst.PI_CTRL.integrator_1_30 ));
    InMux I__1798 (
            .O(N__19172),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ));
    CascadeMux I__1797 (
            .O(N__19169),
            .I(N__19166));
    InMux I__1796 (
            .O(N__19166),
            .I(N__19163));
    LocalMux I__1795 (
            .O(N__19163),
            .I(N__19160));
    Span4Mux_h I__1794 (
            .O(N__19160),
            .I(N__19157));
    Odrv4 I__1793 (
            .O(N__19157),
            .I(\current_shift_inst.PI_CTRL.integrator_1_14 ));
    InMux I__1792 (
            .O(N__19154),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ));
    CascadeMux I__1791 (
            .O(N__19151),
            .I(N__19148));
    InMux I__1790 (
            .O(N__19148),
            .I(N__19145));
    LocalMux I__1789 (
            .O(N__19145),
            .I(N__19142));
    Span4Mux_v I__1788 (
            .O(N__19142),
            .I(N__19139));
    Odrv4 I__1787 (
            .O(N__19139),
            .I(\current_shift_inst.PI_CTRL.integrator_1_15 ));
    InMux I__1786 (
            .O(N__19136),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ));
    CascadeMux I__1785 (
            .O(N__19133),
            .I(N__19130));
    InMux I__1784 (
            .O(N__19130),
            .I(N__19127));
    LocalMux I__1783 (
            .O(N__19127),
            .I(N__19124));
    Span4Mux_v I__1782 (
            .O(N__19124),
            .I(N__19121));
    Odrv4 I__1781 (
            .O(N__19121),
            .I(\current_shift_inst.PI_CTRL.integrator_1_16 ));
    InMux I__1780 (
            .O(N__19118),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ));
    CascadeMux I__1779 (
            .O(N__19115),
            .I(N__19112));
    InMux I__1778 (
            .O(N__19112),
            .I(N__19109));
    LocalMux I__1777 (
            .O(N__19109),
            .I(N__19106));
    Span4Mux_h I__1776 (
            .O(N__19106),
            .I(N__19103));
    Span4Mux_v I__1775 (
            .O(N__19103),
            .I(N__19100));
    Odrv4 I__1774 (
            .O(N__19100),
            .I(\current_shift_inst.PI_CTRL.integrator_1_17 ));
    InMux I__1773 (
            .O(N__19097),
            .I(bfn_3_15_0_));
    CascadeMux I__1772 (
            .O(N__19094),
            .I(N__19091));
    InMux I__1771 (
            .O(N__19091),
            .I(N__19088));
    LocalMux I__1770 (
            .O(N__19088),
            .I(N__19085));
    Span4Mux_v I__1769 (
            .O(N__19085),
            .I(N__19082));
    Odrv4 I__1768 (
            .O(N__19082),
            .I(\current_shift_inst.PI_CTRL.integrator_1_18 ));
    InMux I__1767 (
            .O(N__19079),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ));
    CascadeMux I__1766 (
            .O(N__19076),
            .I(N__19073));
    InMux I__1765 (
            .O(N__19073),
            .I(N__19070));
    LocalMux I__1764 (
            .O(N__19070),
            .I(N__19067));
    Span4Mux_h I__1763 (
            .O(N__19067),
            .I(N__19064));
    Span4Mux_v I__1762 (
            .O(N__19064),
            .I(N__19061));
    Odrv4 I__1761 (
            .O(N__19061),
            .I(\current_shift_inst.PI_CTRL.integrator_1_19 ));
    InMux I__1760 (
            .O(N__19058),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ));
    CascadeMux I__1759 (
            .O(N__19055),
            .I(N__19052));
    InMux I__1758 (
            .O(N__19052),
            .I(N__19049));
    LocalMux I__1757 (
            .O(N__19049),
            .I(N__19046));
    Span12Mux_h I__1756 (
            .O(N__19046),
            .I(N__19043));
    Odrv12 I__1755 (
            .O(N__19043),
            .I(\current_shift_inst.PI_CTRL.integrator_1_20 ));
    InMux I__1754 (
            .O(N__19040),
            .I(N__19037));
    LocalMux I__1753 (
            .O(N__19037),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    InMux I__1752 (
            .O(N__19034),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ));
    CascadeMux I__1751 (
            .O(N__19031),
            .I(N__19028));
    InMux I__1750 (
            .O(N__19028),
            .I(N__19025));
    LocalMux I__1749 (
            .O(N__19025),
            .I(N__19022));
    Span4Mux_v I__1748 (
            .O(N__19022),
            .I(N__19019));
    Odrv4 I__1747 (
            .O(N__19019),
            .I(\current_shift_inst.PI_CTRL.integrator_1_21 ));
    InMux I__1746 (
            .O(N__19016),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ));
    CascadeMux I__1745 (
            .O(N__19013),
            .I(N__19010));
    InMux I__1744 (
            .O(N__19010),
            .I(N__19007));
    LocalMux I__1743 (
            .O(N__19007),
            .I(N__19004));
    Span4Mux_v I__1742 (
            .O(N__19004),
            .I(N__19001));
    Odrv4 I__1741 (
            .O(N__19001),
            .I(\current_shift_inst.PI_CTRL.integrator_1_22 ));
    InMux I__1740 (
            .O(N__18998),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ));
    CascadeMux I__1739 (
            .O(N__18995),
            .I(N__18992));
    InMux I__1738 (
            .O(N__18992),
            .I(N__18989));
    LocalMux I__1737 (
            .O(N__18989),
            .I(N__18986));
    Span4Mux_h I__1736 (
            .O(N__18986),
            .I(N__18983));
    Odrv4 I__1735 (
            .O(N__18983),
            .I(\current_shift_inst.PI_CTRL.integrator_1_6 ));
    InMux I__1734 (
            .O(N__18980),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ));
    CascadeMux I__1733 (
            .O(N__18977),
            .I(N__18974));
    InMux I__1732 (
            .O(N__18974),
            .I(N__18971));
    LocalMux I__1731 (
            .O(N__18971),
            .I(N__18968));
    Span4Mux_h I__1730 (
            .O(N__18968),
            .I(N__18965));
    Odrv4 I__1729 (
            .O(N__18965),
            .I(\current_shift_inst.PI_CTRL.integrator_1_7 ));
    InMux I__1728 (
            .O(N__18962),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ));
    CascadeMux I__1727 (
            .O(N__18959),
            .I(N__18956));
    InMux I__1726 (
            .O(N__18956),
            .I(N__18953));
    LocalMux I__1725 (
            .O(N__18953),
            .I(N__18950));
    Span4Mux_h I__1724 (
            .O(N__18950),
            .I(N__18947));
    Odrv4 I__1723 (
            .O(N__18947),
            .I(\current_shift_inst.PI_CTRL.integrator_1_8 ));
    InMux I__1722 (
            .O(N__18944),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ));
    CascadeMux I__1721 (
            .O(N__18941),
            .I(N__18938));
    InMux I__1720 (
            .O(N__18938),
            .I(N__18935));
    LocalMux I__1719 (
            .O(N__18935),
            .I(N__18932));
    Span4Mux_v I__1718 (
            .O(N__18932),
            .I(N__18929));
    Odrv4 I__1717 (
            .O(N__18929),
            .I(\current_shift_inst.PI_CTRL.integrator_1_9 ));
    CascadeMux I__1716 (
            .O(N__18926),
            .I(N__18923));
    InMux I__1715 (
            .O(N__18923),
            .I(N__18920));
    LocalMux I__1714 (
            .O(N__18920),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    InMux I__1713 (
            .O(N__18917),
            .I(bfn_3_14_0_));
    CascadeMux I__1712 (
            .O(N__18914),
            .I(N__18911));
    InMux I__1711 (
            .O(N__18911),
            .I(N__18908));
    LocalMux I__1710 (
            .O(N__18908),
            .I(N__18905));
    Span4Mux_v I__1709 (
            .O(N__18905),
            .I(N__18902));
    Odrv4 I__1708 (
            .O(N__18902),
            .I(\current_shift_inst.PI_CTRL.integrator_1_10 ));
    InMux I__1707 (
            .O(N__18899),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ));
    CascadeMux I__1706 (
            .O(N__18896),
            .I(N__18893));
    InMux I__1705 (
            .O(N__18893),
            .I(N__18890));
    LocalMux I__1704 (
            .O(N__18890),
            .I(N__18887));
    Span4Mux_v I__1703 (
            .O(N__18887),
            .I(N__18884));
    Odrv4 I__1702 (
            .O(N__18884),
            .I(\current_shift_inst.PI_CTRL.integrator_1_11 ));
    InMux I__1701 (
            .O(N__18881),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ));
    InMux I__1700 (
            .O(N__18878),
            .I(N__18875));
    LocalMux I__1699 (
            .O(N__18875),
            .I(N__18872));
    Span4Mux_h I__1698 (
            .O(N__18872),
            .I(N__18869));
    Odrv4 I__1697 (
            .O(N__18869),
            .I(\current_shift_inst.PI_CTRL.integrator_1_12 ));
    InMux I__1696 (
            .O(N__18866),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ));
    CascadeMux I__1695 (
            .O(N__18863),
            .I(N__18860));
    InMux I__1694 (
            .O(N__18860),
            .I(N__18857));
    LocalMux I__1693 (
            .O(N__18857),
            .I(N__18854));
    Span4Mux_h I__1692 (
            .O(N__18854),
            .I(N__18851));
    Odrv4 I__1691 (
            .O(N__18851),
            .I(\current_shift_inst.PI_CTRL.integrator_1_13 ));
    InMux I__1690 (
            .O(N__18848),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ));
    InMux I__1689 (
            .O(N__18845),
            .I(N__18842));
    LocalMux I__1688 (
            .O(N__18842),
            .I(N__18839));
    Odrv4 I__1687 (
            .O(N__18839),
            .I(rgb_drv_RNOZ0));
    ClkMux I__1686 (
            .O(N__18836),
            .I(N__18830));
    ClkMux I__1685 (
            .O(N__18835),
            .I(N__18830));
    GlobalMux I__1684 (
            .O(N__18830),
            .I(N__18827));
    gio2CtrlBuf I__1683 (
            .O(N__18827),
            .I(delay_hc_input_c_g));
    CascadeMux I__1682 (
            .O(N__18824),
            .I(N__18821));
    InMux I__1681 (
            .O(N__18821),
            .I(N__18817));
    InMux I__1680 (
            .O(N__18820),
            .I(N__18814));
    LocalMux I__1679 (
            .O(N__18817),
            .I(N__18809));
    LocalMux I__1678 (
            .O(N__18814),
            .I(N__18809));
    Span4Mux_v I__1677 (
            .O(N__18809),
            .I(N__18806));
    Odrv4 I__1676 (
            .O(N__18806),
            .I(\current_shift_inst.PI_CTRL.un1_integrator ));
    CascadeMux I__1675 (
            .O(N__18803),
            .I(N__18800));
    InMux I__1674 (
            .O(N__18800),
            .I(N__18797));
    LocalMux I__1673 (
            .O(N__18797),
            .I(N__18794));
    Span4Mux_v I__1672 (
            .O(N__18794),
            .I(N__18791));
    Odrv4 I__1671 (
            .O(N__18791),
            .I(\current_shift_inst.PI_CTRL.integrator_1_2 ));
    InMux I__1670 (
            .O(N__18788),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ));
    CascadeMux I__1669 (
            .O(N__18785),
            .I(N__18782));
    InMux I__1668 (
            .O(N__18782),
            .I(N__18779));
    LocalMux I__1667 (
            .O(N__18779),
            .I(N__18776));
    Span4Mux_v I__1666 (
            .O(N__18776),
            .I(N__18773));
    Odrv4 I__1665 (
            .O(N__18773),
            .I(\current_shift_inst.PI_CTRL.integrator_1_3 ));
    InMux I__1664 (
            .O(N__18770),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ));
    CascadeMux I__1663 (
            .O(N__18767),
            .I(N__18764));
    InMux I__1662 (
            .O(N__18764),
            .I(N__18761));
    LocalMux I__1661 (
            .O(N__18761),
            .I(N__18758));
    Span4Mux_v I__1660 (
            .O(N__18758),
            .I(N__18755));
    Odrv4 I__1659 (
            .O(N__18755),
            .I(\current_shift_inst.PI_CTRL.integrator_1_4 ));
    CascadeMux I__1658 (
            .O(N__18752),
            .I(N__18749));
    InMux I__1657 (
            .O(N__18749),
            .I(N__18746));
    LocalMux I__1656 (
            .O(N__18746),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    InMux I__1655 (
            .O(N__18743),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ));
    CascadeMux I__1654 (
            .O(N__18740),
            .I(N__18737));
    InMux I__1653 (
            .O(N__18737),
            .I(N__18734));
    LocalMux I__1652 (
            .O(N__18734),
            .I(N__18731));
    Span4Mux_h I__1651 (
            .O(N__18731),
            .I(N__18728));
    Odrv4 I__1650 (
            .O(N__18728),
            .I(\current_shift_inst.PI_CTRL.integrator_1_5 ));
    InMux I__1649 (
            .O(N__18725),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ));
    InMux I__1648 (
            .O(N__18722),
            .I(N__18719));
    LocalMux I__1647 (
            .O(N__18719),
            .I(N__18716));
    Span4Mux_v I__1646 (
            .O(N__18716),
            .I(N__18713));
    Odrv4 I__1645 (
            .O(N__18713),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_11 ));
    InMux I__1644 (
            .O(N__18710),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ));
    InMux I__1643 (
            .O(N__18707),
            .I(N__18704));
    LocalMux I__1642 (
            .O(N__18704),
            .I(N__18701));
    Span4Mux_v I__1641 (
            .O(N__18701),
            .I(N__18698));
    Odrv4 I__1640 (
            .O(N__18698),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_12 ));
    InMux I__1639 (
            .O(N__18695),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ));
    InMux I__1638 (
            .O(N__18692),
            .I(N__18689));
    LocalMux I__1637 (
            .O(N__18689),
            .I(N__18686));
    Span4Mux_v I__1636 (
            .O(N__18686),
            .I(N__18683));
    Odrv4 I__1635 (
            .O(N__18683),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_13 ));
    InMux I__1634 (
            .O(N__18680),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ));
    InMux I__1633 (
            .O(N__18677),
            .I(N__18674));
    LocalMux I__1632 (
            .O(N__18674),
            .I(N__18671));
    Span4Mux_v I__1631 (
            .O(N__18671),
            .I(N__18668));
    Odrv4 I__1630 (
            .O(N__18668),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_14 ));
    InMux I__1629 (
            .O(N__18665),
            .I(N__18651));
    CascadeMux I__1628 (
            .O(N__18664),
            .I(N__18648));
    CascadeMux I__1627 (
            .O(N__18663),
            .I(N__18645));
    CascadeMux I__1626 (
            .O(N__18662),
            .I(N__18642));
    CascadeMux I__1625 (
            .O(N__18661),
            .I(N__18639));
    CascadeMux I__1624 (
            .O(N__18660),
            .I(N__18636));
    CascadeMux I__1623 (
            .O(N__18659),
            .I(N__18633));
    CascadeMux I__1622 (
            .O(N__18658),
            .I(N__18630));
    CascadeMux I__1621 (
            .O(N__18657),
            .I(N__18627));
    CascadeMux I__1620 (
            .O(N__18656),
            .I(N__18624));
    CascadeMux I__1619 (
            .O(N__18655),
            .I(N__18621));
    CascadeMux I__1618 (
            .O(N__18654),
            .I(N__18618));
    LocalMux I__1617 (
            .O(N__18651),
            .I(N__18615));
    InMux I__1616 (
            .O(N__18648),
            .I(N__18608));
    InMux I__1615 (
            .O(N__18645),
            .I(N__18608));
    InMux I__1614 (
            .O(N__18642),
            .I(N__18608));
    InMux I__1613 (
            .O(N__18639),
            .I(N__18599));
    InMux I__1612 (
            .O(N__18636),
            .I(N__18599));
    InMux I__1611 (
            .O(N__18633),
            .I(N__18599));
    InMux I__1610 (
            .O(N__18630),
            .I(N__18599));
    InMux I__1609 (
            .O(N__18627),
            .I(N__18594));
    InMux I__1608 (
            .O(N__18624),
            .I(N__18594));
    InMux I__1607 (
            .O(N__18621),
            .I(N__18589));
    InMux I__1606 (
            .O(N__18618),
            .I(N__18589));
    Odrv4 I__1605 (
            .O(N__18615),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    LocalMux I__1604 (
            .O(N__18608),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    LocalMux I__1603 (
            .O(N__18599),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    LocalMux I__1602 (
            .O(N__18594),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    LocalMux I__1601 (
            .O(N__18589),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    InMux I__1600 (
            .O(N__18578),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ));
    InMux I__1599 (
            .O(N__18575),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ));
    InMux I__1598 (
            .O(N__18572),
            .I(N__18569));
    LocalMux I__1597 (
            .O(N__18569),
            .I(N__18566));
    Span4Mux_v I__1596 (
            .O(N__18566),
            .I(N__18563));
    Odrv4 I__1595 (
            .O(N__18563),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_3 ));
    CascadeMux I__1594 (
            .O(N__18560),
            .I(N__18557));
    InMux I__1593 (
            .O(N__18557),
            .I(N__18554));
    LocalMux I__1592 (
            .O(N__18554),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_18 ));
    InMux I__1591 (
            .O(N__18551),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ));
    InMux I__1590 (
            .O(N__18548),
            .I(N__18545));
    LocalMux I__1589 (
            .O(N__18545),
            .I(N__18542));
    Span4Mux_v I__1588 (
            .O(N__18542),
            .I(N__18539));
    Odrv4 I__1587 (
            .O(N__18539),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_4 ));
    InMux I__1586 (
            .O(N__18536),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ));
    InMux I__1585 (
            .O(N__18533),
            .I(N__18530));
    LocalMux I__1584 (
            .O(N__18530),
            .I(N__18527));
    Span4Mux_v I__1583 (
            .O(N__18527),
            .I(N__18524));
    Odrv4 I__1582 (
            .O(N__18524),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_5 ));
    InMux I__1581 (
            .O(N__18521),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ));
    InMux I__1580 (
            .O(N__18518),
            .I(N__18515));
    LocalMux I__1579 (
            .O(N__18515),
            .I(N__18512));
    Span4Mux_v I__1578 (
            .O(N__18512),
            .I(N__18509));
    Odrv4 I__1577 (
            .O(N__18509),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_6 ));
    InMux I__1576 (
            .O(N__18506),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ));
    InMux I__1575 (
            .O(N__18503),
            .I(N__18500));
    LocalMux I__1574 (
            .O(N__18500),
            .I(N__18497));
    Span4Mux_v I__1573 (
            .O(N__18497),
            .I(N__18494));
    Odrv4 I__1572 (
            .O(N__18494),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_7 ));
    InMux I__1571 (
            .O(N__18491),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ));
    InMux I__1570 (
            .O(N__18488),
            .I(N__18485));
    LocalMux I__1569 (
            .O(N__18485),
            .I(N__18482));
    Span4Mux_v I__1568 (
            .O(N__18482),
            .I(N__18479));
    Odrv4 I__1567 (
            .O(N__18479),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_8 ));
    InMux I__1566 (
            .O(N__18476),
            .I(bfn_1_12_0_));
    InMux I__1565 (
            .O(N__18473),
            .I(N__18470));
    LocalMux I__1564 (
            .O(N__18470),
            .I(N__18467));
    Span4Mux_v I__1563 (
            .O(N__18467),
            .I(N__18464));
    Odrv4 I__1562 (
            .O(N__18464),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_9 ));
    InMux I__1561 (
            .O(N__18461),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ));
    InMux I__1560 (
            .O(N__18458),
            .I(N__18455));
    LocalMux I__1559 (
            .O(N__18455),
            .I(N__18452));
    Span4Mux_v I__1558 (
            .O(N__18452),
            .I(N__18449));
    Odrv4 I__1557 (
            .O(N__18449),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_10 ));
    InMux I__1556 (
            .O(N__18446),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ));
    InMux I__1555 (
            .O(N__18443),
            .I(N__18440));
    LocalMux I__1554 (
            .O(N__18440),
            .I(N__18437));
    Span4Mux_v I__1553 (
            .O(N__18437),
            .I(N__18434));
    Odrv4 I__1552 (
            .O(N__18434),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_15 ));
    InMux I__1551 (
            .O(N__18431),
            .I(N__18428));
    LocalMux I__1550 (
            .O(N__18428),
            .I(N__18425));
    Span4Mux_v I__1549 (
            .O(N__18425),
            .I(N__18422));
    Odrv4 I__1548 (
            .O(N__18422),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_0 ));
    CascadeMux I__1547 (
            .O(N__18419),
            .I(N__18416));
    InMux I__1546 (
            .O(N__18416),
            .I(N__18413));
    LocalMux I__1545 (
            .O(N__18413),
            .I(N__18410));
    Odrv4 I__1544 (
            .O(N__18410),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_15 ));
    InMux I__1543 (
            .O(N__18407),
            .I(N__18404));
    LocalMux I__1542 (
            .O(N__18404),
            .I(N__18401));
    Span4Mux_v I__1541 (
            .O(N__18401),
            .I(N__18398));
    Odrv4 I__1540 (
            .O(N__18398),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_1 ));
    CascadeMux I__1539 (
            .O(N__18395),
            .I(N__18392));
    InMux I__1538 (
            .O(N__18392),
            .I(N__18389));
    LocalMux I__1537 (
            .O(N__18389),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_16 ));
    InMux I__1536 (
            .O(N__18386),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ));
    InMux I__1535 (
            .O(N__18383),
            .I(N__18380));
    LocalMux I__1534 (
            .O(N__18380),
            .I(N__18377));
    Span4Mux_v I__1533 (
            .O(N__18377),
            .I(N__18374));
    Odrv4 I__1532 (
            .O(N__18374),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_2 ));
    CascadeMux I__1531 (
            .O(N__18371),
            .I(N__18368));
    InMux I__1530 (
            .O(N__18368),
            .I(N__18365));
    LocalMux I__1529 (
            .O(N__18365),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_17 ));
    InMux I__1528 (
            .O(N__18362),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ));
    IoInMux I__1527 (
            .O(N__18359),
            .I(N__18356));
    LocalMux I__1526 (
            .O(N__18356),
            .I(N__18353));
    Span4Mux_s1_v I__1525 (
            .O(N__18353),
            .I(N__18350));
    Span4Mux_h I__1524 (
            .O(N__18350),
            .I(N__18347));
    Sp12to4 I__1523 (
            .O(N__18347),
            .I(N__18344));
    Span12Mux_s9_v I__1522 (
            .O(N__18344),
            .I(N__18341));
    Span12Mux_v I__1521 (
            .O(N__18341),
            .I(N__18338));
    Odrv12 I__1520 (
            .O(N__18338),
            .I(delay_tr_input_ibuf_gb_io_gb_input));
    IoInMux I__1519 (
            .O(N__18335),
            .I(N__18332));
    LocalMux I__1518 (
            .O(N__18332),
            .I(N__18329));
    IoSpan4Mux I__1517 (
            .O(N__18329),
            .I(N__18326));
    IoSpan4Mux I__1516 (
            .O(N__18326),
            .I(N__18323));
    Odrv4 I__1515 (
            .O(N__18323),
            .I(delay_hc_input_ibuf_gb_io_gb_input));
    defparam IN_MUX_bfv_14_28_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_28_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_28_0_));
    defparam IN_MUX_bfv_14_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_29_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_7 ),
            .carryinitout(bfn_14_29_0_));
    defparam IN_MUX_bfv_14_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_30_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_15 ),
            .carryinitout(bfn_14_30_0_));
    defparam IN_MUX_bfv_14_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_10_0_));
    defparam IN_MUX_bfv_14_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_11_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_14_11_0_));
    defparam IN_MUX_bfv_14_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_12_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_14_12_0_));
    defparam IN_MUX_bfv_14_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_13_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_14_13_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_11_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_12_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_11_12_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_17_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_12_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_17_12_0_));
    defparam IN_MUX_bfv_17_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_13_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_17_13_0_));
    defparam IN_MUX_bfv_17_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_17_14_0_));
    defparam IN_MUX_bfv_12_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_6_0_));
    defparam IN_MUX_bfv_12_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_7_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_12_7_0_));
    defparam IN_MUX_bfv_12_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_8_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_12_8_0_));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_12_9_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_11_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_16_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .carryinitout(bfn_11_16_0_));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_12_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_13_0_));
    defparam IN_MUX_bfv_12_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_14_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .carryinitout(bfn_12_14_0_));
    defparam IN_MUX_bfv_12_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_15_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .carryinitout(bfn_12_15_0_));
    defparam IN_MUX_bfv_12_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_16_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .carryinitout(bfn_12_16_0_));
    defparam IN_MUX_bfv_9_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_16_0_));
    defparam IN_MUX_bfv_9_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_17_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_7 ),
            .carryinitout(bfn_9_17_0_));
    defparam IN_MUX_bfv_9_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_18_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_15 ),
            .carryinitout(bfn_9_18_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_23 ),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_3_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_13_0_));
    defparam IN_MUX_bfv_3_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_14_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .carryinitout(bfn_3_14_0_));
    defparam IN_MUX_bfv_3_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_15_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .carryinitout(bfn_3_15_0_));
    defparam IN_MUX_bfv_3_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_16_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .carryinitout(bfn_3_16_0_));
    defparam IN_MUX_bfv_15_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_23_0_));
    defparam IN_MUX_bfv_15_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_24_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryinitout(bfn_15_24_0_));
    defparam IN_MUX_bfv_15_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_25_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryinitout(bfn_15_25_0_));
    defparam IN_MUX_bfv_15_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_26_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryinitout(bfn_15_26_0_));
    defparam IN_MUX_bfv_13_28_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_28_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_28_0_));
    defparam IN_MUX_bfv_13_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_29_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .carryinitout(bfn_13_29_0_));
    defparam IN_MUX_bfv_13_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_30_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_15 ),
            .carryinitout(bfn_13_30_0_));
    defparam IN_MUX_bfv_13_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_24_0_));
    defparam IN_MUX_bfv_13_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_25_0_ (
            .carryinitin(\pwm_generator_inst.un19_threshold_cry_7 ),
            .carryinitout(bfn_13_25_0_));
    defparam IN_MUX_bfv_14_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_25_0_));
    defparam IN_MUX_bfv_14_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_26_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_1_cry_7 ),
            .carryinitout(bfn_14_26_0_));
    defparam IN_MUX_bfv_14_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_27_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_1_cry_15 ),
            .carryinitout(bfn_14_27_0_));
    defparam IN_MUX_bfv_11_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_23_0_));
    defparam IN_MUX_bfv_11_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_24_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_11_24_0_));
    defparam IN_MUX_bfv_12_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_21_0_));
    defparam IN_MUX_bfv_12_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_22_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_12_22_0_));
    defparam IN_MUX_bfv_14_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_7_0_));
    defparam IN_MUX_bfv_14_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_8_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un4_running_cry_8 ),
            .carryinitout(bfn_14_8_0_));
    defparam IN_MUX_bfv_14_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_9_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un4_running_cry_16 ),
            .carryinitout(bfn_14_9_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_9_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_12_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un4_running_cry_8 ),
            .carryinitout(bfn_9_12_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un4_running_cry_16 ),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_18_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_10_0_));
    defparam IN_MUX_bfv_18_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_11_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un4_running_cry_8 ),
            .carryinitout(bfn_18_11_0_));
    defparam IN_MUX_bfv_18_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_12_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un4_running_cry_16 ),
            .carryinitout(bfn_18_12_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_7_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un4_running_cry_8 ),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un4_running_cry_16 ),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_15_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_14_0_));
    defparam IN_MUX_bfv_15_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_15_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_15_15_0_));
    defparam IN_MUX_bfv_15_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_16_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_15_16_0_));
    defparam IN_MUX_bfv_15_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_17_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_15_17_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_8_12_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_8_10_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_7 ),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_7_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_20_0_));
    defparam IN_MUX_bfv_7_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_21_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_7_21_0_));
    defparam IN_MUX_bfv_7_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_22_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_7_22_0_));
    defparam IN_MUX_bfv_7_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_23_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_7_23_0_));
    defparam IN_MUX_bfv_10_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_18_0_));
    defparam IN_MUX_bfv_10_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_19_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_8 ),
            .carryinitout(bfn_10_19_0_));
    defparam IN_MUX_bfv_10_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_20_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_16 ),
            .carryinitout(bfn_10_20_0_));
    defparam IN_MUX_bfv_10_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_21_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_24 ),
            .carryinitout(bfn_10_21_0_));
    defparam IN_MUX_bfv_8_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_19_0_));
    defparam IN_MUX_bfv_8_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_20_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_8_20_0_));
    defparam IN_MUX_bfv_8_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_21_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_8_21_0_));
    defparam IN_MUX_bfv_8_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_22_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_8_22_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .carryinitout(bfn_7_14_0_));
    ICE_GB delay_tr_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__18359),
            .GLOBALBUFFEROUTPUT(delay_tr_input_c_g));
    ICE_GB delay_hc_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__18335),
            .GLOBALBUFFEROUTPUT(delay_hc_input_c_g));
    ICE_GB \current_shift_inst.timer_s1.running_RNII51H_0  (
            .USERSIGNALTOGLOBALBUFFER(N__32600),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_162_i_g ));
    ICE_GB \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_0  (
            .USERSIGNALTOGLOBALBUFFER(N__36125),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst2.stoper_tr.un1_start_g ));
    ICE_GB \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_0  (
            .USERSIGNALTOGLOBALBUFFER(N__26204),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst2.stoper_hc.un1_start_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__37792),
            .CLKHFEN(N__37794),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__37793),
            .RGB2PWM(N__19346),
            .RGB1(rgb_g),
            .CURREN(N__37913),
            .RGB2(rgb_b),
            .RGB1PWM(N__18845),
            .RGB0PWM(N__48311),
            .RGB0(rgb_r));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_10_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(N__18443),
            .in2(_gnd_net_),
            .in3(N__18665),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_11_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__18431),
            .in2(N__18419),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_16 ),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__18407),
            .in2(N__18395),
            .in3(N__18386),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__18383),
            .in2(N__18371),
            .in3(N__18362),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__18572),
            .in2(N__18560),
            .in3(N__18551),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__18548),
            .in2(N__18654),
            .in3(N__18536),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(N__18533),
            .in2(N__18656),
            .in3(N__18521),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_11_6  (
            .in0(_gnd_net_),
            .in1(N__18518),
            .in2(N__18655),
            .in3(N__18506),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(N__18503),
            .in2(N__18657),
            .in3(N__18491),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__18488),
            .in2(N__18658),
            .in3(N__18476),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_24 ),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(N__18473),
            .in2(N__18662),
            .in3(N__18461),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_12_2  (
            .in0(_gnd_net_),
            .in1(N__18458),
            .in2(N__18659),
            .in3(N__18446),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_12_3  (
            .in0(_gnd_net_),
            .in1(N__18722),
            .in2(N__18663),
            .in3(N__18710),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_12_4  (
            .in0(_gnd_net_),
            .in1(N__18707),
            .in2(N__18660),
            .in3(N__18695),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_12_5  (
            .in0(_gnd_net_),
            .in1(N__18692),
            .in2(N__18664),
            .in3(N__18680),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_12_6  (
            .in0(_gnd_net_),
            .in1(N__18677),
            .in2(N__18661),
            .in3(N__18578),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18575),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_hc_LC_2_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_2_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_hc_LC_2_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29142),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18836),
            .ce(),
            .sr(N__48255));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_2_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_2_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_2_13_6 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_2_13_6  (
            .in0(N__41042),
            .in1(N__20008),
            .in2(N__18752),
            .in3(N__19815),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48794),
            .ce(),
            .sr(N__48261));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_2_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_2_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_2_14_2 .LUT_INIT=16'b0101101001001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_2_14_2  (
            .in0(N__39835),
            .in1(N__20009),
            .in2(N__18824),
            .in3(N__19830),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48785),
            .ce(),
            .sr(N__48264));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_2_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_2_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_2_15_2 .LUT_INIT=16'b1011000010110001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_2_15_2  (
            .in0(N__20001),
            .in1(N__41041),
            .in2(N__18926),
            .in3(N__19802),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48773),
            .ce(),
            .sr(N__48268));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_2_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_2_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_2_15_6 .LUT_INIT=16'b1111111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_2_15_6  (
            .in0(N__20000),
            .in1(N__41040),
            .in2(N__19829),
            .in3(N__19040),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48773),
            .ce(),
            .sr(N__48268));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_2_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_2_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_2_17_3 .LUT_INIT=16'b1111010011100100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_2_17_3  (
            .in0(N__19998),
            .in1(N__41046),
            .in2(N__19235),
            .in3(N__19814),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48755),
            .ce(),
            .sr(N__48277));
    defparam rgb_drv_RNO_LC_2_30_3.C_ON=1'b0;
    defparam rgb_drv_RNO_LC_2_30_3.SEQ_MODE=4'b0000;
    defparam rgb_drv_RNO_LC_2_30_3.LUT_INIT=16'b0000000010101010;
    LogicCell40 rgb_drv_RNO_LC_2_30_3 (
            .in0(N__43025),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48310),
            .lcout(rgb_drv_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_hc_LC_3_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_3_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_hc_LC_3_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_3_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29143),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18835),
            .ce(),
            .sr(N__48247));
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_3_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_3_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_3_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_3_13_0  (
            .in0(_gnd_net_),
            .in1(N__18820),
            .in2(N__39857),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_3_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_3_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_3_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_3_13_1  (
            .in0(_gnd_net_),
            .in1(N__39786),
            .in2(N__18803),
            .in3(N__18788),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_3_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_3_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_3_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_3_13_2  (
            .in0(_gnd_net_),
            .in1(N__39729),
            .in2(N__18785),
            .in3(N__18770),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_3_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_3_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_3_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_3_13_3  (
            .in0(_gnd_net_),
            .in1(N__39666),
            .in2(N__18767),
            .in3(N__18743),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_3_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_3_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_3_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_3_13_4  (
            .in0(_gnd_net_),
            .in1(N__39638),
            .in2(N__18740),
            .in3(N__18725),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_3_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_3_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_3_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_3_13_5  (
            .in0(_gnd_net_),
            .in1(N__39557),
            .in2(N__18995),
            .in3(N__18980),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_3_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_3_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_3_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_3_13_6  (
            .in0(_gnd_net_),
            .in1(N__39512),
            .in2(N__18977),
            .in3(N__18962),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_3_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_3_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_3_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_3_13_7  (
            .in0(_gnd_net_),
            .in1(N__39458),
            .in2(N__18959),
            .in3(N__18944),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_3_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_3_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_3_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_3_14_0  (
            .in0(_gnd_net_),
            .in1(N__40302),
            .in2(N__18941),
            .in3(N__18917),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_3_14_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_3_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_3_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_3_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_3_14_1  (
            .in0(_gnd_net_),
            .in1(N__40254),
            .in2(N__18914),
            .in3(N__18899),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_3_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_3_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_3_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_3_14_2  (
            .in0(_gnd_net_),
            .in1(N__40181),
            .in2(N__18896),
            .in3(N__18881),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_3_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_3_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_3_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_3_14_3  (
            .in0(_gnd_net_),
            .in1(N__18878),
            .in2(N__40118),
            .in3(N__18866),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_3_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_3_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_3_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_3_14_4  (
            .in0(_gnd_net_),
            .in1(N__40067),
            .in2(N__18863),
            .in3(N__18848),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_3_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_3_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_3_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_3_14_5  (
            .in0(_gnd_net_),
            .in1(N__40021),
            .in2(N__19169),
            .in3(N__19154),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_3_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_3_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_3_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_3_14_6  (
            .in0(_gnd_net_),
            .in1(N__39965),
            .in2(N__19151),
            .in3(N__19136),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_3_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_3_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_3_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_3_14_7  (
            .in0(_gnd_net_),
            .in1(N__39920),
            .in2(N__19133),
            .in3(N__19118),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_3_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_3_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_3_15_0  (
            .in0(_gnd_net_),
            .in1(N__40709),
            .in2(N__19115),
            .in3(N__19097),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_3_15_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_3_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_3_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_3_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_3_15_1  (
            .in0(_gnd_net_),
            .in1(N__40665),
            .in2(N__19094),
            .in3(N__19079),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_3_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_3_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_3_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_3_15_2  (
            .in0(_gnd_net_),
            .in1(N__40604),
            .in2(N__19076),
            .in3(N__19058),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_3_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_3_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_3_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_3_15_3  (
            .in0(_gnd_net_),
            .in1(N__40550),
            .in2(N__19055),
            .in3(N__19034),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_3_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_3_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_3_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_3_15_4  (
            .in0(_gnd_net_),
            .in1(N__40514),
            .in2(N__19031),
            .in3(N__19016),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_3_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_3_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_3_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_3_15_5  (
            .in0(_gnd_net_),
            .in1(N__40469),
            .in2(N__19013),
            .in3(N__18998),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_3_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_3_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_3_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_3_15_6  (
            .in0(_gnd_net_),
            .in1(N__40412),
            .in2(N__19325),
            .in3(N__19310),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_3_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_3_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_3_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_3_15_7  (
            .in0(_gnd_net_),
            .in1(N__19307),
            .in2(N__40379),
            .in3(N__19295),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_3_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_3_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_3_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_3_16_0  (
            .in0(_gnd_net_),
            .in1(N__41297),
            .in2(N__19292),
            .in3(N__19274),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(bfn_3_16_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_3_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_3_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_3_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_3_16_1  (
            .in0(_gnd_net_),
            .in1(N__41258),
            .in2(N__19271),
            .in3(N__19256),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_3_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_3_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_3_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_3_16_2  (
            .in0(_gnd_net_),
            .in1(N__41211),
            .in2(N__19253),
            .in3(N__19226),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_3_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_3_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_3_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_3_16_3  (
            .in0(_gnd_net_),
            .in1(N__41169),
            .in2(N__19223),
            .in3(N__19205),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_3_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_3_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_3_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_3_16_4  (
            .in0(_gnd_net_),
            .in1(N__41120),
            .in2(N__19202),
            .in3(N__19187),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_3_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_3_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_3_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_3_16_5  (
            .in0(_gnd_net_),
            .in1(N__19184),
            .in2(N__41088),
            .in3(N__19172),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_3_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_3_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_3_16_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_3_16_6  (
            .in0(N__40971),
            .in1(N__19406),
            .in2(N__19391),
            .in3(N__19376),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_3_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_3_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_3_17_1 .LUT_INIT=16'b1111111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_3_17_1  (
            .in0(N__41008),
            .in1(N__19927),
            .in2(N__19806),
            .in3(N__19373),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48742),
            .ce(),
            .sr(N__48273));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_3_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_3_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_3_17_4 .LUT_INIT=16'b1111010011100100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_3_17_4  (
            .in0(N__19926),
            .in1(N__41010),
            .in2(N__19367),
            .in3(N__19748),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48742),
            .ce(),
            .sr(N__48273));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_3_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_3_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_3_17_6 .LUT_INIT=16'b1111010011100100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_3_17_6  (
            .in0(N__19925),
            .in1(N__41009),
            .in2(N__19358),
            .in3(N__19747),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48742),
            .ce(),
            .sr(N__48273));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_3_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_3_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_3_18_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_3_18_5  (
            .in0(N__41304),
            .in1(N__41207),
            .in2(N__41270),
            .in3(N__41168),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_3_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_3_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_3_19_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_3_19_5  (
            .in0(N__40614),
            .in1(N__40661),
            .in2(N__40725),
            .in3(N__40477),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_drv_RNO_0_LC_3_30_7.C_ON=1'b0;
    defparam rgb_drv_RNO_0_LC_3_30_7.SEQ_MODE=4'b0000;
    defparam rgb_drv_RNO_0_LC_3_30_7.LUT_INIT=16'b1010101001010101;
    LogicCell40 rgb_drv_RNO_0_LC_3_30_7 (
            .in0(N__48309),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43024),
            .lcout(N_38_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_4_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_4_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_4_13_1 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_4_13_1  (
            .in0(N__19981),
            .in1(N__19823),
            .in2(_gnd_net_),
            .in3(N__19337),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48774),
            .ce(),
            .sr(N__48248));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_4_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_4_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_4_13_2 .LUT_INIT=16'b1010100010101000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_4_13_2  (
            .in0(N__19331),
            .in1(N__19980),
            .in2(N__19832),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48774),
            .ce(),
            .sr(N__48248));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_4_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_4_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_4_13_5 .LUT_INIT=16'b1010111100000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_4_13_5  (
            .in0(N__19982),
            .in1(N__19824),
            .in2(N__41050),
            .in3(N__19466),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48774),
            .ce(),
            .sr(N__48248));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_4_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_4_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_4_14_1 .LUT_INIT=16'b1011101100000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_4_14_1  (
            .in0(N__19978),
            .in1(N__41033),
            .in2(N__19821),
            .in3(N__19460),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48765),
            .ce(),
            .sr(N__48256));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_4_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_4_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_4_14_3 .LUT_INIT=16'b1111111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_4_14_3  (
            .in0(N__19977),
            .in1(N__41032),
            .in2(N__19820),
            .in3(N__19454),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48765),
            .ce(),
            .sr(N__48256));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_4_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_4_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_4_14_5 .LUT_INIT=16'b1011101100000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_4_14_5  (
            .in0(N__19979),
            .in1(N__41034),
            .in2(N__19822),
            .in3(N__19448),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48765),
            .ce(),
            .sr(N__48256));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_4_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_4_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_4_14_6 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_4_14_6  (
            .in0(N__41031),
            .in1(N__19976),
            .in2(N__19442),
            .in3(N__19788),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48765),
            .ce(),
            .sr(N__48256));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_4_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_4_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_4_15_0 .LUT_INIT=16'b1111111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_4_15_0  (
            .in0(N__19965),
            .in1(N__41004),
            .in2(N__19817),
            .in3(N__19433),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48756),
            .ce(),
            .sr(N__48262));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_4_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_4_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_4_15_1 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_4_15_1  (
            .in0(N__41002),
            .in1(N__19968),
            .in2(N__19427),
            .in3(N__19778),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48756),
            .ce(),
            .sr(N__48262));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_4_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_4_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_4_15_2 .LUT_INIT=16'b1111111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_4_15_2  (
            .in0(N__19967),
            .in1(N__41005),
            .in2(N__19818),
            .in3(N__19418),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48756),
            .ce(),
            .sr(N__48262));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_4_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_4_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_4_15_4 .LUT_INIT=16'b1111111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_4_15_4  (
            .in0(N__19969),
            .in1(N__41006),
            .in2(N__19819),
            .in3(N__19412),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48756),
            .ce(),
            .sr(N__48262));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_4_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_4_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_4_15_5 .LUT_INIT=16'b1111000011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_4_15_5  (
            .in0(N__41000),
            .in1(N__19776),
            .in2(N__19538),
            .in3(N__19963),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48756),
            .ce(),
            .sr(N__48262));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_4_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_4_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_4_15_6 .LUT_INIT=16'b1111111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_4_15_6  (
            .in0(N__19964),
            .in1(N__41003),
            .in2(N__19816),
            .in3(N__19529),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48756),
            .ce(),
            .sr(N__48262));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_4_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_4_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_4_15_7 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_4_15_7  (
            .in0(N__41001),
            .in1(N__19966),
            .in2(N__19523),
            .in3(N__19777),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48756),
            .ce(),
            .sr(N__48262));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_4_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_4_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_4_16_0 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_4_16_0  (
            .in0(N__40995),
            .in1(N__19958),
            .in2(N__19514),
            .in3(N__19739),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48743),
            .ce(),
            .sr(N__48265));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_4_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_4_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_4_16_2 .LUT_INIT=16'b1111000011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_4_16_2  (
            .in0(N__40997),
            .in1(N__19740),
            .in2(N__19502),
            .in3(N__19961),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48743),
            .ce(),
            .sr(N__48265));
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_4_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_4_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_4_16_3 .LUT_INIT=16'b1111111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_31_LC_4_16_3  (
            .in0(N__19962),
            .in1(N__40998),
            .in2(N__19804),
            .in3(N__19493),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48743),
            .ce(),
            .sr(N__48265));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_4_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_4_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_4_16_5 .LUT_INIT=16'b1101110111001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_4_16_5  (
            .in0(N__19960),
            .in1(N__19487),
            .in2(N__19803),
            .in3(N__40999),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48743),
            .ce(),
            .sr(N__48265));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_4_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_4_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_4_16_6 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_4_16_6  (
            .in0(N__40996),
            .in1(N__19959),
            .in2(N__19481),
            .in3(N__19738),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48743),
            .ce(),
            .sr(N__48265));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_4_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_4_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_4_17_5 .LUT_INIT=16'b1111111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_4_17_5  (
            .in0(N__19895),
            .in1(N__41011),
            .in2(N__19807),
            .in3(N__19472),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48732),
            .ce(),
            .sr(N__48269));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_4_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_4_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_4_18_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_4_18_1  (
            .in0(N__39966),
            .in1(N__40250),
            .in2(N__40081),
            .in3(N__39925),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_4_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_4_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_4_18_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_4_18_2  (
            .in0(N__40194),
            .in1(N__40020),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_4_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_4_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_4_18_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_4_18_3  (
            .in0(N__40129),
            .in1(N__19574),
            .in2(N__19568),
            .in3(N__41078),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_4_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_4_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_4_18_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_4_18_4  (
            .in0(N__20099),
            .in1(N__19565),
            .in2(N__19559),
            .in3(N__19544),
            .lcout(\current_shift_inst.PI_CTRL.N_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_4_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_4_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_4_19_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_4_19_0  (
            .in0(N__39519),
            .in1(N__39472),
            .in2(N__39581),
            .in3(N__40323),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_4_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_4_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_4_19_1 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_4_19_1  (
            .in0(N__39645),
            .in1(N__39690),
            .in2(N__19556),
            .in3(N__39748),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_44_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_4_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_4_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_4_19_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_4_19_2  (
            .in0(N__41136),
            .in1(N__40413),
            .in2(N__19553),
            .in3(N__19550),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_4_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_4_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_4_21_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_4_21_3  (
            .in0(N__39921),
            .in1(N__40016),
            .in2(N__40198),
            .in3(N__40128),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_4_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_4_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_4_22_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_4_22_0  (
            .in0(_gnd_net_),
            .in1(N__41259),
            .in2(_gnd_net_),
            .in3(N__40515),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_4_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_4_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_4_22_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_4_22_2  (
            .in0(N__41179),
            .in1(N__41224),
            .in2(N__41314),
            .in3(N__41092),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_4_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_4_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_4_22_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_4_22_3  (
            .in0(N__40560),
            .in1(N__40383),
            .in2(N__19616),
            .in3(N__19613),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_4_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_4_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_4_22_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_4_22_5  (
            .in0(N__40615),
            .in1(N__40669),
            .in2(N__40735),
            .in3(N__40473),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_4_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_4_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_4_22_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_4_22_6  (
            .in0(N__41013),
            .in1(N__40420),
            .in2(N__19607),
            .in3(N__19604),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_4_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_4_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_4_22_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_4_22_7  (
            .in0(N__20093),
            .in1(N__19598),
            .in2(N__19592),
            .in3(N__19580),
            .lcout(\current_shift_inst.PI_CTRL.N_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_4_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_4_23_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_4_23_4 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_4_23_4  (
            .in0(N__39523),
            .in1(N__39647),
            .in2(_gnd_net_),
            .in3(N__39471),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_4_23_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_4_23_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_4_23_5 .LUT_INIT=16'b0000000000110111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_4_23_5  (
            .in0(N__39796),
            .in1(N__39747),
            .in2(N__39877),
            .in3(N__39694),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_77_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_4_23_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_4_23_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_4_23_6 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_4_23_6  (
            .in0(N__19589),
            .in1(N__40327),
            .in2(N__19583),
            .in3(N__39573),
            .lcout(\current_shift_inst.PI_CTRL.N_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_5_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_5_7_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_5_7_1  (
            .in0(N__23611),
            .in1(N__23589),
            .in2(_gnd_net_),
            .in3(N__41887),
            .lcout(elapsed_time_ns_1_RNI7ADN9_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_5_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_5_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_5_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_29_LC_5_8_7  (
            .in0(N__23610),
            .in1(N__23590),
            .in2(_gnd_net_),
            .in3(N__41816),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48804),
            .ce(N__28504),
            .sr(N__48215));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_5_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_5_9_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_5_9_3  (
            .in0(N__41884),
            .in1(N__23670),
            .in2(_gnd_net_),
            .in3(N__23650),
            .lcout(elapsed_time_ns_1_RNIL73T9_0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_5_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_5_10_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_5_10_0  (
            .in0(N__28283),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28209),
            .lcout(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_5_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_5_10_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_5_10_2  (
            .in0(N__23883),
            .in1(N__23864),
            .in2(_gnd_net_),
            .in3(N__41881),
            .lcout(elapsed_time_ns_1_RNIDV2T9_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_5_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_5_10_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_5_10_4  (
            .in0(N__20055),
            .in1(N__20431),
            .in2(_gnd_net_),
            .in3(N__41883),
            .lcout(elapsed_time_ns_1_RNIUVBN9_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_5_10_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_5_10_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_5_10_6  (
            .in0(N__31533),
            .in1(N__31503),
            .in2(_gnd_net_),
            .in3(N__41882),
            .lcout(elapsed_time_ns_1_RNI03DN9_0_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_5_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_5_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_5_12_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_22_LC_5_12_1  (
            .in0(N__41886),
            .in1(N__31534),
            .in2(_gnd_net_),
            .in3(N__31510),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48775),
            .ce(N__28502),
            .sr(N__48237));
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_5_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_5_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_5_12_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_11_LC_5_12_5  (
            .in0(N__41885),
            .in1(N__20056),
            .in2(_gnd_net_),
            .in3(N__20430),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48775),
            .ce(N__28502),
            .sr(N__48237));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_5_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_5_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_5_13_6 .LUT_INIT=16'b1101000011010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_5_13_6  (
            .in0(N__41036),
            .in1(N__19999),
            .in2(N__20033),
            .in3(N__19828),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48766),
            .ce(),
            .sr(N__48242));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_5_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_5_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_5_14_2 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_5_14_2  (
            .in0(N__41035),
            .in1(N__19997),
            .in2(N__20021),
            .in3(N__19831),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48757),
            .ce(),
            .sr(N__48249));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_5_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_5_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_5_15_4 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_5_15_4  (
            .in0(N__41007),
            .in1(N__19983),
            .in2(N__19847),
            .in3(N__19805),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48744),
            .ce(),
            .sr(N__48257));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_5_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_5_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_5_19_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_5_19_5  (
            .in0(N__40384),
            .in1(N__40573),
            .in2(N__40529),
            .in3(N__41012),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_5_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_5_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_5_22_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_5_22_1  (
            .in0(N__39979),
            .in1(N__40080),
            .in2(N__40261),
            .in3(N__41140),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_5_30_0.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_5_30_0.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_5_30_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_5_30_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20087),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_7_5_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_7_5_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_7_5_1  (
            .in0(N__22971),
            .in1(N__24058),
            .in2(_gnd_net_),
            .in3(N__41878),
            .lcout(elapsed_time_ns_1_RNI68CN9_0_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_7_6_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_7_6_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_7_6_0  (
            .in0(N__23938),
            .in1(N__23379),
            .in2(_gnd_net_),
            .in3(N__41898),
            .lcout(elapsed_time_ns_1_RNI04EN9_0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_7_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_7_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_7_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_19_LC_7_7_7  (
            .in0(N__22972),
            .in1(N__24062),
            .in2(_gnd_net_),
            .in3(N__41899),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48799),
            .ce(N__28508),
            .sr(N__48191));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_7_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_7_8_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_7_8_4  (
            .in0(N__23736),
            .in1(N__23713),
            .in2(_gnd_net_),
            .in3(N__41814),
            .lcout(elapsed_time_ns_1_RNITUBN9_0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_7_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_7_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_7_8_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_11_LC_7_8_7  (
            .in0(N__41815),
            .in1(N__20060),
            .in2(_gnd_net_),
            .in3(N__20432),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48795),
            .ce(N__36595),
            .sr(N__48201));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_7_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_7_9_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_7_9_2  (
            .in0(N__31612),
            .in1(N__31585),
            .in2(_gnd_net_),
            .in3(N__41861),
            .lcout(elapsed_time_ns_1_RNI14DN9_0_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_7_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_7_9_3 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_7_9_3  (
            .in0(N__22021),
            .in1(N__25963),
            .in2(N__25996),
            .in3(N__22000),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_7_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_7_9_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_7_9_5  (
            .in0(_gnd_net_),
            .in1(N__23239),
            .in2(_gnd_net_),
            .in3(N__25080),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_7_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_7_9_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_7_9_6  (
            .in0(N__24916),
            .in1(N__23162),
            .in2(N__20135),
            .in3(N__20132),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_7_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_7_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_7_10_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_12_LC_7_10_1  (
            .in0(N__28706),
            .in1(N__28744),
            .in2(_gnd_net_),
            .in3(N__41903),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48776),
            .ce(N__36444),
            .sr(N__48216));
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_7_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_7_10_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.state_RNIG7JF_2_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(N__31768),
            .in2(_gnd_net_),
            .in3(N__31801),
            .lcout(\phase_controller_inst2.state_RNIG7JFZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_7_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_7_11_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_7_11_4  (
            .in0(N__20414),
            .in1(N__23699),
            .in2(N__28739),
            .in3(N__23636),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_7_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_7_12_0 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_7_12_0  (
            .in0(N__20108),
            .in1(N__20122),
            .in2(N__25886),
            .in3(N__25859),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_7_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_7_12_1 .LUT_INIT=16'b1111011101010001;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_7_12_1  (
            .in0(N__25858),
            .in1(N__25885),
            .in2(N__20123),
            .in3(N__20107),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_7_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_7_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_7_12_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_23_LC_7_12_3  (
            .in0(N__41901),
            .in1(N__31608),
            .in2(_gnd_net_),
            .in3(N__31574),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48758),
            .ce(N__28503),
            .sr(N__48227));
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_7_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_7_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_7_12_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_9_LC_7_12_4  (
            .in0(N__23643),
            .in1(N__23678),
            .in2(_gnd_net_),
            .in3(N__41902),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48758),
            .ce(N__28503),
            .sr(N__48227));
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_7_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_7_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_7_12_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_10_LC_7_12_5  (
            .in0(N__41900),
            .in1(N__23737),
            .in2(_gnd_net_),
            .in3(N__23703),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48758),
            .ce(N__28503),
            .sr(N__48227));
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_7_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_7_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__20162),
            .in2(_gnd_net_),
            .in3(N__22487),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_7_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_7_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_7_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_1_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(N__22475),
            .in2(_gnd_net_),
            .in3(N__20156),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .clk(N__48745),
            .ce(),
            .sr(N__48232));
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_7_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_7_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_7_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(N__22454),
            .in2(_gnd_net_),
            .in3(N__20153),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .clk(N__48745),
            .ce(),
            .sr(N__48232));
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_7_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_7_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_7_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_3_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(N__22439),
            .in2(_gnd_net_),
            .in3(N__20150),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .clk(N__48745),
            .ce(),
            .sr(N__48232));
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_7_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_7_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_7_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_4_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(N__22418),
            .in2(_gnd_net_),
            .in3(N__20147),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .clk(N__48745),
            .ce(),
            .sr(N__48232));
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_7_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_7_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_7_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_5_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(N__22397),
            .in2(_gnd_net_),
            .in3(N__20144),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .clk(N__48745),
            .ce(),
            .sr(N__48232));
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_7_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_7_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_7_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_6_LC_7_13_6  (
            .in0(_gnd_net_),
            .in1(N__22376),
            .in2(_gnd_net_),
            .in3(N__20141),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .clk(N__48745),
            .ce(),
            .sr(N__48232));
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_7_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_7_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_7_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_7_LC_7_13_7  (
            .in0(_gnd_net_),
            .in1(N__22616),
            .in2(_gnd_net_),
            .in3(N__20138),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .clk(N__48745),
            .ce(),
            .sr(N__48232));
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_7_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_7_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_7_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_8_LC_7_14_0  (
            .in0(_gnd_net_),
            .in1(N__22601),
            .in2(_gnd_net_),
            .in3(N__20183),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_8 ),
            .ltout(),
            .carryin(bfn_7_14_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .clk(N__48733),
            .ce(),
            .sr(N__48238));
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_7_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_7_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_7_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_9_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(N__22586),
            .in2(_gnd_net_),
            .in3(N__20180),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .clk(N__48733),
            .ce(),
            .sr(N__48238));
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_7_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_7_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_7_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_10_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(N__22571),
            .in2(_gnd_net_),
            .in3(N__20177),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .clk(N__48733),
            .ce(),
            .sr(N__48238));
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_7_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_7_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_7_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_11_LC_7_14_3  (
            .in0(_gnd_net_),
            .in1(N__22556),
            .in2(_gnd_net_),
            .in3(N__20174),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .clk(N__48733),
            .ce(),
            .sr(N__48238));
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_7_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_7_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_7_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_12_LC_7_14_4  (
            .in0(_gnd_net_),
            .in1(N__22535),
            .in2(_gnd_net_),
            .in3(N__20171),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .clk(N__48733),
            .ce(),
            .sr(N__48238));
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_7_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_7_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_7_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_13_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(N__21059),
            .in2(_gnd_net_),
            .in3(N__20168),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .clk(N__48733),
            .ce(),
            .sr(N__48238));
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_7_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_7_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_7_14_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_14_LC_7_14_6  (
            .in0(_gnd_net_),
            .in1(N__22517),
            .in2(_gnd_net_),
            .in3(N__20165),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48733),
            .ce(),
            .sr(N__48238));
    defparam \phase_controller_inst2.state_1_LC_7_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_1_LC_7_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_1_LC_7_14_7 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \phase_controller_inst2.state_1_LC_7_14_7  (
            .in0(N__27793),
            .in1(N__31830),
            .in2(_gnd_net_),
            .in3(N__31715),
            .lcout(\phase_controller_inst2.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48733),
            .ce(),
            .sr(N__48238));
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_7_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_7_17_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_7_17_0  (
            .in0(N__26911),
            .in1(N__32143),
            .in2(_gnd_net_),
            .in3(N__32112),
            .lcout(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_7_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_7_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_7_17_4 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_7_17_4  (
            .in0(N__26910),
            .in1(N__33695),
            .in2(_gnd_net_),
            .in3(N__33649),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_7_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_7_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32400),
            .lcout(\current_shift_inst.un4_control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_7_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_7_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24231),
            .lcout(\current_shift_inst.un4_control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_7_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_7_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_7_19_2 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_7_19_2  (
            .in0(_gnd_net_),
            .in1(N__29784),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_7_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_7_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_7_19_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(N__32652),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_7_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_7_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_7_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_7_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29600),
            .lcout(\current_shift_inst.un4_control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_7_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_7_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_7_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24421),
            .lcout(\current_shift_inst.un4_control_input_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_7_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_7_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_7_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_7_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29519),
            .lcout(\current_shift_inst.un4_control_input_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_7_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_7_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_7_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_7_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32318),
            .lcout(\current_shift_inst.un4_control_input_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_7_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_7_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_7_20_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_7_20_0  (
            .in0(_gnd_net_),
            .in1(N__21255),
            .in2(N__21232),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_7_20_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__48684),
            .ce(N__33740),
            .sr(N__48270));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_7_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_7_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_7_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_7_20_1  (
            .in0(_gnd_net_),
            .in1(N__23955),
            .in2(N__21208),
            .in3(N__20210),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__48684),
            .ce(N__33740),
            .sr(N__48270));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_7_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_7_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_7_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_7_20_2  (
            .in0(_gnd_net_),
            .in1(N__21447),
            .in2(N__21233),
            .in3(N__20207),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__48684),
            .ce(N__33740),
            .sr(N__48270));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_7_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_7_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_7_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_7_20_3  (
            .in0(_gnd_net_),
            .in1(N__21423),
            .in2(N__21209),
            .in3(N__20204),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__48684),
            .ce(N__33740),
            .sr(N__48270));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_7_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_7_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_7_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_7_20_4  (
            .in0(_gnd_net_),
            .in1(N__21399),
            .in2(N__21452),
            .in3(N__20201),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__48684),
            .ce(N__33740),
            .sr(N__48270));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_7_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_7_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_7_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_7_20_5  (
            .in0(_gnd_net_),
            .in1(N__21375),
            .in2(N__21428),
            .in3(N__20198),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__48684),
            .ce(N__33740),
            .sr(N__48270));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_7_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_7_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_7_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_7_20_6  (
            .in0(_gnd_net_),
            .in1(N__21351),
            .in2(N__21404),
            .in3(N__20195),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__48684),
            .ce(N__33740),
            .sr(N__48270));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_7_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_7_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_7_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_7_20_7  (
            .in0(_gnd_net_),
            .in1(N__21327),
            .in2(N__21380),
            .in3(N__20192),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__48684),
            .ce(N__33740),
            .sr(N__48270));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_7_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_7_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_7_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_7_21_0  (
            .in0(_gnd_net_),
            .in1(N__21303),
            .in2(N__21356),
            .in3(N__20189),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_7_21_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__48679),
            .ce(N__33739),
            .sr(N__48274));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_7_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_7_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_7_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_7_21_1  (
            .in0(_gnd_net_),
            .in1(N__21279),
            .in2(N__21332),
            .in3(N__20186),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__48679),
            .ce(N__33739),
            .sr(N__48274));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_7_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_7_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_7_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_7_21_2  (
            .in0(_gnd_net_),
            .in1(N__21660),
            .in2(N__21308),
            .in3(N__20237),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__48679),
            .ce(N__33739),
            .sr(N__48274));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_7_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_7_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_7_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_7_21_3  (
            .in0(_gnd_net_),
            .in1(N__21636),
            .in2(N__21284),
            .in3(N__20234),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__48679),
            .ce(N__33739),
            .sr(N__48274));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_7_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_7_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_7_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_7_21_4  (
            .in0(_gnd_net_),
            .in1(N__21612),
            .in2(N__21665),
            .in3(N__20231),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__48679),
            .ce(N__33739),
            .sr(N__48274));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_7_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_7_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_7_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_7_21_5  (
            .in0(_gnd_net_),
            .in1(N__21588),
            .in2(N__21641),
            .in3(N__20228),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__48679),
            .ce(N__33739),
            .sr(N__48274));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_7_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_7_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_7_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_7_21_6  (
            .in0(_gnd_net_),
            .in1(N__21564),
            .in2(N__21617),
            .in3(N__20225),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__48679),
            .ce(N__33739),
            .sr(N__48274));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_7_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_7_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_7_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_7_21_7  (
            .in0(_gnd_net_),
            .in1(N__21540),
            .in2(N__21593),
            .in3(N__20222),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__48679),
            .ce(N__33739),
            .sr(N__48274));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_7_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_7_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_7_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_7_22_0  (
            .in0(_gnd_net_),
            .in1(N__21516),
            .in2(N__21569),
            .in3(N__20219),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_7_22_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__48675),
            .ce(N__33738),
            .sr(N__48278));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_7_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_7_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_7_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_7_22_1  (
            .in0(_gnd_net_),
            .in1(N__21492),
            .in2(N__21545),
            .in3(N__20216),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__48675),
            .ce(N__33738),
            .sr(N__48278));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_7_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_7_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_7_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_7_22_2  (
            .in0(_gnd_net_),
            .in1(N__21468),
            .in2(N__21521),
            .in3(N__20213),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__48675),
            .ce(N__33738),
            .sr(N__48278));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_7_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_7_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_7_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_7_22_3  (
            .in0(_gnd_net_),
            .in1(N__21843),
            .in2(N__21497),
            .in3(N__20264),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__48675),
            .ce(N__33738),
            .sr(N__48278));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_7_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_7_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_7_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_7_22_4  (
            .in0(_gnd_net_),
            .in1(N__21819),
            .in2(N__21473),
            .in3(N__20261),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__48675),
            .ce(N__33738),
            .sr(N__48278));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_7_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_7_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_7_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_7_22_5  (
            .in0(_gnd_net_),
            .in1(N__21795),
            .in2(N__21848),
            .in3(N__20258),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__48675),
            .ce(N__33738),
            .sr(N__48278));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_7_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_7_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_7_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_7_22_6  (
            .in0(_gnd_net_),
            .in1(N__21771),
            .in2(N__21824),
            .in3(N__20255),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__48675),
            .ce(N__33738),
            .sr(N__48278));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_7_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_7_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_7_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_7_22_7  (
            .in0(_gnd_net_),
            .in1(N__21747),
            .in2(N__21800),
            .in3(N__20252),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__48675),
            .ce(N__33738),
            .sr(N__48278));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_7_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_7_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_7_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_7_23_0  (
            .in0(_gnd_net_),
            .in1(N__21723),
            .in2(N__21776),
            .in3(N__20249),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_7_23_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__48669),
            .ce(N__33737),
            .sr(N__48281));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_7_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_7_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_7_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_7_23_1  (
            .in0(_gnd_net_),
            .in1(N__21699),
            .in2(N__21752),
            .in3(N__20246),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__48669),
            .ce(N__33737),
            .sr(N__48281));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_7_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_7_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_7_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_7_23_2  (
            .in0(_gnd_net_),
            .in1(N__21679),
            .in2(N__21728),
            .in3(N__20243),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__48669),
            .ce(N__33737),
            .sr(N__48281));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_7_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_7_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_7_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_7_23_3  (
            .in0(_gnd_net_),
            .in1(N__21904),
            .in2(N__21704),
            .in3(N__20240),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__48669),
            .ce(N__33737),
            .sr(N__48281));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_7_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_7_23_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_7_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_7_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20312),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_7_24_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_7_24_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_7_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_7_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20308),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48665),
            .ce(),
            .sr(N__48282));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_8_3_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_8_3_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_8_3_4  (
            .in0(N__21869),
            .in1(N__23292),
            .in2(_gnd_net_),
            .in3(N__41890),
            .lcout(elapsed_time_ns_1_RNI24CN9_0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_5_1.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_5_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_5_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH1_MAX_D1_LC_8_5_1 (
            .in0(N__20282),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_max_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48805),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_8_5_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_8_5_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_8_5_5  (
            .in0(N__22948),
            .in1(N__24023),
            .in2(_gnd_net_),
            .in3(N__41825),
            .lcout(elapsed_time_ns_1_RNI57CN9_0_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_8_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_8_6_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_8_6_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_14_LC_8_6_5  (
            .in0(N__30725),
            .in1(N__30767),
            .in2(_gnd_net_),
            .in3(N__41833),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48800),
            .ce(N__28511),
            .sr(N__48173));
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_8_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_8_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_8_6_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_18_LC_8_6_6  (
            .in0(N__41832),
            .in1(N__22944),
            .in2(_gnd_net_),
            .in3(N__24021),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48800),
            .ce(N__28511),
            .sr(N__48173));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_8_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_8_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_8_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_8_7_0  (
            .in0(N__29116),
            .in1(N__21951),
            .in2(_gnd_net_),
            .in3(N__20273),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__48796),
            .ce(N__29219),
            .sr(N__48182));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_8_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_8_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_8_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_8_7_1  (
            .in0(N__29112),
            .in1(N__21927),
            .in2(_gnd_net_),
            .in3(N__20270),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__48796),
            .ce(N__29219),
            .sr(N__48182));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_8_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_8_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_8_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_8_7_2  (
            .in0(N__29117),
            .in1(N__20607),
            .in2(_gnd_net_),
            .in3(N__20267),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__48796),
            .ce(N__29219),
            .sr(N__48182));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_8_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_8_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_8_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_8_7_3  (
            .in0(N__29113),
            .in1(N__20581),
            .in2(_gnd_net_),
            .in3(N__20339),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__48796),
            .ce(N__29219),
            .sr(N__48182));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_8_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_8_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_8_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_8_7_4  (
            .in0(N__29118),
            .in1(N__20556),
            .in2(_gnd_net_),
            .in3(N__20336),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__48796),
            .ce(N__29219),
            .sr(N__48182));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_8_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_8_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_8_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_8_7_5  (
            .in0(N__29114),
            .in1(N__20529),
            .in2(_gnd_net_),
            .in3(N__20333),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__48796),
            .ce(N__29219),
            .sr(N__48182));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_8_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_8_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_8_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_8_7_6  (
            .in0(N__29119),
            .in1(N__20503),
            .in2(_gnd_net_),
            .in3(N__20330),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__48796),
            .ce(N__29219),
            .sr(N__48182));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_8_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_8_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_8_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_8_7_7  (
            .in0(N__29115),
            .in1(N__20479),
            .in2(_gnd_net_),
            .in3(N__20327),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__48796),
            .ce(N__29219),
            .sr(N__48182));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_8_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_8_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_8_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_8_8_0  (
            .in0(N__29111),
            .in1(N__20448),
            .in2(_gnd_net_),
            .in3(N__20324),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__48786),
            .ce(N__29218),
            .sr(N__48192));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_8_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_8_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_8_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_8_8_1  (
            .in0(N__29123),
            .in1(N__20829),
            .in2(_gnd_net_),
            .in3(N__20321),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__48786),
            .ce(N__29218),
            .sr(N__48192));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_8_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_8_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_8_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_8_8_2  (
            .in0(N__29108),
            .in1(N__20800),
            .in2(_gnd_net_),
            .in3(N__20318),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__48786),
            .ce(N__29218),
            .sr(N__48192));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_8_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_8_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_8_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_8_8_3  (
            .in0(N__29120),
            .in1(N__20781),
            .in2(_gnd_net_),
            .in3(N__20315),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__48786),
            .ce(N__29218),
            .sr(N__48192));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_8_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_8_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_8_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_8_8_4  (
            .in0(N__29109),
            .in1(N__20754),
            .in2(_gnd_net_),
            .in3(N__20366),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__48786),
            .ce(N__29218),
            .sr(N__48192));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_8_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_8_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_8_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_8_8_5  (
            .in0(N__29121),
            .in1(N__20727),
            .in2(_gnd_net_),
            .in3(N__20363),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__48786),
            .ce(N__29218),
            .sr(N__48192));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_8_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_8_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_8_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_8_8_6  (
            .in0(N__29110),
            .in1(N__20697),
            .in2(_gnd_net_),
            .in3(N__20360),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__48786),
            .ce(N__29218),
            .sr(N__48192));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_8_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_8_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_8_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_8_8_7  (
            .in0(N__29122),
            .in1(N__20667),
            .in2(_gnd_net_),
            .in3(N__20357),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__48786),
            .ce(N__29218),
            .sr(N__48192));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_8_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_8_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_8_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_8_9_0  (
            .in0(N__29100),
            .in1(N__20643),
            .in2(_gnd_net_),
            .in3(N__20354),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__48777),
            .ce(N__29217),
            .sr(N__48202));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_8_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_8_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_8_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_8_9_1  (
            .in0(N__29104),
            .in1(N__21042),
            .in2(_gnd_net_),
            .in3(N__20351),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__48777),
            .ce(N__29217),
            .sr(N__48202));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_8_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_8_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_8_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_8_9_2  (
            .in0(N__29101),
            .in1(N__21018),
            .in2(_gnd_net_),
            .in3(N__20348),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__48777),
            .ce(N__29217),
            .sr(N__48202));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_8_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_8_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_8_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_8_9_3  (
            .in0(N__29105),
            .in1(N__20994),
            .in2(_gnd_net_),
            .in3(N__20345),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__48777),
            .ce(N__29217),
            .sr(N__48202));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_8_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_8_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_8_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_8_9_4  (
            .in0(N__29102),
            .in1(N__20973),
            .in2(_gnd_net_),
            .in3(N__20342),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__48777),
            .ce(N__29217),
            .sr(N__48202));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_8_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_8_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_8_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_8_9_5  (
            .in0(N__29106),
            .in1(N__20949),
            .in2(_gnd_net_),
            .in3(N__20393),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__48777),
            .ce(N__29217),
            .sr(N__48202));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_8_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_8_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_8_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_8_9_6  (
            .in0(N__29103),
            .in1(N__20914),
            .in2(_gnd_net_),
            .in3(N__20390),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__48777),
            .ce(N__29217),
            .sr(N__48202));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_8_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_8_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_8_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_8_9_7  (
            .in0(N__29107),
            .in1(N__20889),
            .in2(_gnd_net_),
            .in3(N__20387),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__48777),
            .ce(N__29217),
            .sr(N__48202));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_8_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_8_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_8_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_8_10_0  (
            .in0(N__29058),
            .in1(N__20859),
            .in2(_gnd_net_),
            .in3(N__20384),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__48767),
            .ce(N__29210),
            .sr(N__48209));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_8_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_8_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_8_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_8_10_1  (
            .in0(N__29062),
            .in1(N__21165),
            .in2(_gnd_net_),
            .in3(N__20381),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__48767),
            .ce(N__29210),
            .sr(N__48209));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_8_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_8_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_8_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_8_10_2  (
            .in0(N__29059),
            .in1(N__21126),
            .in2(_gnd_net_),
            .in3(N__20378),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__48767),
            .ce(N__29210),
            .sr(N__48209));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_8_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_8_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_8_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_8_10_3  (
            .in0(N__29063),
            .in1(N__21084),
            .in2(_gnd_net_),
            .in3(N__20375),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__48767),
            .ce(N__29210),
            .sr(N__48209));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_8_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_8_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_8_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_8_10_4  (
            .in0(N__29060),
            .in1(N__21145),
            .in2(_gnd_net_),
            .in3(N__20372),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__48767),
            .ce(N__29210),
            .sr(N__48209));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_8_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_8_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_8_10_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_8_10_5  (
            .in0(N__21103),
            .in1(N__29061),
            .in2(_gnd_net_),
            .in3(N__20369),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48767),
            .ce(N__29210),
            .sr(N__48209));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_8_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_8_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_8_11_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(N__21956),
            .in2(N__20618),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__48759),
            .ce(N__29882),
            .sr(N__48217));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_8_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_8_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_8_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__20587),
            .in2(N__21935),
            .in3(N__20621),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__48759),
            .ce(N__29882),
            .sr(N__48217));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_8_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_8_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_8_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(N__20617),
            .in2(N__20563),
            .in3(N__20591),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__48759),
            .ce(N__29882),
            .sr(N__48217));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_8_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_8_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_8_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__20588),
            .in2(N__20536),
            .in3(N__20567),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__48759),
            .ce(N__29882),
            .sr(N__48217));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_8_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_8_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_8_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(N__20509),
            .in2(N__20564),
            .in3(N__20540),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__48759),
            .ce(N__29882),
            .sr(N__48217));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_8_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_8_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_8_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(N__20485),
            .in2(N__20537),
            .in3(N__20513),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__48759),
            .ce(N__29882),
            .sr(N__48217));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_8_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_8_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_8_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(N__20510),
            .in2(N__20461),
            .in3(N__20489),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__48759),
            .ce(N__29882),
            .sr(N__48217));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_8_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_8_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_8_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(N__20486),
            .in2(N__20836),
            .in3(N__20465),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__48759),
            .ce(N__29882),
            .sr(N__48217));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_8_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_8_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_8_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_8_12_0  (
            .in0(_gnd_net_),
            .in1(N__20806),
            .in2(N__20462),
            .in3(N__20396),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_8_12_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__48746),
            .ce(N__29887),
            .sr(N__48221));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_8_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_8_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_8_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(N__20782),
            .in2(N__20840),
            .in3(N__20810),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__48746),
            .ce(N__29887),
            .sr(N__48221));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_8_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_8_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_8_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(N__20807),
            .in2(N__20761),
            .in3(N__20786),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__48746),
            .ce(N__29887),
            .sr(N__48221));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_8_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_8_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_8_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(N__20783),
            .in2(N__20734),
            .in3(N__20765),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__48746),
            .ce(N__29887),
            .sr(N__48221));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_8_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_8_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_8_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_8_12_4  (
            .in0(_gnd_net_),
            .in1(N__20704),
            .in2(N__20762),
            .in3(N__20738),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__48746),
            .ce(N__29887),
            .sr(N__48221));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_8_12_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_8_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_8_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_8_12_5  (
            .in0(_gnd_net_),
            .in1(N__20674),
            .in2(N__20735),
            .in3(N__20711),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__48746),
            .ce(N__29887),
            .sr(N__48221));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_8_12_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_8_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_8_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_8_12_6  (
            .in0(_gnd_net_),
            .in1(N__20644),
            .in2(N__20708),
            .in3(N__20681),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__48746),
            .ce(N__29887),
            .sr(N__48221));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_8_12_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_8_12_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_8_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_8_12_7  (
            .in0(_gnd_net_),
            .in1(N__21049),
            .in2(N__20678),
            .in3(N__20651),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__48746),
            .ce(N__29887),
            .sr(N__48221));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_8_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_8_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_8_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(N__21019),
            .in2(N__20648),
            .in3(N__20624),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__48734),
            .ce(N__29886),
            .sr(N__48228));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_8_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_8_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_8_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__20995),
            .in2(N__21053),
            .in3(N__21026),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__48734),
            .ce(N__29886),
            .sr(N__48228));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_8_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_8_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_8_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__20974),
            .in2(N__21023),
            .in3(N__20999),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__48734),
            .ce(N__29886),
            .sr(N__48228));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_8_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_8_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_8_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(N__20996),
            .in2(N__20954),
            .in3(N__20978),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__48734),
            .ce(N__29886),
            .sr(N__48228));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_8_13_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_8_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_8_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__20975),
            .in2(N__20926),
            .in3(N__20957),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__48734),
            .ce(N__29886),
            .sr(N__48228));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_8_13_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_8_13_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_8_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_8_13_5  (
            .in0(_gnd_net_),
            .in1(N__20953),
            .in2(N__20896),
            .in3(N__20930),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__48734),
            .ce(N__29886),
            .sr(N__48228));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_8_13_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_8_13_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_8_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_8_13_6  (
            .in0(_gnd_net_),
            .in1(N__20866),
            .in2(N__20927),
            .in3(N__20900),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__48734),
            .ce(N__29886),
            .sr(N__48228));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_8_13_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_8_13_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_8_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_8_13_7  (
            .in0(_gnd_net_),
            .in1(N__21172),
            .in2(N__20897),
            .in3(N__20873),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__48734),
            .ce(N__29886),
            .sr(N__48228));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_8_14_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_8_14_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_8_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_8_14_0  (
            .in0(_gnd_net_),
            .in1(N__21127),
            .in2(N__20870),
            .in3(N__20843),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__48724),
            .ce(N__29875),
            .sr(N__48233));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_8_14_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_8_14_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_8_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_8_14_1  (
            .in0(_gnd_net_),
            .in1(N__21085),
            .in2(N__21176),
            .in3(N__21149),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__48724),
            .ce(N__29875),
            .sr(N__48233));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_8_14_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_8_14_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_8_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_8_14_2  (
            .in0(_gnd_net_),
            .in1(N__21146),
            .in2(N__21131),
            .in3(N__21107),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__48724),
            .ce(N__29875),
            .sr(N__48233));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_8_14_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_8_14_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_8_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_8_14_3  (
            .in0(_gnd_net_),
            .in1(N__21104),
            .in2(N__21089),
            .in3(N__21065),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__48724),
            .ce(N__29875),
            .sr(N__48233));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_8_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_8_14_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_8_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21062),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48724),
            .ce(N__29875),
            .sr(N__48233));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_8_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_8_15_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_8_15_0  (
            .in0(N__26375),
            .in1(N__28865),
            .in2(_gnd_net_),
            .in3(N__29309),
            .lcout(\current_shift_inst.control_input_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_8_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_8_15_2 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_8_15_2  (
            .in0(N__26435),
            .in1(N__28967),
            .in2(_gnd_net_),
            .in3(N__29306),
            .lcout(\current_shift_inst.control_input_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_8_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_8_15_3 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_8_15_3  (
            .in0(N__29310),
            .in1(N__26360),
            .in2(_gnd_net_),
            .in3(N__28838),
            .lcout(\current_shift_inst.control_input_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_8_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_8_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_8_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22510),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_8_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_8_15_5 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_8_15_5  (
            .in0(N__29308),
            .in1(N__28898),
            .in2(_gnd_net_),
            .in3(N__26390),
            .lcout(\current_shift_inst.control_input_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_8_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_8_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_8_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29311),
            .lcout(\current_shift_inst.control_input_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_8_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_8_15_7 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_8_15_7  (
            .in0(N__29307),
            .in1(N__28928),
            .in2(_gnd_net_),
            .in3(N__26405),
            .lcout(\current_shift_inst.control_input_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_8_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_8_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_8_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33648),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_8_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_8_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_8_16_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_8_16_2  (
            .in0(N__21260),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48704),
            .ce(N__33742),
            .sr(N__48243));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_8_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_8_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_8_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_8_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33772),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48704),
            .ce(N__33742),
            .sr(N__48243));
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_8_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_8_16_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_inv_LC_8_16_6  (
            .in0(N__37879),
            .in1(N__21185),
            .in2(_gnd_net_),
            .in3(N__22636),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_31 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_8_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_8_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_8_16_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_8_16_7  (
            .in0(_gnd_net_),
            .in1(N__37880),
            .in2(N__21179),
            .in3(N__29446),
            .lcout(\current_shift_inst.un38_control_input_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_8_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_8_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_8_17_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_8_17_2  (
            .in0(N__27126),
            .in1(N__33611),
            .in2(_gnd_net_),
            .in3(N__27086),
            .lcout(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_8_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_8_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_8_17_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_8_17_3  (
            .in0(N__33615),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33272),
            .lcout(\current_shift_inst.un38_control_input_axb_31_s0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_8_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_8_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_8_17_5 .LUT_INIT=16'b1100010111000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_8_17_5  (
            .in0(N__24148),
            .in1(N__24787),
            .in2(N__33617),
            .in3(N__33273),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_8_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_8_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_8_17_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_8_17_6  (
            .in0(N__26922),
            .in1(N__24147),
            .in2(_gnd_net_),
            .in3(N__24786),
            .lcout(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_8_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_8_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_8_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_8_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33771),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48696),
            .ce(N__33741),
            .sr(N__48250));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_8_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_8_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_8_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_8_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26549),
            .lcout(\current_shift_inst.un4_control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_8_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_8_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_8_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_8_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24378),
            .lcout(\current_shift_inst.un4_control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_8_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_8_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_8_18_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_8_18_4  (
            .in0(N__26550),
            .in1(N__26921),
            .in2(_gnd_net_),
            .in3(N__26528),
            .lcout(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_8_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_8_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_8_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_8_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29675),
            .lcout(\current_shift_inst.un4_control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.counter_0_LC_8_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_8_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_8_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_8_19_0  (
            .in0(N__34219),
            .in1(N__21256),
            .in2(_gnd_net_),
            .in3(N__21239),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_19_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__48685),
            .ce(N__32582),
            .sr(N__48263));
    defparam \current_shift_inst.timer_s1.counter_1_LC_8_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_8_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_8_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_8_19_1  (
            .in0(N__34223),
            .in1(N__23956),
            .in2(_gnd_net_),
            .in3(N__21236),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__48685),
            .ce(N__32582),
            .sr(N__48263));
    defparam \current_shift_inst.timer_s1.counter_2_LC_8_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_8_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_8_19_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_8_19_2  (
            .in0(N__34220),
            .in1(N__21231),
            .in2(_gnd_net_),
            .in3(N__21212),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__48685),
            .ce(N__32582),
            .sr(N__48263));
    defparam \current_shift_inst.timer_s1.counter_3_LC_8_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_8_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_8_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_8_19_3  (
            .in0(N__34224),
            .in1(N__21207),
            .in2(_gnd_net_),
            .in3(N__21188),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__48685),
            .ce(N__32582),
            .sr(N__48263));
    defparam \current_shift_inst.timer_s1.counter_4_LC_8_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_8_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_8_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_8_19_4  (
            .in0(N__34221),
            .in1(N__21451),
            .in2(_gnd_net_),
            .in3(N__21431),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__48685),
            .ce(N__32582),
            .sr(N__48263));
    defparam \current_shift_inst.timer_s1.counter_5_LC_8_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_8_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_8_19_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_8_19_5  (
            .in0(N__34225),
            .in1(N__21427),
            .in2(_gnd_net_),
            .in3(N__21407),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__48685),
            .ce(N__32582),
            .sr(N__48263));
    defparam \current_shift_inst.timer_s1.counter_6_LC_8_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_8_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_8_19_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_8_19_6  (
            .in0(N__34222),
            .in1(N__21403),
            .in2(_gnd_net_),
            .in3(N__21383),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__48685),
            .ce(N__32582),
            .sr(N__48263));
    defparam \current_shift_inst.timer_s1.counter_7_LC_8_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_8_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_8_19_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_8_19_7  (
            .in0(N__34226),
            .in1(N__21379),
            .in2(_gnd_net_),
            .in3(N__21359),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__48685),
            .ce(N__32582),
            .sr(N__48263));
    defparam \current_shift_inst.timer_s1.counter_8_LC_8_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_8_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_8_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_8_20_0  (
            .in0(N__34157),
            .in1(N__21355),
            .in2(_gnd_net_),
            .in3(N__21335),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_20_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__48680),
            .ce(N__32584),
            .sr(N__48266));
    defparam \current_shift_inst.timer_s1.counter_9_LC_8_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_8_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_8_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_8_20_1  (
            .in0(N__34161),
            .in1(N__21331),
            .in2(_gnd_net_),
            .in3(N__21311),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__48680),
            .ce(N__32584),
            .sr(N__48266));
    defparam \current_shift_inst.timer_s1.counter_10_LC_8_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_8_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_8_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_8_20_2  (
            .in0(N__34154),
            .in1(N__21307),
            .in2(_gnd_net_),
            .in3(N__21287),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__48680),
            .ce(N__32584),
            .sr(N__48266));
    defparam \current_shift_inst.timer_s1.counter_11_LC_8_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_8_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_8_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_8_20_3  (
            .in0(N__34158),
            .in1(N__21283),
            .in2(_gnd_net_),
            .in3(N__21263),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__48680),
            .ce(N__32584),
            .sr(N__48266));
    defparam \current_shift_inst.timer_s1.counter_12_LC_8_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_8_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_8_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_8_20_4  (
            .in0(N__34155),
            .in1(N__21664),
            .in2(_gnd_net_),
            .in3(N__21644),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__48680),
            .ce(N__32584),
            .sr(N__48266));
    defparam \current_shift_inst.timer_s1.counter_13_LC_8_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_8_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_8_20_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_8_20_5  (
            .in0(N__34159),
            .in1(N__21640),
            .in2(_gnd_net_),
            .in3(N__21620),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__48680),
            .ce(N__32584),
            .sr(N__48266));
    defparam \current_shift_inst.timer_s1.counter_14_LC_8_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_8_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_8_20_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_8_20_6  (
            .in0(N__34156),
            .in1(N__21616),
            .in2(_gnd_net_),
            .in3(N__21596),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__48680),
            .ce(N__32584),
            .sr(N__48266));
    defparam \current_shift_inst.timer_s1.counter_15_LC_8_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_8_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_8_20_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_8_20_7  (
            .in0(N__34160),
            .in1(N__21592),
            .in2(_gnd_net_),
            .in3(N__21572),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__48680),
            .ce(N__32584),
            .sr(N__48266));
    defparam \current_shift_inst.timer_s1.counter_16_LC_8_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_8_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_8_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_8_21_0  (
            .in0(N__34191),
            .in1(N__21568),
            .in2(_gnd_net_),
            .in3(N__21548),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_8_21_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__48676),
            .ce(N__32583),
            .sr(N__48271));
    defparam \current_shift_inst.timer_s1.counter_17_LC_8_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_8_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_8_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_8_21_1  (
            .in0(N__34121),
            .in1(N__21544),
            .in2(_gnd_net_),
            .in3(N__21524),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__48676),
            .ce(N__32583),
            .sr(N__48271));
    defparam \current_shift_inst.timer_s1.counter_18_LC_8_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_8_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_8_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_8_21_2  (
            .in0(N__34192),
            .in1(N__21520),
            .in2(_gnd_net_),
            .in3(N__21500),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__48676),
            .ce(N__32583),
            .sr(N__48271));
    defparam \current_shift_inst.timer_s1.counter_19_LC_8_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_8_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_8_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_8_21_3  (
            .in0(N__34122),
            .in1(N__21496),
            .in2(_gnd_net_),
            .in3(N__21476),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__48676),
            .ce(N__32583),
            .sr(N__48271));
    defparam \current_shift_inst.timer_s1.counter_20_LC_8_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_8_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_8_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_8_21_4  (
            .in0(N__34193),
            .in1(N__21472),
            .in2(_gnd_net_),
            .in3(N__21851),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__48676),
            .ce(N__32583),
            .sr(N__48271));
    defparam \current_shift_inst.timer_s1.counter_21_LC_8_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_8_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_8_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_8_21_5  (
            .in0(N__34123),
            .in1(N__21847),
            .in2(_gnd_net_),
            .in3(N__21827),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__48676),
            .ce(N__32583),
            .sr(N__48271));
    defparam \current_shift_inst.timer_s1.counter_22_LC_8_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_8_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_8_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_8_21_6  (
            .in0(N__34194),
            .in1(N__21823),
            .in2(_gnd_net_),
            .in3(N__21803),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__48676),
            .ce(N__32583),
            .sr(N__48271));
    defparam \current_shift_inst.timer_s1.counter_23_LC_8_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_8_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_8_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_8_21_7  (
            .in0(N__34124),
            .in1(N__21799),
            .in2(_gnd_net_),
            .in3(N__21779),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__48676),
            .ce(N__32583),
            .sr(N__48271));
    defparam \current_shift_inst.timer_s1.counter_24_LC_8_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_8_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_8_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_8_22_0  (
            .in0(N__34204),
            .in1(N__21775),
            .in2(_gnd_net_),
            .in3(N__21755),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_8_22_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__48670),
            .ce(N__32588),
            .sr(N__48275));
    defparam \current_shift_inst.timer_s1.counter_25_LC_8_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_8_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_8_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_8_22_1  (
            .in0(N__34208),
            .in1(N__21751),
            .in2(_gnd_net_),
            .in3(N__21731),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__48670),
            .ce(N__32588),
            .sr(N__48275));
    defparam \current_shift_inst.timer_s1.counter_26_LC_8_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_8_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_8_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_8_22_2  (
            .in0(N__34205),
            .in1(N__21727),
            .in2(_gnd_net_),
            .in3(N__21707),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__48670),
            .ce(N__32588),
            .sr(N__48275));
    defparam \current_shift_inst.timer_s1.counter_27_LC_8_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_8_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_8_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_8_22_3  (
            .in0(N__34209),
            .in1(N__21703),
            .in2(_gnd_net_),
            .in3(N__21683),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__48670),
            .ce(N__32588),
            .sr(N__48275));
    defparam \current_shift_inst.timer_s1.counter_28_LC_8_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_8_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_8_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_8_22_4  (
            .in0(N__34206),
            .in1(N__21680),
            .in2(_gnd_net_),
            .in3(N__21668),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__48670),
            .ce(N__32588),
            .sr(N__48275));
    defparam \current_shift_inst.timer_s1.counter_29_LC_8_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_8_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_8_22_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_8_22_5  (
            .in0(N__21905),
            .in1(N__34207),
            .in2(_gnd_net_),
            .in3(N__21908),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48670),
            .ce(N__32588),
            .sr(N__48275));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_8_23_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_8_23_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_8_23_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_8_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30286),
            .lcout(\current_shift_inst.un4_control_input_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_8_23_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_8_23_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_8_23_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_8_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30555),
            .lcout(\current_shift_inst.un4_control_input_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.S2_LC_8_29_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.S2_LC_8_29_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S2_LC_8_29_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S2_LC_8_29_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31732),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48648),
            .ce(),
            .sr(N__48286));
    defparam GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_8_30_2.C_ON=1'b0;
    defparam GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_8_30_2.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_8_30_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_8_30_2 (
            .in0(N__48812),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_clock_output_0_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_2_5.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_2_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_2_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH1_MIN_D1_LC_9_2_5 (
            .in0(N__21878),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_min_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48808),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_9_3_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_9_3_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_9_3_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_15_LC_9_3_5  (
            .in0(N__21867),
            .in1(N__23293),
            .in2(_gnd_net_),
            .in3(N__41891),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48807),
            .ce(N__28514),
            .sr(N__48141));
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_9_4_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_9_4_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_9_4_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_15_LC_9_4_1  (
            .in0(N__21868),
            .in1(N__23294),
            .in2(_gnd_net_),
            .in3(N__41895),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48806),
            .ce(N__36608),
            .sr(N__48149));
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_9_5_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_9_5_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_9_5_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_20_LC_9_5_7  (
            .in0(N__31374),
            .in1(N__31357),
            .in2(_gnd_net_),
            .in3(N__41879),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48801),
            .ce(N__28513),
            .sr(N__48157));
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_9_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_9_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_9_6_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_7_LC_9_6_3  (
            .in0(N__41850),
            .in1(N__25058),
            .in2(_gnd_net_),
            .in3(N__25102),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48797),
            .ce(N__28512),
            .sr(N__48166));
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_9_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_9_6_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_9_6_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_5_LC_9_6_7  (
            .in0(N__41849),
            .in1(N__23178),
            .in2(_gnd_net_),
            .in3(N__23134),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48797),
            .ce(N__28512),
            .sr(N__48166));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_9_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_9_7_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_9_7_3  (
            .in0(N__31584),
            .in1(N__31502),
            .in2(N__41943),
            .in3(N__38249),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_9_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_9_7_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_9_7_4  (
            .in0(N__23579),
            .in1(N__28577),
            .in2(N__23439),
            .in3(N__28640),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_9_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_9_7_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_9_7_5  (
            .in0(N__21968),
            .in1(N__23981),
            .in2(N__21962),
            .in3(N__23249),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_9_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_9_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_9_7_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_13_LC_9_7_6  (
            .in0(N__23532),
            .in1(N__41668),
            .in2(_gnd_net_),
            .in3(N__23513),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48787),
            .ce(N__36601),
            .sr(N__48174));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_9_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_9_8_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_9_8_0  (
            .in0(N__22997),
            .in1(N__23039),
            .in2(N__23098),
            .in3(N__23852),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_9_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_9_8_1 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(N__31878),
            .in2(N__21959),
            .in3(N__28166),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_9_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_9_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_9_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21955),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48778),
            .ce(N__29888),
            .sr(N__48183));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_9_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_9_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_9_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21928),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48778),
            .ce(N__29888),
            .sr(N__48183));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_9_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_9_8_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_9_8_5  (
            .in0(N__23040),
            .in1(N__23066),
            .in2(_gnd_net_),
            .in3(N__41743),
            .lcout(elapsed_time_ns_1_RNIE03T9_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_9_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_9_8_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_9_8_6  (
            .in0(N__22998),
            .in1(N__41653),
            .in2(_gnd_net_),
            .in3(N__23021),
            .lcout(elapsed_time_ns_1_RNIF13T9_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_9_8_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_9_8_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_9_8_7  (
            .in0(N__23093),
            .in1(N__23117),
            .in2(_gnd_net_),
            .in3(N__41742),
            .lcout(elapsed_time_ns_1_RNIG23T9_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_9_0 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_9_0  (
            .in0(N__22022),
            .in1(N__25964),
            .in2(N__25997),
            .in3(N__22004),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_9_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_9_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_9_9_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_2_LC_9_9_4  (
            .in0(N__23041),
            .in1(N__23064),
            .in2(_gnd_net_),
            .in3(N__41666),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48768),
            .ce(N__28509),
            .sr(N__48193));
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_9_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_9_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_9_9_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_3_LC_9_9_5  (
            .in0(N__41665),
            .in1(N__23019),
            .in2(_gnd_net_),
            .in3(N__22999),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48768),
            .ce(N__28509),
            .sr(N__48193));
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_9_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_9_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_9_9_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_4_LC_9_9_6  (
            .in0(N__23115),
            .in1(N__23097),
            .in2(_gnd_net_),
            .in3(N__41667),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48768),
            .ce(N__28509),
            .sr(N__48193));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_9_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_9_10_0 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_9_10_0  (
            .in0(N__25936),
            .in1(N__23542),
            .in2(N__25913),
            .in3(N__21983),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_9_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_9_10_1 .LUT_INIT=16'b1011000011111011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_9_10_1  (
            .in0(N__21982),
            .in1(N__25937),
            .in2(N__23546),
            .in3(N__25912),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_9_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_9_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_9_10_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_6_LC_9_10_4  (
            .in0(N__41787),
            .in1(N__24909),
            .in2(_gnd_net_),
            .in3(N__24944),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48760),
            .ce(N__28505),
            .sr(N__48203));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_9_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_9_10_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_9_10_5  (
            .in0(N__23234),
            .in1(N__41786),
            .in2(_gnd_net_),
            .in3(N__23212),
            .lcout(elapsed_time_ns_1_RNIK63T9_0_8),
            .ltout(elapsed_time_ns_1_RNIK63T9_0_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_9_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_9_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_9_10_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_8_LC_9_10_6  (
            .in0(N__41788),
            .in1(_gnd_net_),
            .in2(N__22124),
            .in3(N__23235),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48760),
            .ce(N__28505),
            .sr(N__48203));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_9_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_9_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(N__23831),
            .in2(N__22121),
            .in3(N__25416),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_9_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_9_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_9_11_1  (
            .in0(_gnd_net_),
            .in1(N__22112),
            .in2(N__22103),
            .in3(N__25682),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_9_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_9_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(N__22082),
            .in2(N__22094),
            .in3(N__25655),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_9_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_9_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(N__22076),
            .in2(N__22067),
            .in3(N__25637),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_9_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_9_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(N__22058),
            .in2(N__22046),
            .in3(N__25616),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_9_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_9_11_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_9_11_5  (
            .in0(N__25598),
            .in1(N__22037),
            .in2(N__22031),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_9_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_9_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_9_11_6  (
            .in0(_gnd_net_),
            .in1(N__22262),
            .in2(N__22253),
            .in3(N__25580),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_9_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_9_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_9_11_7  (
            .in0(_gnd_net_),
            .in1(N__22244),
            .in2(N__22235),
            .in3(N__25559),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_9_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_9_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(N__22214),
            .in2(N__22226),
            .in3(N__25541),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_9_12_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_9_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_9_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__22202),
            .in2(N__22193),
            .in3(N__25826),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_9_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_9_12_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_9_12_2  (
            .in0(N__25808),
            .in1(N__22184),
            .in2(N__22175),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_9_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_9_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(N__22163),
            .in2(N__28679),
            .in3(N__25790),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_9_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_9_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(N__23474),
            .in2(N__22157),
            .in3(N__25772),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_9_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_9_12_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_9_12_5  (
            .in0(N__25754),
            .in1(N__22145),
            .in2(N__22133),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_9_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_9_12_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_9_12_6  (
            .in0(N__25736),
            .in1(N__22361),
            .in2(N__22349),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_9_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_9_12_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_9_12_7  (
            .in0(_gnd_net_),
            .in1(N__24068),
            .in2(N__24164),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_9_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_9_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__22340),
            .in2(N__22331),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_9_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_9_13_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(N__22313),
            .in2(N__22304),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_9_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_9_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__22289),
            .in2(N__22277),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_9_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_9_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__27953),
            .in2(N__28004),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_9_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_9_13_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(N__24197),
            .in2(N__28382),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_9_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_9_13_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(N__28103),
            .in2(N__28019),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_9_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_9_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__23765),
            .in2(N__23810),
            .in3(N__22493),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_9_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_9_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22490),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_9_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_9_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__24293),
            .in2(N__24284),
            .in3(N__24282),
            .lcout(\current_shift_inst.control_input_18 ),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\current_shift_inst.control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_9_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_9_14_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__22499),
            .in2(_gnd_net_),
            .in3(N__22463),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_0 ),
            .carryout(\current_shift_inst.control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_9_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_9_14_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(N__22460),
            .in2(_gnd_net_),
            .in3(N__22442),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_1 ),
            .carryout(\current_shift_inst.control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_9_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_9_14_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__22649),
            .in2(_gnd_net_),
            .in3(N__22427),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_2 ),
            .carryout(\current_shift_inst.control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_9_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_9_14_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(N__22424),
            .in2(_gnd_net_),
            .in3(N__22406),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_3 ),
            .carryout(\current_shift_inst.control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_9_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_9_14_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(N__22403),
            .in2(_gnd_net_),
            .in3(N__22385),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_4 ),
            .carryout(\current_shift_inst.control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_9_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_9_14_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__22382),
            .in2(_gnd_net_),
            .in3(N__22364),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_5 ),
            .carryout(\current_shift_inst.control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_9_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_9_14_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(N__22622),
            .in2(_gnd_net_),
            .in3(N__22604),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_6 ),
            .carryout(\current_shift_inst.control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_9_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_9_15_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__29366),
            .in2(_gnd_net_),
            .in3(N__22589),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\current_shift_inst.control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_9_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_9_15_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__29342),
            .in2(_gnd_net_),
            .in3(N__22574),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_8 ),
            .carryout(\current_shift_inst.control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_9_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_9_15_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__29231),
            .in2(_gnd_net_),
            .in3(N__22559),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_9 ),
            .carryout(\current_shift_inst.control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_9_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_9_15_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__29390),
            .in2(_gnd_net_),
            .in3(N__22544),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_10 ),
            .carryout(\current_shift_inst.control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_9_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_9_15_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(N__22541),
            .in2(_gnd_net_),
            .in3(N__22523),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_11 ),
            .carryout(\current_shift_inst.control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_9_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_9_15_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(N__29305),
            .in2(_gnd_net_),
            .in3(N__22520),
            .lcout(\current_shift_inst.control_input_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_9_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_9_15_6 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_9_15_6  (
            .in0(N__29303),
            .in1(N__26450),
            .in2(_gnd_net_),
            .in3(N__28979),
            .lcout(\current_shift_inst.control_input_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_9_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_9_15_7 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_9_15_7  (
            .in0(N__26420),
            .in1(N__28955),
            .in2(_gnd_net_),
            .in3(N__29304),
            .lcout(\current_shift_inst.control_input_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_9_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_9_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(N__31958),
            .in2(N__22643),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_16_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_9_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_9_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(N__37866),
            .in2(N__24215),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_0 ),
            .carryout(\current_shift_inst.un10_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_9_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_9_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(N__24320),
            .in2(N__37906),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_1 ),
            .carryout(\current_shift_inst.un10_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_9_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_9_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(N__37870),
            .in2(N__24587),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_2 ),
            .carryout(\current_shift_inst.un10_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_9_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_9_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(N__24326),
            .in2(N__37907),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_3 ),
            .carryout(\current_shift_inst.un10_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_9_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_9_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_LC_9_16_5  (
            .in0(_gnd_net_),
            .in1(N__37874),
            .in2(N__24356),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_4 ),
            .carryout(\current_shift_inst.un10_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_9_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_9_16_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(N__24170),
            .in2(N__37908),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_5 ),
            .carryout(\current_shift_inst.un10_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_9_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_9_16_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_LC_9_16_7  (
            .in0(_gnd_net_),
            .in1(N__37878),
            .in2(N__24347),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_6 ),
            .carryout(\current_shift_inst.un10_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_9_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_9_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_LC_9_17_0  (
            .in0(_gnd_net_),
            .in1(N__22667),
            .in2(N__37905),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_17_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_9_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_9_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_LC_9_17_1  (
            .in0(_gnd_net_),
            .in1(N__37865),
            .in2(N__24308),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_8 ),
            .carryout(\current_shift_inst.un10_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_9_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_9_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_LC_9_17_2  (
            .in0(_gnd_net_),
            .in1(N__22754),
            .in2(N__37902),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_9 ),
            .carryout(\current_shift_inst.un10_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_9_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_9_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_LC_9_17_3  (
            .in0(_gnd_net_),
            .in1(N__37853),
            .in2(N__24335),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_10 ),
            .carryout(\current_shift_inst.un10_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_9_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_9_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_LC_9_17_4  (
            .in0(_gnd_net_),
            .in1(N__22739),
            .in2(N__37903),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_11 ),
            .carryout(\current_shift_inst.un10_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_9_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_9_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_LC_9_17_5  (
            .in0(_gnd_net_),
            .in1(N__37857),
            .in2(N__22661),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_12 ),
            .carryout(\current_shift_inst.un10_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_9_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_9_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_LC_9_17_6  (
            .in0(_gnd_net_),
            .in1(N__24314),
            .in2(N__37904),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_13 ),
            .carryout(\current_shift_inst.un10_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_9_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_9_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_LC_9_17_7  (
            .in0(_gnd_net_),
            .in1(N__37861),
            .in2(N__24404),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_14 ),
            .carryout(\current_shift_inst.un10_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_9_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_9_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(N__37834),
            .in2(N__22775),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_18_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_9_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_9_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_LC_9_18_1  (
            .in0(_gnd_net_),
            .in1(N__26855),
            .in2(N__37898),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_16 ),
            .carryout(\current_shift_inst.un10_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_9_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_9_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_LC_9_18_2  (
            .in0(_gnd_net_),
            .in1(N__37838),
            .in2(N__22817),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_17 ),
            .carryout(\current_shift_inst.un10_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_9_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_9_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_9_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_LC_9_18_3  (
            .in0(_gnd_net_),
            .in1(N__26660),
            .in2(N__37899),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_18 ),
            .carryout(\current_shift_inst.un10_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_9_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_9_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_LC_9_18_4  (
            .in0(_gnd_net_),
            .in1(N__37842),
            .in2(N__26687),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_19 ),
            .carryout(\current_shift_inst.un10_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_9_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_9_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_LC_9_18_5  (
            .in0(_gnd_net_),
            .in1(N__22673),
            .in2(N__37900),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_20 ),
            .carryout(\current_shift_inst.un10_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_9_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_9_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_LC_9_18_6  (
            .in0(_gnd_net_),
            .in1(N__37846),
            .in2(N__26702),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_21 ),
            .carryout(\current_shift_inst.un10_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_9_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_9_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(N__22730),
            .in2(N__37901),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_22 ),
            .carryout(\current_shift_inst.un10_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_9_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_9_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__37717),
            .in2(N__22688),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_9_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_9_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__22694),
            .in2(N__37831),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_24 ),
            .carryout(\current_shift_inst.un10_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_9_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_9_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(N__37721),
            .in2(N__22721),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_25 ),
            .carryout(\current_shift_inst.un10_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_9_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_9_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(N__22679),
            .in2(N__37832),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_26 ),
            .carryout(\current_shift_inst.un10_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_9_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_9_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(N__37725),
            .in2(N__22709),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_27 ),
            .carryout(\current_shift_inst.un10_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_9_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_9_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_LC_9_19_5  (
            .in0(_gnd_net_),
            .in1(N__22745),
            .in2(N__37833),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_28 ),
            .carryout(\current_shift_inst.un10_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_9_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_9_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(N__37729),
            .in2(N__22763),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_29 ),
            .carryout(\current_shift_inst.un10_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_9_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_9_19_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(N__33589),
            .in2(_gnd_net_),
            .in3(N__22697),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_9_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_9_20_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_9_20_0  (
            .in0(N__33607),
            .in1(N__27189),
            .in2(_gnd_net_),
            .in3(N__27148),
            .lcout(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_9_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_9_20_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_9_20_1  (
            .in0(N__26984),
            .in1(N__27051),
            .in2(_gnd_net_),
            .in3(N__27009),
            .lcout(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_9_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_9_20_2 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_9_20_2  (
            .in0(N__33608),
            .in1(N__33849),
            .in2(N__33811),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_9_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_9_20_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_9_20_3  (
            .in0(N__29532),
            .in1(N__26983),
            .in2(_gnd_net_),
            .in3(N__29478),
            .lcout(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_9_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_9_20_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_9_20_4  (
            .in0(N__33610),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31999),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_9_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_9_20_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_9_20_5  (
            .in0(N__30405),
            .in1(N__26981),
            .in2(_gnd_net_),
            .in3(N__30369),
            .lcout(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_9_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_9_20_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_9_20_6  (
            .in0(N__33609),
            .in1(N__30573),
            .in2(_gnd_net_),
            .in3(N__30525),
            .lcout(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_9_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_9_20_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_9_20_7  (
            .in0(N__32328),
            .in1(N__26982),
            .in2(_gnd_net_),
            .in3(N__32283),
            .lcout(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_9_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_9_21_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_9_21_0  (
            .in0(N__26977),
            .in1(N__30069),
            .in2(_gnd_net_),
            .in3(N__30090),
            .lcout(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_9_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_9_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_9_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32139),
            .lcout(\current_shift_inst.un4_control_input_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_9_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_9_21_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_9_21_2  (
            .in0(N__33547),
            .in1(N__26643),
            .in2(_gnd_net_),
            .in3(N__26604),
            .lcout(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_9_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_9_21_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_9_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27044),
            .lcout(\current_shift_inst.un4_control_input_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_9_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_9_21_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30396),
            .lcout(\current_shift_inst.un4_control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_9_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_9_21_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_9_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30159),
            .lcout(\current_shift_inst.un4_control_input_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_9_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_9_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_9_21_6 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_9_21_6  (
            .in0(N__26976),
            .in1(N__29964),
            .in2(_gnd_net_),
            .in3(N__30007),
            .lcout(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_9_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_9_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_9_21_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_9_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32459),
            .lcout(\current_shift_inst.un4_control_input_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_9_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_9_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_9_22_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_9_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24135),
            .lcout(\current_shift_inst.un4_control_input_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_9_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_9_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_9_22_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_9_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27180),
            .lcout(\current_shift_inst.un4_control_input_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_9_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_9_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_9_22_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_9_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30056),
            .lcout(\current_shift_inst.un4_control_input_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_9_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_9_22_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_9_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27119),
            .lcout(\current_shift_inst.un4_control_input_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_9_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_9_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_9_22_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_9_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30236),
            .lcout(\current_shift_inst.un4_control_input_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_9_23_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_9_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_9_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_2_LC_9_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22805),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48661),
            .ce(),
            .sr(N__48276));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_9_23_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_9_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_9_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_9_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22928),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48661),
            .ce(),
            .sr(N__48276));
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_9_23_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_9_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_9_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_1_LC_9_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22901),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48661),
            .ce(),
            .sr(N__48276));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_9_24_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_9_24_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_9_24_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_9_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22871),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48658),
            .ce(),
            .sr(N__48279));
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_9_24_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_9_24_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_9_24_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_13_LC_9_24_6  (
            .in0(N__22847),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48658),
            .ce(),
            .sr(N__48279));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_10_4_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_10_4_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_10_4_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_10_4_4  (
            .in0(N__31378),
            .in1(N__31356),
            .in2(_gnd_net_),
            .in3(N__41779),
            .lcout(elapsed_time_ns_1_RNIU0DN9_0_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_10_5_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_10_5_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_10_5_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_10_5_1  (
            .in0(N__23335),
            .in1(N__27709),
            .in2(N__27743),
            .in3(N__23197),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_10_5_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_10_5_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_10_5_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_10_5_5  (
            .in0(N__41783),
            .in1(N__23179),
            .in2(_gnd_net_),
            .in3(N__23135),
            .lcout(elapsed_time_ns_1_RNIH33T9_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_10_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_10_6_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_10_6_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_30_LC_10_6_2  (
            .in0(N__41771),
            .in1(N__23463),
            .in2(_gnd_net_),
            .in3(N__23440),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48780),
            .ce(N__36597),
            .sr(N__48150));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_10_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_10_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_10_6_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_LC_10_6_3  (
            .in0(N__25101),
            .in1(N__25053),
            .in2(_gnd_net_),
            .in3(N__41775),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48780),
            .ce(N__36597),
            .sr(N__48150));
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_10_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_10_6_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_10_6_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_31_LC_10_6_4  (
            .in0(N__41772),
            .in1(N__23939),
            .in2(_gnd_net_),
            .in3(N__23380),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48780),
            .ce(N__36597),
            .sr(N__48150));
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_10_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_10_6_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_10_6_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_24_LC_10_6_5  (
            .in0(N__38200),
            .in1(N__38260),
            .in2(_gnd_net_),
            .in3(N__41774),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48780),
            .ce(N__36597),
            .sr(N__48150));
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_10_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_10_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_10_6_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_5_LC_10_6_6  (
            .in0(N__41773),
            .in1(N__23180),
            .in2(_gnd_net_),
            .in3(N__23133),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48780),
            .ce(N__36597),
            .sr(N__48150));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_10_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_10_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_10_7_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_LC_10_7_0  (
            .in0(N__23116),
            .in1(N__23099),
            .in2(_gnd_net_),
            .in3(N__41659),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48769),
            .ce(N__36605),
            .sr(N__48158));
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_10_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_10_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_10_7_1 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_2_LC_10_7_1  (
            .in0(N__41655),
            .in1(N__23065),
            .in2(N__23048),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48769),
            .ce(N__36605),
            .sr(N__48158));
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_10_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_10_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_10_7_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_3_LC_10_7_3  (
            .in0(N__41656),
            .in1(N__23020),
            .in2(_gnd_net_),
            .in3(N__23003),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48769),
            .ce(N__36605),
            .sr(N__48158));
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_10_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_10_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_10_7_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_19_LC_10_7_4  (
            .in0(N__22976),
            .in1(N__24057),
            .in2(_gnd_net_),
            .in3(N__41658),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48769),
            .ce(N__36605),
            .sr(N__48158));
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_10_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_10_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_10_7_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_1_LC_10_7_5  (
            .in0(N__41654),
            .in1(N__23891),
            .in2(_gnd_net_),
            .in3(N__23856),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48769),
            .ce(N__36605),
            .sr(N__48158));
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_10_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_10_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_10_7_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_18_LC_10_7_6  (
            .in0(N__22952),
            .in1(N__24022),
            .in2(_gnd_net_),
            .in3(N__41657),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48769),
            .ce(N__36605),
            .sr(N__48158));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_10_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_10_8_0 .LUT_INIT=16'b0100110101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_10_8_0  (
            .in0(N__27776),
            .in1(N__23350),
            .in2(N__27554),
            .in3(N__23360),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_10_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_10_8_1 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_10_8_1  (
            .in0(N__23359),
            .in1(N__27775),
            .in2(N__23351),
            .in3(N__27553),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_10_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_10_8_2 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_10_8_2  (
            .in0(N__27739),
            .in1(N__23339),
            .in2(N__23201),
            .in3(N__27710),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_10_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_10_8_3 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_10_8_3  (
            .in0(N__23937),
            .in1(N__23324),
            .in2(N__23318),
            .in3(N__23303),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_10_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_10_8_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_10_8_4  (
            .in0(N__27297),
            .in1(_gnd_net_),
            .in2(N__23297),
            .in3(N__27327),
            .lcout(elapsed_time_ns_1_RNI35CN9_0_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_10_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_10_8_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_10_8_5  (
            .in0(N__41652),
            .in1(N__23465),
            .in2(_gnd_net_),
            .in3(N__23432),
            .lcout(elapsed_time_ns_1_RNIV2EN9_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_10_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_10_8_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_10_8_6  (
            .in0(N__23511),
            .in1(N__23533),
            .in2(_gnd_net_),
            .in3(N__41651),
            .lcout(elapsed_time_ns_1_RNI02CN9_0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_10_8_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_10_8_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_10_8_7  (
            .in0(N__23282),
            .in1(N__23510),
            .in2(N__30769),
            .in3(N__27296),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_10_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_10_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_10_9_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_8_LC_10_9_0  (
            .in0(N__23243),
            .in1(N__41663),
            .in2(_gnd_net_),
            .in3(N__23213),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48748),
            .ce(N__36606),
            .sr(N__48175));
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_10_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_10_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_10_9_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_25_LC_10_9_1  (
            .in0(N__41660),
            .in1(N__28662),
            .in2(_gnd_net_),
            .in3(N__28645),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48748),
            .ce(N__36606),
            .sr(N__48175));
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_10_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_10_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_10_9_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_10_LC_10_9_2  (
            .in0(N__23741),
            .in1(N__23714),
            .in2(_gnd_net_),
            .in3(N__41664),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48748),
            .ce(N__36606),
            .sr(N__48175));
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_10_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_10_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_10_9_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_9_LC_10_9_3  (
            .in0(N__41662),
            .in1(N__23677),
            .in2(_gnd_net_),
            .in3(N__23651),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48748),
            .ce(N__36606),
            .sr(N__48175));
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_10_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_10_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_10_9_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_29_LC_10_9_7  (
            .in0(N__41661),
            .in1(N__23618),
            .in2(_gnd_net_),
            .in3(N__23591),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48748),
            .ce(N__36606),
            .sr(N__48175));
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_10_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_10_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_10_10_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_21_LC_10_10_0  (
            .in0(N__41419),
            .in1(N__41942),
            .in2(_gnd_net_),
            .in3(N__41794),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48736),
            .ce(N__28506),
            .sr(N__48184));
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_10_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_10_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_10_10_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_16_LC_10_10_2  (
            .in0(N__27328),
            .in1(N__27301),
            .in2(_gnd_net_),
            .in3(N__41793),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48736),
            .ce(N__28506),
            .sr(N__48184));
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_10_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_10_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_10_10_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_17_LC_10_10_3  (
            .in0(N__41789),
            .in1(N__25127),
            .in2(_gnd_net_),
            .in3(N__25165),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48736),
            .ce(N__28506),
            .sr(N__48184));
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_10_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_10_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_10_10_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_13_LC_10_10_4  (
            .in0(N__23534),
            .in1(N__41792),
            .in2(_gnd_net_),
            .in3(N__23512),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48736),
            .ce(N__28506),
            .sr(N__48184));
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_10_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_10_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_10_10_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_30_LC_10_10_5  (
            .in0(N__41791),
            .in1(N__23464),
            .in2(_gnd_net_),
            .in3(N__23441),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48736),
            .ce(N__28506),
            .sr(N__48184));
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_10_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_10_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_10_10_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_31_LC_10_10_6  (
            .in0(N__41795),
            .in1(N__23384),
            .in2(_gnd_net_),
            .in3(N__23933),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48736),
            .ce(N__28506),
            .sr(N__48184));
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_10_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_10_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_10_10_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_1_LC_10_10_7  (
            .in0(N__41790),
            .in1(N__23884),
            .in2(_gnd_net_),
            .in3(N__23863),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48736),
            .ce(N__28506),
            .sr(N__48184));
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_30_LC_10_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_30_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_30_LC_10_11_0 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_RNISIH31_30_LC_10_11_0  (
            .in0(N__23776),
            .in1(N__26232),
            .in2(N__26045),
            .in3(N__23788),
            .lcout(),
            .ltout(\phase_controller_inst2.stoper_hc.un4_running_df30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIEABO2_28_LC_10_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIEABO2_28_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIEABO2_28_LC_10_11_1 .LUT_INIT=16'b1111110101011101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIEABO2_28_LC_10_11_1  (
            .in0(N__28210),
            .in1(N__23800),
            .in2(N__23825),
            .in3(N__23822),
            .lcout(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_10_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_10_11_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_10_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23813),
            .in3(N__28256),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_0_30_LC_10_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_0_30_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_0_30_LC_10_11_3 .LUT_INIT=16'b0000100011001110;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_RNISIH31_0_30_LC_10_11_3  (
            .in0(N__23787),
            .in1(N__26040),
            .in2(N__26236),
            .in3(N__23775),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3_28_LC_10_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3_28_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3_28_LC_10_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3_28_LC_10_11_4  (
            .in0(_gnd_net_),
            .in1(N__28257),
            .in2(_gnd_net_),
            .in3(N__23752),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_10_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_10_11_5 .LUT_INIT=16'b1000110011101111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_10_11_5  (
            .in0(N__23789),
            .in1(N__26044),
            .in2(N__26237),
            .in3(N__23777),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_10_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_10_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_10_11_6 .LUT_INIT=16'b0001010001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_10_11_6  (
            .in0(N__26203),
            .in1(N__25420),
            .in2(N__23756),
            .in3(N__28261),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48726),
            .ce(),
            .sr(N__48194));
    defparam \phase_controller_inst2.stoper_hc.running_LC_10_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_LC_10_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.running_LC_10_11_7 .LUT_INIT=16'b1101111101010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_LC_10_11_7  (
            .in0(N__28211),
            .in1(N__28237),
            .in2(N__28262),
            .in3(N__28297),
            .lcout(\phase_controller_inst2.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48726),
            .ce(),
            .sr(N__48194));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_10_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_10_12_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_10_12_0  (
            .in0(N__33606),
            .in1(N__30259),
            .in2(N__33278),
            .in3(N__30212),
            .lcout(\current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_10_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_10_12_1 .LUT_INIT=16'b0010001010110010;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_10_12_1  (
            .in0(N__24098),
            .in1(N__25699),
            .in2(N__24085),
            .in3(N__25717),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_10_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_10_12_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_10_12_2  (
            .in0(N__33605),
            .in1(N__24152),
            .in2(N__33277),
            .in3(N__24788),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D2_LC_10_12_4.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_10_12_4.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_10_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D2_LC_10_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24113),
            .lcout(il_min_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48716),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_10_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_10_12_5 .LUT_INIT=16'b1011001010111011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_10_12_5  (
            .in0(N__24097),
            .in1(N__25698),
            .in2(N__24086),
            .in3(N__25716),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_10_12_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_10_12_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_10_12_7  (
            .in0(N__24042),
            .in1(N__25154),
            .in2(N__31346),
            .in3(N__24005),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_10_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_10_13_0 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_10_13_0  (
            .in0(N__33603),
            .in1(N__24568),
            .in2(N__28331),
            .in3(N__24187),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_10_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_10_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_10_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23966),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48706),
            .ce(N__33743),
            .sr(N__48210));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_10_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_10_13_3 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_10_13_3  (
            .in0(N__24569),
            .in1(N__33604),
            .in2(N__24191),
            .in3(N__28330),
            .lcout(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_10_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_10_13_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_10_13_4  (
            .in0(N__26985),
            .in1(N__24567),
            .in2(_gnd_net_),
            .in3(N__24186),
            .lcout(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_10_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_10_14_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_10_14_0  (
            .in0(N__33551),
            .in1(N__24262),
            .in2(N__33280),
            .in3(N__24697),
            .lcout(\current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_10_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_10_14_1 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_10_14_1  (
            .in0(N__32426),
            .in1(N__33550),
            .in2(N__32384),
            .in3(N__33228),
            .lcout(\current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_10_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_10_14_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_10_14_2  (
            .in0(N__33553),
            .in1(N__24440),
            .in2(N__33279),
            .in3(N__24620),
            .lcout(\current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_10_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_10_14_3 .LUT_INIT=16'b1111000001010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_10_14_3  (
            .in0(N__24394),
            .in1(N__33229),
            .in2(N__24500),
            .in3(N__33549),
            .lcout(\current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_14_4 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_14_4  (
            .in0(N__28469),
            .in1(N__28449),
            .in2(N__28426),
            .in3(N__28400),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_10_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_10_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_10_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24185),
            .lcout(\current_shift_inst.un4_control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_10_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_10_14_7 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_10_14_7  (
            .in0(N__29582),
            .in1(N__33230),
            .in2(N__29636),
            .in3(N__33552),
            .lcout(\current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_10_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_10_15_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_10_15_0  (
            .in0(N__26964),
            .in1(N__29628),
            .in2(_gnd_net_),
            .in3(N__29574),
            .lcout(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_10_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_10_15_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_10_15_2  (
            .in0(N__26965),
            .in1(N__24249),
            .in2(_gnd_net_),
            .in3(N__24696),
            .lcout(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_10_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_10_15_4 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_10_15_4  (
            .in0(N__26312),
            .in1(N__28796),
            .in2(_gnd_net_),
            .in3(N__29301),
            .lcout(\current_shift_inst.control_input_axb_0 ),
            .ltout(\current_shift_inst.control_input_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_10_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_10_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_10_15_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_0_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24287),
            .in3(N__24283),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48689),
            .ce(),
            .sr(N__48222));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_10_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_10_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29302),
            .lcout(\current_shift_inst.N_1288_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_10_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_10_16_0 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_10_16_0  (
            .in0(N__33555),
            .in1(N__24395),
            .in2(N__24499),
            .in3(N__33209),
            .lcout(\current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_10_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_10_16_1 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_10_16_1  (
            .in0(N__24619),
            .in1(N__33560),
            .in2(N__33276),
            .in3(N__24436),
            .lcout(\current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_10_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_10_16_2 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_10_16_2  (
            .in0(N__33556),
            .in1(N__33210),
            .in2(N__29693),
            .in3(N__29719),
            .lcout(\current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_10_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_10_16_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_10_16_3  (
            .in0(N__30500),
            .in1(N__33558),
            .in2(N__33274),
            .in3(N__30452),
            .lcout(\current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_10_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_10_16_4 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_10_16_4  (
            .in0(N__33554),
            .in1(N__33208),
            .in2(N__29816),
            .in3(N__29768),
            .lcout(\current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_10_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_10_16_5 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_10_16_5  (
            .in0(N__33211),
            .in1(N__24698),
            .in2(N__24263),
            .in3(N__33557),
            .lcout(\current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_10_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_10_16_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_10_16_6  (
            .in0(N__24435),
            .in1(N__26993),
            .in2(_gnd_net_),
            .in3(N__24618),
            .lcout(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_10_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_10_16_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_10_16_7  (
            .in0(N__32338),
            .in1(N__33559),
            .in2(N__33275),
            .in3(N__32290),
            .lcout(\current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_10_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_10_17_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_10_17_0  (
            .in0(N__24387),
            .in1(N__26939),
            .in2(_gnd_net_),
            .in3(N__24483),
            .lcout(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_10_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_10_17_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_10_17_1  (
            .in0(N__33234),
            .in1(N__33561),
            .in2(N__26566),
            .in3(N__26526),
            .lcout(\current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_10_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_10_17_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_10_17_2  (
            .in0(N__29691),
            .in1(N__26940),
            .in2(_gnd_net_),
            .in3(N__29709),
            .lcout(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_10_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_10_17_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_10_17_3  (
            .in0(N__26941),
            .in1(N__30495),
            .in2(_gnd_net_),
            .in3(N__30450),
            .lcout(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_10_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_10_17_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_10_17_4  (
            .in0(N__32418),
            .in1(N__26938),
            .in2(_gnd_net_),
            .in3(N__32362),
            .lcout(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_17_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_17_5  (
            .in0(N__26936),
            .in1(N__32667),
            .in2(_gnd_net_),
            .in3(N__32625),
            .lcout(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_17_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_17_6  (
            .in0(N__32238),
            .in1(N__26942),
            .in2(_gnd_net_),
            .in3(N__32187),
            .lcout(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_10_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_10_17_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_10_17_7  (
            .in0(N__26937),
            .in1(N__29802),
            .in2(_gnd_net_),
            .in3(N__29760),
            .lcout(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_10_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_10_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_10_18_0  (
            .in0(_gnd_net_),
            .in1(N__24578),
            .in2(N__33712),
            .in3(N__33708),
            .lcout(\current_shift_inst.un4_control_input1_2 ),
            .ltout(),
            .carryin(bfn_10_18_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_10_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_10_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_10_18_1  (
            .in0(_gnd_net_),
            .in1(N__24554),
            .in2(_gnd_net_),
            .in3(N__24542),
            .lcout(\current_shift_inst.un4_control_input1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_10_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_10_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_10_18_2  (
            .in0(_gnd_net_),
            .in1(N__24539),
            .in2(_gnd_net_),
            .in3(N__24527),
            .lcout(\current_shift_inst.un4_control_input1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_10_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_10_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_10_18_3  (
            .in0(_gnd_net_),
            .in1(N__24524),
            .in2(_gnd_net_),
            .in3(N__24512),
            .lcout(\current_shift_inst.un4_control_input1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_10_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_10_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_10_18_4  (
            .in0(_gnd_net_),
            .in1(N__24509),
            .in2(_gnd_net_),
            .in3(N__24470),
            .lcout(\current_shift_inst.un4_control_input1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_10_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_10_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_10_18_5  (
            .in0(_gnd_net_),
            .in1(N__24467),
            .in2(_gnd_net_),
            .in3(N__24455),
            .lcout(\current_shift_inst.un4_control_input1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_10_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_10_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_10_18_6  (
            .in0(_gnd_net_),
            .in1(N__24452),
            .in2(_gnd_net_),
            .in3(N__24443),
            .lcout(\current_shift_inst.un4_control_input1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_10_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_10_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_10_18_7  (
            .in0(_gnd_net_),
            .in1(N__24719),
            .in2(_gnd_net_),
            .in3(N__24710),
            .lcout(\current_shift_inst.un4_control_input1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_10_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_10_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_10_19_0  (
            .in0(_gnd_net_),
            .in1(N__24707),
            .in2(_gnd_net_),
            .in3(N__24674),
            .lcout(\current_shift_inst.un4_control_input1_10 ),
            .ltout(),
            .carryin(bfn_10_19_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_10_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_10_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_10_19_1  (
            .in0(_gnd_net_),
            .in1(N__24671),
            .in2(_gnd_net_),
            .in3(N__24662),
            .lcout(\current_shift_inst.un4_control_input1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_10_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_10_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_10_19_2  (
            .in0(_gnd_net_),
            .in1(N__26495),
            .in2(_gnd_net_),
            .in3(N__24659),
            .lcout(\current_shift_inst.un4_control_input1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_10_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_10_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(N__24656),
            .in2(_gnd_net_),
            .in3(N__24647),
            .lcout(\current_shift_inst.un4_control_input1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_10_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_10_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_10_19_4  (
            .in0(_gnd_net_),
            .in1(N__24644),
            .in2(_gnd_net_),
            .in3(N__24635),
            .lcout(\current_shift_inst.un4_control_input1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_10_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_10_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_10_19_5  (
            .in0(_gnd_net_),
            .in1(N__26489),
            .in2(_gnd_net_),
            .in3(N__24632),
            .lcout(\current_shift_inst.un4_control_input1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_10_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_10_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_10_19_6  (
            .in0(_gnd_net_),
            .in1(N__24629),
            .in2(_gnd_net_),
            .in3(N__24602),
            .lcout(\current_shift_inst.un4_control_input1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_10_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_10_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_10_19_7  (
            .in0(_gnd_net_),
            .in1(N__24599),
            .in2(_gnd_net_),
            .in3(N__24590),
            .lcout(\current_shift_inst.un4_control_input1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_10_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_10_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_10_20_0  (
            .in0(_gnd_net_),
            .in1(N__24833),
            .in2(_gnd_net_),
            .in3(N__24827),
            .lcout(\current_shift_inst.un4_control_input1_18 ),
            .ltout(),
            .carryin(bfn_10_20_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_10_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_10_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_10_20_1  (
            .in0(_gnd_net_),
            .in1(N__24845),
            .in2(_gnd_net_),
            .in3(N__24824),
            .lcout(\current_shift_inst.un4_control_input1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_10_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_10_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_10_20_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_10_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24821),
            .in3(N__24809),
            .lcout(\current_shift_inst.un4_control_input1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_10_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_10_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_10_20_3  (
            .in0(_gnd_net_),
            .in1(N__24806),
            .in2(_gnd_net_),
            .in3(N__24800),
            .lcout(\current_shift_inst.un4_control_input1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_10_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_10_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_10_20_4  (
            .in0(_gnd_net_),
            .in1(N__24797),
            .in2(_gnd_net_),
            .in3(N__24758),
            .lcout(\current_shift_inst.un4_control_input1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_10_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_10_20_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_10_20_5  (
            .in0(_gnd_net_),
            .in1(N__24755),
            .in2(_gnd_net_),
            .in3(N__24743),
            .lcout(\current_shift_inst.un4_control_input1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_10_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_10_20_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_10_20_6  (
            .in0(_gnd_net_),
            .in1(N__24740),
            .in2(_gnd_net_),
            .in3(N__24731),
            .lcout(\current_shift_inst.un4_control_input1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_10_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_10_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_10_20_7  (
            .in0(_gnd_net_),
            .in1(N__24728),
            .in2(_gnd_net_),
            .in3(N__24722),
            .lcout(\current_shift_inst.un4_control_input1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_10_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_10_21_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_10_21_0  (
            .in0(_gnd_net_),
            .in1(N__24890),
            .in2(_gnd_net_),
            .in3(N__24884),
            .lcout(\current_shift_inst.un4_control_input1_26 ),
            .ltout(),
            .carryin(bfn_10_21_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_10_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_10_21_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_10_21_1  (
            .in0(_gnd_net_),
            .in1(N__24959),
            .in2(_gnd_net_),
            .in3(N__24881),
            .lcout(\current_shift_inst.un4_control_input1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_10_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_10_21_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_10_21_2  (
            .in0(_gnd_net_),
            .in1(N__24839),
            .in2(_gnd_net_),
            .in3(N__24878),
            .lcout(\current_shift_inst.un4_control_input1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_10_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_10_21_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_10_21_3  (
            .in0(_gnd_net_),
            .in1(N__24875),
            .in2(_gnd_net_),
            .in3(N__24869),
            .lcout(\current_shift_inst.un4_control_input1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_10_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_10_21_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_10_21_4  (
            .in0(_gnd_net_),
            .in1(N__24866),
            .in2(_gnd_net_),
            .in3(N__24854),
            .lcout(\current_shift_inst.un4_control_input1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_10_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_10_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_10_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24851),
            .lcout(\current_shift_inst.un4_control_input1_31_THRU_CO ),
            .ltout(\current_shift_inst.un4_control_input1_31_THRU_CO_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_10_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_10_21_6 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_10_21_6  (
            .in0(N__33548),
            .in1(N__33292),
            .in2(N__24848),
            .in3(N__31982),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_10_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_10_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_10_21_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_10_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30005),
            .lcout(\current_shift_inst.un4_control_input_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_10_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_10_22_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_10_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33848),
            .lcout(\current_shift_inst.un4_control_input_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_10_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_10_22_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_10_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26642),
            .lcout(\current_shift_inst.un4_control_input_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_11_4_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_11_4_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_11_4_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_27_LC_11_4_1  (
            .in0(N__28178),
            .in1(N__28126),
            .in2(_gnd_net_),
            .in3(N__41897),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48788),
            .ce(N__36596),
            .sr(N__48131));
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_11_4_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_11_4_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_11_4_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_17_LC_11_4_7  (
            .in0(N__25123),
            .in1(N__25172),
            .in2(_gnd_net_),
            .in3(N__41896),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48788),
            .ce(N__36596),
            .sr(N__48131));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_11_5_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_11_5_0 .LUT_INIT=16'b0010101100100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_11_5_0  (
            .in0(N__24952),
            .in1(N__27931),
            .in2(N__27677),
            .in3(N__27341),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_11_5_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_11_5_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_11_5_1  (
            .in0(N__27340),
            .in1(N__27676),
            .in2(N__27932),
            .in3(N__24953),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_11_5_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_11_5_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_11_5_4  (
            .in0(N__41781),
            .in1(N__28534),
            .in2(_gnd_net_),
            .in3(N__28592),
            .lcout(elapsed_time_ns_1_RNI47DN9_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_11_5_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_11_5_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_11_5_5  (
            .in0(N__24922),
            .in1(N__41780),
            .in2(_gnd_net_),
            .in3(N__24937),
            .lcout(elapsed_time_ns_1_RNII43T9_0_6),
            .ltout(elapsed_time_ns_1_RNII43T9_0_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_11_5_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_11_5_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_11_5_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_LC_11_5_6  (
            .in0(N__41782),
            .in1(_gnd_net_),
            .in2(N__24926),
            .in3(N__24923),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48781),
            .ce(N__36607),
            .sr(N__48136));
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_0_30_LC_11_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_0_30_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_0_30_LC_11_6_0 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_RNIO0241_0_30_LC_11_6_0  (
            .in0(N__27897),
            .in1(N__25035),
            .in2(N__27871),
            .in3(N__25020),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_11_6_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_11_6_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_11_6_1  (
            .in0(N__41769),
            .in1(N__28174),
            .in2(_gnd_net_),
            .in3(N__28125),
            .lcout(elapsed_time_ns_1_RNI58DN9_0_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_11_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_11_6_3 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_11_6_3  (
            .in0(N__25037),
            .in1(N__27870),
            .in2(N__25025),
            .in3(N__27899),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_11_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_11_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_11_6_4  (
            .in0(N__25122),
            .in1(N__25164),
            .in2(_gnd_net_),
            .in3(N__41768),
            .lcout(elapsed_time_ns_1_RNI46CN9_0_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_11_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_11_6_5 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_11_6_5  (
            .in0(N__41770),
            .in1(N__25057),
            .in2(N__25103),
            .in3(_gnd_net_),
            .lcout(elapsed_time_ns_1_RNIJ53T9_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_30_LC_11_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_30_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_30_LC_11_6_6 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_RNIO0241_30_LC_11_6_6  (
            .in0(N__27898),
            .in1(N__25036),
            .in2(N__27872),
            .in3(N__25021),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un4_running_df30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI4E6P2_28_LC_11_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI4E6P2_28_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI4E6P2_28_LC_11_6_7 .LUT_INIT=16'b1111110101011101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI4E6P2_28_LC_11_6_7  (
            .in0(N__42355),
            .in1(N__25459),
            .in2(N__25010),
            .in3(N__25448),
            .lcout(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_11_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_11_7_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_11_7_0  (
            .in0(N__27814),
            .in1(N__25007),
            .in2(N__25001),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_11_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_11_7_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_11_7_1  (
            .in0(N__27529),
            .in1(N__24992),
            .in2(N__24986),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_11_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_11_7_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_11_7_2  (
            .in0(N__27502),
            .in1(N__24974),
            .in2(N__24968),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_11_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_11_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(N__25307),
            .in2(N__25301),
            .in3(N__27487),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_11_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_11_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_11_7_4  (
            .in0(_gnd_net_),
            .in1(N__25283),
            .in2(N__25292),
            .in3(N__27472),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_11_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_11_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(N__25277),
            .in2(N__25268),
            .in3(N__27457),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_11_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_11_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_11_7_6  (
            .in0(_gnd_net_),
            .in1(N__25259),
            .in2(N__25250),
            .in3(N__27442),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_11_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_11_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_11_7_7  (
            .in0(_gnd_net_),
            .in1(N__25229),
            .in2(N__25241),
            .in3(N__27427),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_11_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_11_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(N__25223),
            .in2(N__25217),
            .in3(N__27412),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_11_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_11_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__25208),
            .in2(N__25202),
            .in3(N__27649),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_11_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_11_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(N__25193),
            .in2(N__25184),
            .in3(N__27634),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_11_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_11_8_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_11_8_3  (
            .in0(N__27619),
            .in1(N__25400),
            .in2(N__25388),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_11_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_11_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__25376),
            .in2(N__25364),
            .in3(N__27604),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_11_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_11_8_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_11_8_5  (
            .in0(N__27589),
            .in1(N__27353),
            .in2(N__25355),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_11_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_11_8_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_11_8_6  (
            .in0(N__27574),
            .in1(N__25331),
            .in2(N__25346),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_11_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_11_8_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(N__30782),
            .in2(N__31142),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_11_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_11_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__25322),
            .in2(N__25316),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_11_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_11_9_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__31457),
            .in2(N__31409),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_11_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_11_9_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__31625),
            .in2(N__31028),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_11_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_11_9_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__25523),
            .in2(N__25511),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_11_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_11_9_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__25502),
            .in2(N__25493),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_11_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_11_9_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(N__25433),
            .in2(N__31247),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_11_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_11_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(N__25478),
            .in2(N__25469),
            .in3(N__25439),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_11_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_11_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25436),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_11_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_11_10_4 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_11_10_4  (
            .in0(N__31859),
            .in1(N__31303),
            .in2(N__31285),
            .in3(N__31264),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_11_10_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_11_10_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_11_10_6  (
            .in0(N__41784),
            .in1(N__28701),
            .in2(_gnd_net_),
            .in3(N__28745),
            .lcout(elapsed_time_ns_1_RNIV0CN9_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_11_10_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_11_10_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_11_10_7  (
            .in0(N__28666),
            .in1(N__28641),
            .in2(_gnd_net_),
            .in3(N__41785),
            .lcout(elapsed_time_ns_1_RNI36DN9_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_11_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_11_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__25427),
            .in2(N__25421),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_11_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_11_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_11_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_11_11_1  (
            .in0(N__26153),
            .in1(N__25681),
            .in2(_gnd_net_),
            .in3(N__25667),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__48717),
            .ce(),
            .sr(N__48185));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_11_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_11_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_11_11_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_11_11_2  (
            .in0(N__26196),
            .in1(N__25654),
            .in2(N__25664),
            .in3(N__25640),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__48717),
            .ce(),
            .sr(N__48185));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_11_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_11_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_11_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_11_11_3  (
            .in0(N__26154),
            .in1(N__25633),
            .in2(_gnd_net_),
            .in3(N__25619),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__48717),
            .ce(),
            .sr(N__48185));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_11_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_11_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_11_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_11_11_4  (
            .in0(N__26197),
            .in1(N__25615),
            .in2(_gnd_net_),
            .in3(N__25601),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__48717),
            .ce(),
            .sr(N__48185));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_11_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_11_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_11_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_11_11_5  (
            .in0(N__26155),
            .in1(N__25597),
            .in2(_gnd_net_),
            .in3(N__25583),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__48717),
            .ce(),
            .sr(N__48185));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_11_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_11_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_11_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_11_11_6  (
            .in0(N__26198),
            .in1(N__25576),
            .in2(_gnd_net_),
            .in3(N__25562),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__48717),
            .ce(),
            .sr(N__48185));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_11_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_11_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_11_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_11_11_7  (
            .in0(N__26156),
            .in1(N__25558),
            .in2(_gnd_net_),
            .in3(N__25544),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__48717),
            .ce(),
            .sr(N__48185));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_11_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_11_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_11_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_11_12_0  (
            .in0(N__26202),
            .in1(N__25540),
            .in2(_gnd_net_),
            .in3(N__25526),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_11_12_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__48707),
            .ce(),
            .sr(N__48195));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_11_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_11_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_11_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_11_12_1  (
            .in0(N__26192),
            .in1(N__25825),
            .in2(_gnd_net_),
            .in3(N__25811),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__48707),
            .ce(),
            .sr(N__48195));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_11_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_11_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_11_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_11_12_2  (
            .in0(N__26199),
            .in1(N__25807),
            .in2(_gnd_net_),
            .in3(N__25793),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__48707),
            .ce(),
            .sr(N__48195));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_11_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_11_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_11_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_11_12_3  (
            .in0(N__26193),
            .in1(N__25789),
            .in2(_gnd_net_),
            .in3(N__25775),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__48707),
            .ce(),
            .sr(N__48195));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_11_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_11_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_11_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_11_12_4  (
            .in0(N__26200),
            .in1(N__25771),
            .in2(_gnd_net_),
            .in3(N__25757),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__48707),
            .ce(),
            .sr(N__48195));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_11_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_11_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_11_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_11_12_5  (
            .in0(N__26194),
            .in1(N__25753),
            .in2(_gnd_net_),
            .in3(N__25739),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__48707),
            .ce(),
            .sr(N__48195));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_11_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_11_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_11_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_11_12_6  (
            .in0(N__26201),
            .in1(N__25735),
            .in2(_gnd_net_),
            .in3(N__25721),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__48707),
            .ce(),
            .sr(N__48195));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_11_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_11_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_11_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_11_12_7  (
            .in0(N__26195),
            .in1(N__25718),
            .in2(_gnd_net_),
            .in3(N__25703),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__48707),
            .ce(),
            .sr(N__48195));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_11_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_11_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_11_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_11_13_0  (
            .in0(N__26145),
            .in1(N__25700),
            .in2(_gnd_net_),
            .in3(N__25685),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__48698),
            .ce(),
            .sr(N__48204));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_11_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_11_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_11_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_11_13_1  (
            .in0(N__26157),
            .in1(N__25983),
            .in2(_gnd_net_),
            .in3(N__25967),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__48698),
            .ce(),
            .sr(N__48204));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_11_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_11_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_11_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_11_13_2  (
            .in0(N__26146),
            .in1(N__25956),
            .in2(_gnd_net_),
            .in3(N__25940),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(N__48698),
            .ce(),
            .sr(N__48204));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_11_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_11_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_11_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_11_13_3  (
            .in0(N__26158),
            .in1(N__25930),
            .in2(_gnd_net_),
            .in3(N__25916),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(N__48698),
            .ce(),
            .sr(N__48204));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_11_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_11_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_11_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_11_13_4  (
            .in0(N__26147),
            .in1(N__25903),
            .in2(_gnd_net_),
            .in3(N__25889),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ),
            .clk(N__48698),
            .ce(),
            .sr(N__48204));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_11_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_11_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_11_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_11_13_5  (
            .in0(N__26159),
            .in1(N__25876),
            .in2(_gnd_net_),
            .in3(N__25862),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ),
            .clk(N__48698),
            .ce(),
            .sr(N__48204));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_11_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_11_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_11_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_11_13_6  (
            .in0(N__26148),
            .in1(N__25852),
            .in2(_gnd_net_),
            .in3(N__25838),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ),
            .clk(N__48698),
            .ce(),
            .sr(N__48204));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_11_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_11_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_11_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_11_13_7  (
            .in0(N__26160),
            .in1(N__27989),
            .in2(_gnd_net_),
            .in3(N__25835),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ),
            .clk(N__48698),
            .ce(),
            .sr(N__48204));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_11_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_11_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_11_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_11_14_0  (
            .in0(N__26149),
            .in1(N__27969),
            .in2(_gnd_net_),
            .in3(N__25832),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ),
            .clk(N__48690),
            .ce(),
            .sr(N__48211));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_11_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_11_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_11_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_11_14_1  (
            .in0(N__26142),
            .in1(N__28422),
            .in2(_gnd_net_),
            .in3(N__25829),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ),
            .clk(N__48690),
            .ce(),
            .sr(N__48211));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_11_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_11_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_11_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_11_14_2  (
            .in0(N__26150),
            .in1(N__28450),
            .in2(_gnd_net_),
            .in3(N__26246),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ),
            .clk(N__48690),
            .ce(),
            .sr(N__48211));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_11_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_11_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_11_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_11_14_3  (
            .in0(N__26143),
            .in1(N__28042),
            .in2(_gnd_net_),
            .in3(N__26243),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ),
            .clk(N__48690),
            .ce(),
            .sr(N__48211));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_11_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_11_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_11_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_11_14_4  (
            .in0(N__26151),
            .in1(N__28089),
            .in2(_gnd_net_),
            .in3(N__26240),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ),
            .clk(N__48690),
            .ce(),
            .sr(N__48211));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_11_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_11_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_11_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_11_14_5  (
            .in0(N__26144),
            .in1(N__26221),
            .in2(_gnd_net_),
            .in3(N__26207),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ),
            .clk(N__48690),
            .ce(),
            .sr(N__48211));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_11_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_11_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_11_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_11_14_6  (
            .in0(N__26152),
            .in1(N__26032),
            .in2(_gnd_net_),
            .in3(N__26048),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48690),
            .ce(),
            .sr(N__48211));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_11_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_11_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__28366),
            .in2(N__29447),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_11_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_11_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__28326),
            .in2(N__26018),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_11_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_11_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(N__32612),
            .in2(N__33121),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_11_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_11_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__32916),
            .in2(N__26006),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_11_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_11_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__26300),
            .in2(N__33122),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_11_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_11_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(N__32920),
            .in2(N__26294),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_11_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_11_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(N__26285),
            .in2(N__33123),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_11_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_11_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(N__32924),
            .in2(N__26279),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_11_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_11_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_LC_11_16_0  (
            .in0(_gnd_net_),
            .in1(N__26270),
            .in2(N__33124),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_16_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_11_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_11_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(N__32928),
            .in2(N__26264),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_11_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_11_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(N__26471),
            .in2(N__33125),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_11_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_11_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_LC_11_16_3  (
            .in0(_gnd_net_),
            .in1(N__32932),
            .in2(N__26255),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_11_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_11_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(N__26342),
            .in2(N__33126),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_11_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_11_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(N__32936),
            .in2(N__32084),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_11_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_11_16_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__32165),
            .in2(N__33127),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_11_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_11_16_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_LC_11_16_7  (
            .in0(_gnd_net_),
            .in1(N__32940),
            .in2(N__26336),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_11_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_11_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_LC_11_17_0  (
            .in0(_gnd_net_),
            .in1(N__26729),
            .in2(N__33259),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_11_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_11_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(N__33135),
            .in2(N__29825),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_11_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_11_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(N__26720),
            .in2(N__33260),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_11_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_11_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(N__33139),
            .in2(N__26327),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_11_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_11_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(N__26711),
            .in2(N__33261),
            .in3(N__26303),
            .lcout(\current_shift_inst.un38_control_input_0_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_11_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_11_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(N__33143),
            .in2(N__26462),
            .in3(N__26438),
            .lcout(\current_shift_inst.un38_control_input_0_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_11_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_11_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(N__26738),
            .in2(N__33262),
            .in3(N__26423),
            .lcout(\current_shift_inst.un38_control_input_0_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_11_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_11_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(N__33147),
            .in2(N__26507),
            .in3(N__26408),
            .lcout(\current_shift_inst.un38_control_input_0_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_11_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_11_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(N__33148),
            .in2(N__26483),
            .in3(N__26393),
            .lcout(\current_shift_inst.un38_control_input_0_s1_24 ),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_11_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_11_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(N__27137),
            .in2(N__33263),
            .in3(N__26378),
            .lcout(\current_shift_inst.un38_control_input_0_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_11_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_11_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(N__33152),
            .in2(N__27203),
            .in3(N__26363),
            .lcout(\current_shift_inst.un38_control_input_0_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_11_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_11_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(N__33788),
            .in2(N__33264),
            .in3(N__26348),
            .lcout(\current_shift_inst.un38_control_input_0_s1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_11_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_11_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(N__33156),
            .in2(N__26672),
            .in3(N__26345),
            .lcout(\current_shift_inst.un38_control_input_0_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_11_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_11_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(N__26843),
            .in2(N__33265),
            .in3(N__26591),
            .lcout(\current_shift_inst.un38_control_input_0_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_11_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_11_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(N__33160),
            .in2(N__26588),
            .in3(N__26573),
            .lcout(\current_shift_inst.un38_control_input_0_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_11_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_11_18_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_11_18_7  (
            .in0(N__33161),
            .in1(N__33492),
            .in2(_gnd_net_),
            .in3(N__26570),
            .lcout(\current_shift_inst.un38_control_input_0_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_11_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_11_19_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_11_19_0  (
            .in0(N__33186),
            .in1(N__33567),
            .in2(N__26567),
            .in3(N__26527),
            .lcout(\current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_11_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_11_19_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_11_19_1  (
            .in0(N__33571),
            .in1(N__33180),
            .in2(N__30073),
            .in3(N__30094),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_11_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_11_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30491),
            .lcout(\current_shift_inst.un4_control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_11_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_11_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32234),
            .lcout(\current_shift_inst.un4_control_input_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_11_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_11_19_4 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_11_19_4  (
            .in0(N__27011),
            .in1(N__33572),
            .in2(N__33270),
            .in3(N__27055),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_11_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_11_19_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_11_19_5  (
            .in0(N__33568),
            .in1(N__33184),
            .in2(N__30416),
            .in3(N__30370),
            .lcout(\current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_11_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_11_19_6 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_11_19_6  (
            .in0(N__33179),
            .in1(N__33570),
            .in2(N__30337),
            .in3(N__30311),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_11_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_11_19_7 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_11_19_7  (
            .in0(N__33569),
            .in1(N__33185),
            .in2(N__29488),
            .in3(N__29533),
            .lcout(\current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_11_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_11_20_0 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_11_20_0  (
            .in0(N__33590),
            .in1(N__29965),
            .in2(N__33271),
            .in3(N__30006),
            .lcout(\current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_11_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_11_20_1 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_11_20_1  (
            .in0(N__30130),
            .in1(N__33591),
            .in2(N__33293),
            .in3(N__30169),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_11_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_11_20_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_11_20_2  (
            .in0(N__30303),
            .in1(N__26988),
            .in2(_gnd_net_),
            .in3(N__30327),
            .lcout(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_11_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_11_20_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_11_20_3  (
            .in0(N__26987),
            .in1(N__30168),
            .in2(_gnd_net_),
            .in3(N__30126),
            .lcout(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_11_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_11_20_4 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_11_20_4  (
            .in0(N__33594),
            .in1(N__27128),
            .in2(N__27085),
            .in3(N__33281),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_11_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_11_20_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_11_20_5  (
            .in0(N__26986),
            .in1(N__30249),
            .in2(_gnd_net_),
            .in3(N__30195),
            .lcout(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_11_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_11_20_6 .LUT_INIT=16'b1000110110001101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_11_20_6  (
            .in0(N__33592),
            .in1(N__26605),
            .in2(N__26648),
            .in3(N__33285),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_11_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_11_20_7 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_11_20_7  (
            .in0(N__26647),
            .in1(N__33593),
            .in2(N__26609),
            .in3(N__33187),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_11_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_11_21_0 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_11_21_0  (
            .in0(N__33290),
            .in1(N__33596),
            .in2(N__27158),
            .in3(N__27190),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_11_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_11_21_1 .LUT_INIT=16'b1111010100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_11_21_1  (
            .in0(N__27191),
            .in1(N__33291),
            .in2(N__33616),
            .in3(N__27154),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_11_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_11_21_2 .LUT_INIT=16'b1111000000110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_11_21_2  (
            .in0(N__33287),
            .in1(N__27127),
            .in2(N__27084),
            .in3(N__33602),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_11_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_11_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_11_21_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_11_21_3  (
            .in0(N__33595),
            .in1(N__33289),
            .in2(N__27056),
            .in3(N__27010),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_11_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_11_21_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_11_21_4  (
            .in0(N__26992),
            .in1(N__32460),
            .in2(_gnd_net_),
            .in3(N__32499),
            .lcout(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_11_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_11_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_11_21_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_11_21_6  (
            .in0(N__33286),
            .in1(N__33600),
            .in2(N__33859),
            .in3(N__33810),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_11_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_11_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_11_21_7 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_11_21_7  (
            .in0(N__33601),
            .in1(N__30580),
            .in2(N__30539),
            .in3(N__33288),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_11_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_11_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_11_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_14_LC_11_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26818),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48656),
            .ce(),
            .sr(N__48258));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_11_23_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_11_23_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_11_23_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_11_23_0  (
            .in0(N__34337),
            .in1(N__27257),
            .in2(N__31004),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_11_23_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_11_23_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_11_23_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_11_23_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_11_23_1  (
            .in0(_gnd_net_),
            .in1(N__27251),
            .in2(N__31013),
            .in3(N__34271),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_11_23_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_11_23_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_11_23_2  (
            .in0(N__34313),
            .in1(N__27245),
            .in2(N__30992),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_11_23_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_11_23_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_11_23_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_11_23_3  (
            .in0(_gnd_net_),
            .in1(N__27239),
            .in2(N__30656),
            .in3(N__34247),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_11_23_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_11_23_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_11_23_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_11_23_4  (
            .in0(_gnd_net_),
            .in1(N__27233),
            .in2(N__30647),
            .in3(N__34292),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_11_23_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_11_23_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_11_23_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_11_23_5  (
            .in0(N__34004),
            .in1(N__27227),
            .in2(N__30638),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_11_23_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_11_23_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_11_23_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_11_23_6  (
            .in0(_gnd_net_),
            .in1(N__27221),
            .in2(N__30629),
            .in3(N__34025),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_11_23_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_11_23_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_11_23_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_11_23_7  (
            .in0(N__34046),
            .in1(N__27215),
            .in2(N__30617),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_11_24_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_11_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_11_24_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_11_24_0  (
            .in0(N__34067),
            .in1(N__27209),
            .in2(N__30983),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_11_24_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_11_24_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_11_24_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_11_24_1  (
            .in0(_gnd_net_),
            .in1(N__27398),
            .in2(N__30806),
            .in3(N__34088),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_11_24_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_11_24_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_11_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_11_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27392),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48650),
            .ce(),
            .sr(N__48267));
    defparam \phase_controller_inst2.S1_LC_11_27_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.S1_LC_11_27_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S1_LC_11_27_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S1_LC_11_27_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31085),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48646),
            .ce(),
            .sr(N__48280));
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_12_4_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_12_4_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_12_4_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_14_LC_12_4_1  (
            .in0(N__30714),
            .in1(N__30770),
            .in2(_gnd_net_),
            .in3(N__41893),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48779),
            .ce(N__36593),
            .sr(N__48127));
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_12_4_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_12_4_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_12_4_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_26_LC_12_4_6  (
            .in0(N__41892),
            .in1(N__28530),
            .in2(_gnd_net_),
            .in3(N__28591),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48779),
            .ce(N__36593),
            .sr(N__48127));
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_12_4_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_12_4_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_12_4_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_16_LC_12_4_7  (
            .in0(N__27332),
            .in1(N__27305),
            .in2(_gnd_net_),
            .in3(N__41894),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48779),
            .ce(N__36593),
            .sr(N__48127));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_12_5_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_12_5_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_12_5_4  (
            .in0(_gnd_net_),
            .in1(N__35075),
            .in2(_gnd_net_),
            .in3(N__27834),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3_28_LC_12_5_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3_28_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3_28_LC_12_5_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3_28_LC_12_5_5  (
            .in0(N__35076),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27835),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_12_6_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_12_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_12_6_0  (
            .in0(_gnd_net_),
            .in1(N__27818),
            .in2(N__27266),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_6_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_12_6_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_12_6_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_12_6_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_12_6_1  (
            .in0(N__36542),
            .in1(N__27530),
            .in2(_gnd_net_),
            .in3(N__27518),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__48761),
            .ce(),
            .sr(N__48137));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_12_6_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_12_6_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_12_6_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_12_6_2  (
            .in0(N__36546),
            .in1(N__27503),
            .in2(N__27515),
            .in3(N__27491),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__48761),
            .ce(),
            .sr(N__48137));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_12_6_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_12_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_12_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_12_6_3  (
            .in0(N__36543),
            .in1(N__27488),
            .in2(_gnd_net_),
            .in3(N__27476),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__48761),
            .ce(),
            .sr(N__48137));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_12_6_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_12_6_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_12_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_12_6_4  (
            .in0(N__36547),
            .in1(N__27473),
            .in2(_gnd_net_),
            .in3(N__27461),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__48761),
            .ce(),
            .sr(N__48137));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_12_6_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_12_6_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_12_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_12_6_5  (
            .in0(N__36544),
            .in1(N__27458),
            .in2(_gnd_net_),
            .in3(N__27446),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__48761),
            .ce(),
            .sr(N__48137));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_12_6_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_12_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_12_6_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_12_6_6  (
            .in0(N__36548),
            .in1(N__27443),
            .in2(_gnd_net_),
            .in3(N__27431),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__48761),
            .ce(),
            .sr(N__48137));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_12_6_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_12_6_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_12_6_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_12_6_7  (
            .in0(N__36545),
            .in1(N__27428),
            .in2(_gnd_net_),
            .in3(N__27416),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__48761),
            .ce(),
            .sr(N__48137));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_12_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_12_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_12_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_12_7_0  (
            .in0(N__36573),
            .in1(N__27413),
            .in2(_gnd_net_),
            .in3(N__27401),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_12_7_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__48747),
            .ce(),
            .sr(N__48142));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_12_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_12_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_12_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_12_7_1  (
            .in0(N__36558),
            .in1(N__27650),
            .in2(_gnd_net_),
            .in3(N__27638),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__48747),
            .ce(),
            .sr(N__48142));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_12_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_12_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_12_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_12_7_2  (
            .in0(N__36570),
            .in1(N__27635),
            .in2(_gnd_net_),
            .in3(N__27623),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__48747),
            .ce(),
            .sr(N__48142));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_12_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_12_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_12_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_12_7_3  (
            .in0(N__36559),
            .in1(N__27620),
            .in2(_gnd_net_),
            .in3(N__27608),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__48747),
            .ce(),
            .sr(N__48142));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_12_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_12_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_12_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_12_7_4  (
            .in0(N__36571),
            .in1(N__27605),
            .in2(_gnd_net_),
            .in3(N__27593),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__48747),
            .ce(),
            .sr(N__48142));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_12_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_12_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_12_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_12_7_5  (
            .in0(N__36560),
            .in1(N__27590),
            .in2(_gnd_net_),
            .in3(N__27578),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__48747),
            .ce(),
            .sr(N__48142));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_12_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_12_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_12_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_12_7_6  (
            .in0(N__36572),
            .in1(N__27575),
            .in2(_gnd_net_),
            .in3(N__27563),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__48747),
            .ce(),
            .sr(N__48142));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_12_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_12_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_12_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_12_7_7  (
            .in0(N__36561),
            .in1(N__31164),
            .in2(_gnd_net_),
            .in3(N__27560),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__48747),
            .ce(),
            .sr(N__48142));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_12_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_12_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_12_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_12_8_0  (
            .in0(N__36562),
            .in1(N__31218),
            .in2(_gnd_net_),
            .in3(N__27557),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_12_8_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__48735),
            .ce(),
            .sr(N__48151));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_12_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_12_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_12_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_12_8_1  (
            .in0(N__36577),
            .in1(N__27549),
            .in2(_gnd_net_),
            .in3(N__27533),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__48735),
            .ce(),
            .sr(N__48151));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_12_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_12_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_12_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_12_8_2  (
            .in0(N__36563),
            .in1(N__27774),
            .in2(_gnd_net_),
            .in3(N__27758),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(N__48735),
            .ce(),
            .sr(N__48151));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_12_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_12_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_12_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_12_8_3  (
            .in0(N__36578),
            .in1(N__31425),
            .in2(_gnd_net_),
            .in3(N__27755),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(N__48735),
            .ce(),
            .sr(N__48151));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_12_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_12_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_12_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_12_8_4  (
            .in0(N__36564),
            .in1(N__31445),
            .in2(_gnd_net_),
            .in3(N__27752),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ),
            .clk(N__48735),
            .ce(),
            .sr(N__48151));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_12_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_12_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_12_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_12_8_5  (
            .in0(N__36579),
            .in1(N__31660),
            .in2(_gnd_net_),
            .in3(N__27749),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ),
            .clk(N__48735),
            .ce(),
            .sr(N__48151));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_12_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_12_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_12_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_12_8_6  (
            .in0(N__36565),
            .in1(N__31642),
            .in2(_gnd_net_),
            .in3(N__27746),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ),
            .clk(N__48735),
            .ce(),
            .sr(N__48151));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_12_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_12_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_12_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_12_8_7  (
            .in0(N__36580),
            .in1(N__27735),
            .in2(_gnd_net_),
            .in3(N__27713),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ),
            .clk(N__48735),
            .ce(),
            .sr(N__48151));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_12_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_12_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_12_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_12_9_0  (
            .in0(N__36566),
            .in1(N__27702),
            .in2(_gnd_net_),
            .in3(N__27680),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ),
            .clk(N__48725),
            .ce(),
            .sr(N__48159));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_12_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_12_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_12_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_12_9_1  (
            .in0(N__36574),
            .in1(N__27667),
            .in2(_gnd_net_),
            .in3(N__27653),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ),
            .clk(N__48725),
            .ce(),
            .sr(N__48159));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_12_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_12_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_12_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_12_9_2  (
            .in0(N__36567),
            .in1(N__27922),
            .in2(_gnd_net_),
            .in3(N__27908),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ),
            .clk(N__48725),
            .ce(),
            .sr(N__48159));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_12_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_12_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_12_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_12_9_3  (
            .in0(N__36575),
            .in1(N__31265),
            .in2(_gnd_net_),
            .in3(N__27905),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ),
            .clk(N__48725),
            .ce(),
            .sr(N__48159));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_12_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_12_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_12_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_12_9_4  (
            .in0(N__36568),
            .in1(N__31304),
            .in2(_gnd_net_),
            .in3(N__27902),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ),
            .clk(N__48725),
            .ce(),
            .sr(N__48159));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_12_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_12_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_12_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_12_9_5  (
            .in0(N__36576),
            .in1(N__27896),
            .in2(_gnd_net_),
            .in3(N__27878),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ),
            .clk(N__48725),
            .ce(),
            .sr(N__48159));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_12_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_12_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_12_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_12_9_6  (
            .in0(N__36569),
            .in1(N__27856),
            .in2(_gnd_net_),
            .in3(N__27875),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48725),
            .ce(),
            .sr(N__48159));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_12_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_12_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_12_10_1 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_12_10_1  (
            .in0(N__46202),
            .in1(N__42284),
            .in2(N__44733),
            .in3(N__46701),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48715),
            .ce(),
            .sr(N__48167));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_12_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_12_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_12_10_2 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_12_10_2  (
            .in0(N__36469),
            .in1(N__27842),
            .in2(N__35093),
            .in3(N__27813),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48715),
            .ce(),
            .sr(N__48167));
    defparam \phase_controller_inst2.start_timer_hc_LC_12_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_LC_12_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_hc_LC_12_10_3 .LUT_INIT=16'b1100110011001110;
    LogicCell40 \phase_controller_inst2.start_timer_hc_LC_12_10_3  (
            .in0(N__28278),
            .in1(N__31097),
            .in2(N__42968),
            .in3(N__27794),
            .lcout(\phase_controller_inst2.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48715),
            .ce(),
            .sr(N__48167));
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_12_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_12_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_12_10_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_LC_12_10_5  (
            .in0(N__28279),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48715),
            .ce(),
            .sr(N__48167));
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_12_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_12_10_6 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_12_10_6  (
            .in0(N__28196),
            .in1(N__28301),
            .in2(_gnd_net_),
            .in3(N__28277),
            .lcout(\phase_controller_inst2.stoper_hc.un2_start_0 ),
            .ltout(\phase_controller_inst2.stoper_hc.un2_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_12_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_12_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_12_10_7 .LUT_INIT=16'b1011101000001010;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_LC_12_10_7  (
            .in0(N__31800),
            .in1(N__28238),
            .in2(N__28214),
            .in3(N__28197),
            .lcout(\phase_controller_inst2.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48715),
            .ce(),
            .sr(N__48167));
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_12_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_12_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_12_11_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_27_LC_12_11_1  (
            .in0(N__28173),
            .in1(N__28130),
            .in2(_gnd_net_),
            .in3(N__41854),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48705),
            .ce(N__28510),
            .sr(N__48176));
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_12_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_12_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_12_11_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_28_LC_12_11_2  (
            .in0(N__41853),
            .in1(N__31890),
            .in2(_gnd_net_),
            .in3(N__31910),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48705),
            .ce(N__28510),
            .sr(N__48176));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_12_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_12_11_3 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_12_11_3  (
            .in0(N__28027),
            .in1(N__28090),
            .in2(N__28073),
            .in3(N__28051),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_12_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_12_11_4 .LUT_INIT=16'b0100110101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_12_11_4  (
            .in0(N__28091),
            .in1(N__28069),
            .in2(N__28052),
            .in3(N__28028),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_12_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_12_12_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_12_12_0  (
            .in0(N__27987),
            .in1(N__27970),
            .in2(N__28604),
            .in3(N__27941),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_12_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_12_12_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_12_12_1  (
            .in0(N__27940),
            .in1(N__27988),
            .in2(N__27974),
            .in3(N__28600),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_12_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_12_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_12_12_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_24_LC_12_12_2  (
            .in0(N__38204),
            .in1(N__38256),
            .in2(_gnd_net_),
            .in3(N__41857),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48697),
            .ce(N__28507),
            .sr(N__48186));
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_12_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_12_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_12_12_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_12_LC_12_12_4  (
            .in0(N__28743),
            .in1(N__28705),
            .in2(_gnd_net_),
            .in3(N__41856),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48697),
            .ce(N__28507),
            .sr(N__48186));
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_12_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_12_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_12_12_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_25_LC_12_12_5  (
            .in0(N__41855),
            .in1(N__28667),
            .in2(_gnd_net_),
            .in3(N__28646),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48697),
            .ce(N__28507),
            .sr(N__48186));
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_12_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_12_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_12_12_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_26_LC_12_12_6  (
            .in0(N__28584),
            .in1(N__28538),
            .in2(_gnd_net_),
            .in3(N__41858),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48697),
            .ce(N__28507),
            .sr(N__48186));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_12_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_12_12_7 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_12_12_7  (
            .in0(N__28462),
            .in1(N__28451),
            .in2(N__28430),
            .in3(N__28393),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_12_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_12_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(N__28367),
            .in2(N__33632),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_13_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_12_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_12_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(N__28317),
            .in2(N__28343),
            .in3(N__31983),
            .lcout(\current_shift_inst.un38_control_input_5_1 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_12_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_12_13_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_12_13_2  (
            .in0(N__31984),
            .in1(N__32756),
            .in2(N__29735),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un38_control_input_5_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_12_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_12_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(N__29744),
            .in2(N__32910),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_12_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_12_13_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(N__32760),
            .in2(N__32351),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_12_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_12_13_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(N__28784),
            .in2(N__32911),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_12_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_12_13_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(N__32764),
            .in2(N__29552),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_12_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_12_13_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_LC_12_13_7  (
            .in0(_gnd_net_),
            .in1(N__29648),
            .in2(N__32912),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_12_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_12_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(N__32851),
            .in2(N__28772),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_14_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_12_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_12_14_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(N__28754),
            .in2(N__33065),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_12_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_12_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_LC_12_14_2  (
            .in0(_gnd_net_),
            .in1(N__32855),
            .in2(N__30353),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_12_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_12_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_LC_12_14_3  (
            .in0(_gnd_net_),
            .in1(N__30425),
            .in2(N__33066),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_12_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_12_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_LC_12_14_4  (
            .in0(_gnd_net_),
            .in1(N__32859),
            .in2(N__32267),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_12_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_12_14_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(N__32522),
            .in2(N__33067),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_12_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_12_14_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_LC_12_14_6  (
            .in0(_gnd_net_),
            .in1(N__32863),
            .in2(N__32531),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_12_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_12_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(N__28805),
            .in2(N__33068),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_12_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_12_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(N__32941),
            .in2(N__29462),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_15_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_12_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_12_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(N__32432),
            .in2(N__33128),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_12_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_12_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(N__32945),
            .in2(N__29948),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_12_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_12_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(N__30182),
            .in2(N__33129),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_12_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_12_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(N__32949),
            .in2(N__30110),
            .in3(N__28787),
            .lcout(\current_shift_inst.un38_control_input_0_s0_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_12_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_12_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_12_15_5  (
            .in0(_gnd_net_),
            .in1(N__28991),
            .in2(N__33130),
            .in3(N__28970),
            .lcout(\current_shift_inst.un38_control_input_0_s0_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_12_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_12_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(N__32953),
            .in2(N__30275),
            .in3(N__28958),
            .lcout(\current_shift_inst.un38_control_input_0_s0_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_12_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_12_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(N__30026),
            .in2(N__33131),
            .in3(N__28946),
            .lcout(\current_shift_inst.un38_control_input_0_s0_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_12_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_12_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__33029),
            .in2(N__28943),
            .in3(N__28913),
            .lcout(\current_shift_inst.un38_control_input_0_s0_24 ),
            .ltout(),
            .carryin(bfn_12_16_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_12_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_12_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__28910),
            .in2(N__33191),
            .in3(N__28883),
            .lcout(\current_shift_inst.un38_control_input_0_s0_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_12_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_12_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(N__33033),
            .in2(N__28880),
            .in3(N__28853),
            .lcout(\current_shift_inst.un38_control_input_0_s0_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_12_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_12_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(N__28850),
            .in2(N__33192),
            .in3(N__28826),
            .lcout(\current_shift_inst.un38_control_input_0_s0_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_12_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_12_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_12_16_4  (
            .in0(_gnd_net_),
            .in1(N__33037),
            .in2(N__28823),
            .in3(N__28808),
            .lcout(\current_shift_inst.un38_control_input_0_s0_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_12_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_12_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(N__30509),
            .in2(N__33193),
            .in3(N__29420),
            .lcout(\current_shift_inst.un38_control_input_0_s0_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_12_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_12_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_12_16_6  (
            .in0(_gnd_net_),
            .in1(N__33041),
            .in2(N__32540),
            .in3(N__29417),
            .lcout(\current_shift_inst.un38_control_input_0_s0_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_12_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_12_16_7 .LUT_INIT=16'b1010001101010011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_12_16_7  (
            .in0(N__29414),
            .in1(N__29402),
            .in2(N__29318),
            .in3(N__29393),
            .lcout(\current_shift_inst.control_input_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_12_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_12_17_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_12_17_0  (
            .in0(N__29378),
            .in1(N__29372),
            .in2(_gnd_net_),
            .in3(N__29312),
            .lcout(\current_shift_inst.control_input_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_12_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_12_17_1 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_12_17_1  (
            .in0(N__29313),
            .in1(N__29354),
            .in2(_gnd_net_),
            .in3(N__29348),
            .lcout(\current_shift_inst.control_input_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_12_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_12_17_2 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_12_17_2  (
            .in0(N__29330),
            .in1(N__29324),
            .in2(_gnd_net_),
            .in3(N__29314),
            .lcout(\current_shift_inst.control_input_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_12_17_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_12_17_3 .LUT_INIT=16'b0011111100001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(N__29928),
            .in2(N__29915),
            .in3(N__29158),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_199_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_12_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_12_17_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_12_17_4 .LUT_INIT=16'b0000101011111010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_12_17_4  (
            .in0(N__29159),
            .in1(_gnd_net_),
            .in2(N__29933),
            .in3(N__29914),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48671),
            .ce(),
            .sr(N__48223));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_12_17_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_12_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_12_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29927),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_12_17_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_12_17_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_12_17_6  (
            .in0(N__29929),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29910),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_198_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_12_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_12_18_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_12_18_1  (
            .in0(N__33166),
            .in1(N__33406),
            .in2(N__32482),
            .in3(N__32515),
            .lcout(\current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_12_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_12_18_2 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_12_18_2  (
            .in0(N__33401),
            .in1(N__33167),
            .in2(N__29815),
            .in3(N__29767),
            .lcout(\current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_18_3 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_18_3  (
            .in0(N__32632),
            .in1(N__33400),
            .in2(N__33266),
            .in3(N__32674),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_12_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_12_18_4 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_12_18_4  (
            .in0(N__33404),
            .in1(N__33169),
            .in2(N__29720),
            .in3(N__29692),
            .lcout(\current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_12_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_12_18_5 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_12_18_5  (
            .in0(N__33168),
            .in1(N__33403),
            .in2(N__29635),
            .in3(N__29575),
            .lcout(\current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_12_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_12_18_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_12_18_6  (
            .in0(N__33405),
            .in1(N__33165),
            .in2(N__29537),
            .in3(N__29489),
            .lcout(\current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_12_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_12_18_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_12_18_7  (
            .in0(N__33668),
            .in1(N__33402),
            .in2(_gnd_net_),
            .in3(N__33677),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_12_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_12_19_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_12_19_0  (
            .in0(N__33435),
            .in1(N__30581),
            .in2(N__33267),
            .in3(N__30538),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_12_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_12_19_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_12_19_2  (
            .in0(N__33434),
            .in1(N__30499),
            .in2(N__33269),
            .in3(N__30451),
            .lcout(\current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_12_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_12_19_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_12_19_6  (
            .in0(N__33433),
            .in1(N__30412),
            .in2(N__33268),
            .in3(N__30374),
            .lcout(\current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_12_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_12_20_0 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_12_20_0  (
            .in0(N__33453),
            .in1(N__33114),
            .in2(N__30338),
            .in3(N__30310),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_12_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_12_20_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_12_20_1  (
            .in0(N__33120),
            .in1(N__33451),
            .in2(N__30260),
            .in3(N__30202),
            .lcout(\current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_12_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_12_20_2 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_12_20_2  (
            .in0(N__33452),
            .in1(N__33118),
            .in2(N__30170),
            .in3(N__30131),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_12_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_12_20_3 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_12_20_3  (
            .in0(N__30095),
            .in1(N__33454),
            .in2(N__33258),
            .in3(N__30074),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_12_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_12_20_4 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_12_20_4  (
            .in0(N__33450),
            .in1(N__33119),
            .in2(N__30014),
            .in3(N__29969),
            .lcout(\current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_0_LC_12_21_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_12_21_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_12_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_12_21_0  (
            .in0(N__33971),
            .in1(N__34333),
            .in2(_gnd_net_),
            .in3(N__30608),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_12_21_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__48655),
            .ce(),
            .sr(N__48244));
    defparam \pwm_generator_inst.counter_1_LC_12_21_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_12_21_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_12_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_12_21_1  (
            .in0(N__33965),
            .in1(N__34270),
            .in2(_gnd_net_),
            .in3(N__30605),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__48655),
            .ce(),
            .sr(N__48244));
    defparam \pwm_generator_inst.counter_2_LC_12_21_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_12_21_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_12_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_12_21_2  (
            .in0(N__33972),
            .in1(N__34312),
            .in2(_gnd_net_),
            .in3(N__30602),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__48655),
            .ce(),
            .sr(N__48244));
    defparam \pwm_generator_inst.counter_3_LC_12_21_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_12_21_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_12_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_12_21_3  (
            .in0(N__33966),
            .in1(N__34246),
            .in2(_gnd_net_),
            .in3(N__30599),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__48655),
            .ce(),
            .sr(N__48244));
    defparam \pwm_generator_inst.counter_4_LC_12_21_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_12_21_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_12_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_12_21_4  (
            .in0(N__33973),
            .in1(N__34291),
            .in2(_gnd_net_),
            .in3(N__30596),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__48655),
            .ce(),
            .sr(N__48244));
    defparam \pwm_generator_inst.counter_5_LC_12_21_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_12_21_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_12_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_12_21_5  (
            .in0(N__33967),
            .in1(N__34002),
            .in2(_gnd_net_),
            .in3(N__30593),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__48655),
            .ce(),
            .sr(N__48244));
    defparam \pwm_generator_inst.counter_6_LC_12_21_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_12_21_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_12_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_12_21_6  (
            .in0(N__33974),
            .in1(N__34023),
            .in2(_gnd_net_),
            .in3(N__30590),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__48655),
            .ce(),
            .sr(N__48244));
    defparam \pwm_generator_inst.counter_7_LC_12_21_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_12_21_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_12_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_12_21_7  (
            .in0(N__33968),
            .in1(N__34045),
            .in2(_gnd_net_),
            .in3(N__30587),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__48655),
            .ce(),
            .sr(N__48244));
    defparam \pwm_generator_inst.counter_8_LC_12_22_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_12_22_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_12_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_12_22_0  (
            .in0(N__33970),
            .in1(N__34066),
            .in2(_gnd_net_),
            .in3(N__30584),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_12_22_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__48652),
            .ce(),
            .sr(N__48251));
    defparam \pwm_generator_inst.counter_9_LC_12_22_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_12_22_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_12_22_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \pwm_generator_inst.counter_9_LC_12_22_1  (
            .in0(N__34087),
            .in1(N__33969),
            .in2(_gnd_net_),
            .in3(N__30698),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48652),
            .ce(),
            .sr(N__48251));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_12_23_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_12_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_12_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_12_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48958),
            .lcout(N_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48649),
            .ce(),
            .sr(N__48259));
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_12_23_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_12_23_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_12_23_2  (
            .in0(N__35321),
            .in1(N__30679),
            .in2(_gnd_net_),
            .in3(N__30859),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_12_23_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_12_23_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_12_23_3 .LUT_INIT=16'b1001010101101010;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_12_23_3  (
            .in0(N__30695),
            .in1(N__30680),
            .in2(N__30895),
            .in3(N__35320),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_12_23_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_12_23_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_12_23_7 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_12_23_7  (
            .in0(N__47463),
            .in1(N__47537),
            .in2(N__30896),
            .in3(N__34397),
            .lcout(\pwm_generator_inst.threshold_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_12_24_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_12_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_12_24_0 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_12_24_0  (
            .in0(N__47472),
            .in1(N__47541),
            .in2(N__30899),
            .in3(N__34388),
            .lcout(\pwm_generator_inst.threshold_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_12_24_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_12_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_12_24_1 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_12_24_1  (
            .in0(N__47542),
            .in1(N__47473),
            .in2(N__34379),
            .in3(N__30877),
            .lcout(\pwm_generator_inst.threshold_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_12_24_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_12_24_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_12_24_2 .LUT_INIT=16'b1111111101010011;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_12_24_2  (
            .in0(N__47474),
            .in1(N__47543),
            .in2(N__30898),
            .in3(N__34367),
            .lcout(\pwm_generator_inst.un14_counter_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_12_24_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_12_24_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_12_24_3 .LUT_INIT=16'b1111111100110101;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_12_24_3  (
            .in0(N__47544),
            .in1(N__47475),
            .in2(N__30900),
            .in3(N__34358),
            .lcout(\pwm_generator_inst.un14_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_12_24_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_12_24_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_12_24_5 .LUT_INIT=16'b1111001111110101;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_12_24_5  (
            .in0(N__47539),
            .in1(N__47470),
            .in2(N__34421),
            .in3(N__30869),
            .lcout(\pwm_generator_inst.un14_counter_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_12_24_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_12_24_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_12_24_6 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_12_24_6  (
            .in0(N__47469),
            .in1(N__47538),
            .in2(N__30897),
            .in3(N__33869),
            .lcout(\pwm_generator_inst.threshold_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_12_24_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_12_24_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_12_24_7 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_12_24_7  (
            .in0(N__47540),
            .in1(N__47471),
            .in2(N__34409),
            .in3(N__30870),
            .lcout(\pwm_generator_inst.threshold_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_12_25_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_12_25_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_12_25_1 .LUT_INIT=16'b1111000111111101;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_12_25_1  (
            .in0(N__47545),
            .in1(N__30891),
            .in2(N__34349),
            .in3(N__47477),
            .lcout(\pwm_generator_inst.un14_counter_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_12_25_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_12_25_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_12_25_6 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_12_25_6  (
            .in0(N__47476),
            .in1(N__47546),
            .in2(N__30939),
            .in3(N__34472),
            .lcout(\pwm_generator_inst.threshold_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_26_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_26_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_26_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_26_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_7 .C_ON=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_7 .SEQ_MODE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48308),
            .lcout(\pll_inst.red_c_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_13_4_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_13_4_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_13_4_4 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_13_4_4  (
            .in0(N__31234),
            .in1(N__31223),
            .in2(N__31195),
            .in3(N__31169),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_13_4_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_13_4_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_13_4_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_13_4_5  (
            .in0(N__30718),
            .in1(N__30768),
            .in2(_gnd_net_),
            .in3(N__41889),
            .lcout(elapsed_time_ns_1_RNI13CN9_0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_13_5_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_13_5_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_13_5_0 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_13_5_0  (
            .in0(N__31235),
            .in1(N__31222),
            .in2(N__31196),
            .in3(N__31168),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_0_LC_13_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_0_LC_13_6_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_0_LC_13_6_0 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \phase_controller_inst2.state_0_LC_13_6_0  (
            .in0(N__31733),
            .in1(N__31837),
            .in2(N__31115),
            .in3(N__31127),
            .lcout(\phase_controller_inst2.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48770),
            .ce(),
            .sr(N__48132));
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_13_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_13_6_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_13_6_1 .LUT_INIT=16'b1011000010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_LC_13_6_1  (
            .in0(N__31126),
            .in1(N__35603),
            .in2(N__35237),
            .in3(N__35174),
            .lcout(\phase_controller_inst2.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48770),
            .ce(),
            .sr(N__48132));
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_13_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_13_6_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_13_6_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.state_RNI9M3O_0_LC_13_6_2  (
            .in0(_gnd_net_),
            .in1(N__31125),
            .in2(_gnd_net_),
            .in3(N__31111),
            .lcout(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ),
            .ltout(\phase_controller_inst2.state_RNI9M3OZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_3_LC_13_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_3_LC_13_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_3_LC_13_6_3 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \phase_controller_inst2.state_3_LC_13_6_3  (
            .in0(N__31069),
            .in1(N__31052),
            .in2(N__31100),
            .in3(N__36283),
            .lcout(\phase_controller_inst2.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48770),
            .ce(),
            .sr(N__48132));
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_13_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_13_6_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_13_6_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_RNO_0_LC_13_6_4  (
            .in0(N__31050),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31067),
            .lcout(\phase_controller_inst2.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_13_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_13_6_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_13_6_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.state_ns_i_a3_1_LC_13_6_5  (
            .in0(_gnd_net_),
            .in1(N__43006),
            .in2(_gnd_net_),
            .in3(N__42941),
            .lcout(state_ns_i_a3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_2_LC_13_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_2_LC_13_6_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_2_LC_13_6_7 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \phase_controller_inst2.state_2_LC_13_6_7  (
            .in0(N__31068),
            .in1(N__31051),
            .in2(N__31761),
            .in3(N__31805),
            .lcout(\phase_controller_inst2.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48770),
            .ce(),
            .sr(N__48132));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_13_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_13_7_0 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_13_7_0  (
            .in0(N__31550),
            .in1(N__31466),
            .in2(N__31661),
            .in3(N__31641),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_13_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_13_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_13_7_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_13_7_1  (
            .in0(N__31465),
            .in1(N__31659),
            .in2(N__31643),
            .in3(N__31549),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_13_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_13_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_13_7_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_23_LC_13_7_3  (
            .in0(N__31613),
            .in1(N__31589),
            .in2(_gnd_net_),
            .in3(N__41860),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48762),
            .ce(N__36531),
            .sr(N__48138));
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_13_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_13_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_13_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_22_LC_13_7_5  (
            .in0(N__31541),
            .in1(N__31511),
            .in2(_gnd_net_),
            .in3(N__41859),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48762),
            .ce(N__36531),
            .sr(N__48138));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_13_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_13_8_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_13_8_0  (
            .in0(N__31444),
            .in1(N__31426),
            .in2(N__31394),
            .in3(N__31313),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_13_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_13_8_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_13_8_1  (
            .in0(N__31312),
            .in1(N__31443),
            .in2(N__31430),
            .in3(N__31390),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_13_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_13_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_13_8_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_21_LC_13_8_3  (
            .in0(N__41420),
            .in1(N__41945),
            .in2(_gnd_net_),
            .in3(N__41821),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48749),
            .ce(N__36538),
            .sr(N__48143));
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_13_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_13_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_13_8_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_20_LC_13_8_5  (
            .in0(N__31382),
            .in1(N__31358),
            .in2(_gnd_net_),
            .in3(N__41820),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48749),
            .ce(N__36538),
            .sr(N__48143));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_13_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_13_9_1 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_13_9_1  (
            .in0(N__31852),
            .in1(N__31302),
            .in2(N__31286),
            .in3(N__31263),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_13_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_13_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_13_9_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_13_9_6  (
            .in0(N__31891),
            .in1(N__31906),
            .in2(_gnd_net_),
            .in3(N__41851),
            .lcout(elapsed_time_ns_1_RNI69DN9_0_28),
            .ltout(elapsed_time_ns_1_RNI69DN9_0_28_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_13_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_13_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_13_9_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_28_LC_13_9_7  (
            .in0(N__41852),
            .in1(_gnd_net_),
            .in2(N__31895),
            .in3(N__31892),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48737),
            .ce(N__36594),
            .sr(N__48152));
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_13_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_13_10_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \phase_controller_inst2.start_timer_tr_RNO_0_LC_13_10_0  (
            .in0(N__31841),
            .in1(N__31799),
            .in2(N__31772),
            .in3(N__31731),
            .lcout(),
            .ltout(\phase_controller_inst2.start_timer_tr_RNO_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_tr_LC_13_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_LC_13_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_tr_LC_13_10_1 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \phase_controller_inst2.start_timer_tr_LC_13_10_1  (
            .in0(N__35190),
            .in1(N__31685),
            .in2(N__31676),
            .in3(N__42966),
            .lcout(\phase_controller_inst2.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48727),
            .ce(),
            .sr(N__48160));
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_13_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_13_10_2 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_13_10_2  (
            .in0(N__35216),
            .in1(N__31672),
            .in2(_gnd_net_),
            .in3(N__35189),
            .lcout(\phase_controller_inst2.stoper_tr.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.running_LC_13_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_LC_13_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.running_LC_13_10_3 .LUT_INIT=16'b1000101011111010;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_LC_13_10_3  (
            .in0(N__31673),
            .in1(N__35599),
            .in2(N__35172),
            .in3(N__35218),
            .lcout(\phase_controller_inst2.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48727),
            .ce(),
            .sr(N__48160));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNISIOB3_28_LC_13_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNISIOB3_28_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNISIOB3_28_LC_13_10_4 .LUT_INIT=16'b1111110101110101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNISIOB3_28_LC_13_10_4  (
            .in0(N__35217),
            .in1(N__32033),
            .in2(N__35638),
            .in3(N__35615),
            .lcout(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_13_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_13_10_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_13_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31664),
            .in3(N__35156),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_13_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_13_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_13_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_LC_13_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35191),
            .lcout(\phase_controller_inst2.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48727),
            .ce(),
            .sr(N__48160));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34_28_LC_13_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34_28_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34_28_LC_13_10_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34_28_LC_13_10_7  (
            .in0(_gnd_net_),
            .in1(N__35157),
            .in2(_gnd_net_),
            .in3(N__35131),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_13_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_13_11_0 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_13_11_0  (
            .in0(N__31921),
            .in1(N__31934),
            .in2(N__35885),
            .in3(N__35863),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_13_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_13_11_1 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_13_11_1  (
            .in0(N__31933),
            .in1(N__35862),
            .in2(N__31925),
            .in3(N__35883),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_13_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_13_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_13_11_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_16_LC_13_11_2  (
            .in0(N__42266),
            .in1(N__42170),
            .in2(_gnd_net_),
            .in3(N__47120),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48718),
            .ce(N__46110),
            .sr(N__48168));
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_13_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_13_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_13_11_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_2_LC_13_11_6  (
            .in0(N__43622),
            .in1(N__43592),
            .in2(_gnd_net_),
            .in3(N__47121),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48718),
            .ce(N__46110),
            .sr(N__48168));
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_13_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_13_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_13_12_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_17_LC_13_12_0  (
            .in0(N__47116),
            .in1(N__42224),
            .in2(_gnd_net_),
            .in3(N__42527),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48708),
            .ce(N__46112),
            .sr(N__48177));
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_13_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_13_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_13_12_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_15_LC_13_12_1  (
            .in0(N__43409),
            .in1(N__43383),
            .in2(_gnd_net_),
            .in3(N__47117),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48708),
            .ce(N__46112),
            .sr(N__48177));
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_13_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_13_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_13_12_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_29_LC_13_12_3  (
            .in0(N__42449),
            .in1(N__42425),
            .in2(_gnd_net_),
            .in3(N__47119),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48708),
            .ce(N__46112),
            .sr(N__48177));
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_13_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_13_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_13_12_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_19_LC_13_12_7  (
            .in0(N__44813),
            .in1(N__44787),
            .in2(_gnd_net_),
            .in3(N__47118),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48708),
            .ce(N__46112),
            .sr(N__48177));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_13_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_13_13_0 .LUT_INIT=16'b0100110101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_13_13_0  (
            .in0(N__35958),
            .in1(N__32054),
            .in2(N__35984),
            .in3(N__32042),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_13_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_13_13_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_13_13_1  (
            .in0(N__32041),
            .in1(N__35982),
            .in2(N__35963),
            .in3(N__32053),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_13_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_13_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_13_13_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_28_LC_13_13_2  (
            .in0(N__44232),
            .in1(N__43808),
            .in2(_gnd_net_),
            .in3(N__47122),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48699),
            .ce(N__46113),
            .sr(N__48187));
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_0_30_LC_13_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_0_30_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_0_30_LC_13_14_0 .LUT_INIT=16'b0100111100000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_0_30_LC_13_14_0  (
            .in0(N__36213),
            .in1(N__32023),
            .in2(N__44138),
            .in3(N__36041),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_30_LC_13_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_30_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_30_LC_13_14_1 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_30_LC_13_14_1  (
            .in0(N__32022),
            .in1(N__44136),
            .in2(N__36046),
            .in3(N__36212),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_df30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_13_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_13_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_13_14_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_30_LC_13_14_2  (
            .in0(N__45788),
            .in1(N__45806),
            .in2(_gnd_net_),
            .in3(N__47115),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48691),
            .ce(N__46115),
            .sr(N__48196));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_13_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_13_14_3 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_13_14_3  (
            .in0(N__32024),
            .in1(N__44137),
            .in2(N__36047),
            .in3(N__36214),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_13_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_13_14_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_13_14_4  (
            .in0(N__42199),
            .in1(N__38584),
            .in2(_gnd_net_),
            .in3(N__47112),
            .lcout(elapsed_time_ns_1_RNI0AOBB_0_13),
            .ltout(elapsed_time_ns_1_RNI0AOBB_0_13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_13_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_13_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_13_14_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_13_LC_13_14_5  (
            .in0(N__47113),
            .in1(_gnd_net_),
            .in2(N__32012),
            .in3(N__42200),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48691),
            .ce(N__46115),
            .sr(N__48196));
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_13_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_13_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_13_14_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_14_LC_13_14_7  (
            .in0(N__47114),
            .in1(N__46298),
            .in2(_gnd_net_),
            .in3(N__46337),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48691),
            .ce(N__46115),
            .sr(N__48196));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_13_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_13_15_0 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_13_15_0  (
            .in0(N__32009),
            .in1(N__33079),
            .in2(N__31988),
            .in3(N__33470),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_13_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_13_15_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_13_15_1  (
            .in0(N__33468),
            .in1(N__32248),
            .in2(N__33219),
            .in3(N__32194),
            .lcout(\current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_13_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_13_15_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_13_15_3  (
            .in0(N__33467),
            .in1(N__32156),
            .in2(N__33218),
            .in3(N__32117),
            .lcout(\current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_13_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_13_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_13_15_4 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_13_15_4  (
            .in0(N__32516),
            .in1(N__33075),
            .in2(N__32483),
            .in3(N__33469),
            .lcout(\current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_13_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_13_15_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_13_15_5  (
            .in0(N__33466),
            .in1(N__32422),
            .in2(N__33220),
            .in3(N__32374),
            .lcout(\current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_13_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_13_16_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_13_16_0  (
            .in0(N__33515),
            .in1(N__32339),
            .in2(N__33221),
            .in3(N__32294),
            .lcout(\current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_13_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_13_16_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_13_16_1  (
            .in0(N__33086),
            .in1(N__33517),
            .in2(N__32252),
            .in3(N__32195),
            .lcout(\current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_13_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_13_16_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_13_16_4  (
            .in0(N__33516),
            .in1(N__32155),
            .in2(N__33222),
            .in3(N__32113),
            .lcout(\current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D2_LC_13_16_6.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_13_16_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_13_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D2_LC_13_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32072),
            .lcout(il_max_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48681),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_13_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_13_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_13_17_2 .LUT_INIT=16'b1101000011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_13_17_2  (
            .in0(N__35120),
            .in1(N__42699),
            .in2(N__42340),
            .in3(N__35092),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48677),
            .ce(),
            .sr(N__48218));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_13_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_13_18_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_13_18_2  (
            .in0(N__33223),
            .in1(N__33385),
            .in2(N__33863),
            .in3(N__33815),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_13_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_13_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_13_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_13_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33779),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48672),
            .ce(N__33736),
            .sr(N__48224));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_13_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_13_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_13_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33713),
            .lcout(\current_shift_inst.un4_control_input1_1 ),
            .ltout(\current_shift_inst.un4_control_input1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_13_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_13_18_6 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_13_18_6  (
            .in0(_gnd_net_),
            .in1(N__33383),
            .in2(N__33671),
            .in3(N__33667),
            .lcout(\current_shift_inst.un38_control_input_cry_0_s0_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_13_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_13_18_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_13_18_7  (
            .in0(N__33384),
            .in1(N__33224),
            .in2(N__32678),
            .in3(N__32636),
            .lcout(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_21_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNII51H_LC_13_21_1  (
            .in0(_gnd_net_),
            .in1(N__36845),
            .in2(_gnd_net_),
            .in3(N__36866),
            .lcout(\current_shift_inst.timer_s1.N_162_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_21_4 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_21_4  (
            .in0(N__36847),
            .in1(N__36867),
            .in2(_gnd_net_),
            .in3(N__39335),
            .lcout(\current_shift_inst.timer_s1.N_163_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_13_21_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_13_21_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_13_21_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pwm_generator_inst.counter_RNISQD2_0_LC_13_21_5  (
            .in0(_gnd_net_),
            .in1(N__34332),
            .in2(_gnd_net_),
            .in3(N__34308),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_13_21_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_13_21_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_13_21_6 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_1_LC_13_21_6  (
            .in0(N__34290),
            .in1(N__34269),
            .in2(N__34250),
            .in3(N__34245),
            .lcout(\pwm_generator_inst.un1_counterlt9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_13_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_13_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_13_21_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_13_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36846),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_13_22_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_13_22_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_13_22_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIVDL3_9_LC_13_22_4  (
            .in0(N__34086),
            .in1(N__34062),
            .in2(_gnd_net_),
            .in3(N__34044),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto9_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_13_22_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_13_22_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_5_LC_13_22_5  (
            .in0(N__34024),
            .in1(N__34003),
            .in2(N__33983),
            .in3(N__33980),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_13_23_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_13_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_13_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_13_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33935),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48653),
            .ce(),
            .sr(N__48252));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_13_23_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_13_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_13_23_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_13_23_5  (
            .in0(_gnd_net_),
            .in1(N__39893),
            .in2(_gnd_net_),
            .in3(N__39873),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48653),
            .ce(),
            .sr(N__48252));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_13_23_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_13_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_13_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_13_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33902),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48653),
            .ce(),
            .sr(N__48252));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_13_24_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_13_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_13_24_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_13_24_0  (
            .in0(_gnd_net_),
            .in1(N__34442),
            .in2(N__37310),
            .in3(N__37305),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ),
            .ltout(),
            .carryin(bfn_13_24_0_),
            .carryout(\pwm_generator_inst.un19_threshold_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_13_24_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_13_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_13_24_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_13_24_1  (
            .in0(_gnd_net_),
            .in1(N__37223),
            .in2(_gnd_net_),
            .in3(N__34412),
            .lcout(\pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_0 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_13_24_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_13_24_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_13_24_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_13_24_2  (
            .in0(_gnd_net_),
            .in1(N__34430),
            .in2(_gnd_net_),
            .in3(N__34400),
            .lcout(\pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_1 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_13_24_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_13_24_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_13_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_13_24_3  (
            .in0(_gnd_net_),
            .in1(N__34460),
            .in2(_gnd_net_),
            .in3(N__34391),
            .lcout(\pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_2 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_13_24_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_13_24_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_13_24_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_13_24_4  (
            .in0(_gnd_net_),
            .in1(N__34448),
            .in2(_gnd_net_),
            .in3(N__34382),
            .lcout(\pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_3 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_13_24_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_13_24_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_13_24_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_13_24_5  (
            .in0(_gnd_net_),
            .in1(N__34466),
            .in2(_gnd_net_),
            .in3(N__34370),
            .lcout(\pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_4 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_13_24_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_13_24_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_13_24_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_13_24_6  (
            .in0(_gnd_net_),
            .in1(N__34454),
            .in2(_gnd_net_),
            .in3(N__34361),
            .lcout(\pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_5 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_13_24_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_13_24_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_13_24_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_13_24_7  (
            .in0(_gnd_net_),
            .in1(N__34763),
            .in2(_gnd_net_),
            .in3(N__34352),
            .lcout(\pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_6 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_13_25_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_13_25_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_13_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_13_25_0  (
            .in0(_gnd_net_),
            .in1(N__34436),
            .in2(_gnd_net_),
            .in3(N__34340),
            .lcout(\pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ),
            .ltout(),
            .carryin(bfn_13_25_0_),
            .carryout(\pwm_generator_inst.un19_threshold_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_13_25_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_13_25_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_13_25_1 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_13_25_1  (
            .in0(N__37481),
            .in1(N__37514),
            .in2(N__37309),
            .in3(N__34475),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_13_25_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_13_25_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_13_25_2 .LUT_INIT=16'b1011100001110100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_13_25_2  (
            .in0(N__37439),
            .in1(N__37298),
            .in2(N__37985),
            .in3(N__37184),
            .lcout(\pwm_generator_inst.un19_threshold_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_13_25_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_13_25_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_13_25_3 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_13_25_3  (
            .in0(N__37202),
            .in1(N__40778),
            .in2(N__40763),
            .in3(N__37288),
            .lcout(\pwm_generator_inst.un19_threshold_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_13_25_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_13_25_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_13_25_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_13_25_4  (
            .in0(N__37952),
            .in1(N__37154),
            .in2(N__37307),
            .in3(N__37175),
            .lcout(\pwm_generator_inst.un19_threshold_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_13_25_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_13_25_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_13_25_6 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_13_25_6  (
            .in0(N__37193),
            .in1(N__41375),
            .in2(N__37306),
            .in3(N__41393),
            .lcout(\pwm_generator_inst.un19_threshold_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_13_25_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_13_25_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_13_25_7 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_13_25_7  (
            .in0(N__44423),
            .in1(N__37319),
            .in2(N__44402),
            .in3(N__37284),
            .lcout(\pwm_generator_inst.un19_threshold_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_13_26_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_13_26_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_13_26_0 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_13_26_0  (
            .in0(N__37538),
            .in1(N__37297),
            .in2(N__37472),
            .in3(N__37133),
            .lcout(\pwm_generator_inst.un19_threshold_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_13_26_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_13_26_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_13_26_6 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_13_26_6  (
            .in0(N__37358),
            .in1(N__37211),
            .in2(N__37418),
            .in3(N__37296),
            .lcout(\pwm_generator_inst.un19_threshold_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_13_27_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_13_27_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_13_27_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_13_27_5  (
            .in0(N__37948),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37174),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_13_27_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_13_27_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_13_27_7 .LUT_INIT=16'b1010110001011100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_13_27_7  (
            .in0(N__37142),
            .in1(N__37928),
            .in2(N__37308),
            .in3(N__37454),
            .lcout(\pwm_generator_inst.un19_threshold_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_13_28_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_13_28_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_13_28_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_axb_4_LC_13_28_0  (
            .in0(_gnd_net_),
            .in1(N__34754),
            .in2(N__34733),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_axbZ0Z_4 ),
            .ltout(),
            .carryin(bfn_13_28_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_13_28_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_13_28_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_13_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_13_28_1  (
            .in0(_gnd_net_),
            .in1(N__34715),
            .in2(N__34697),
            .in3(N__34679),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_13_28_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_13_28_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_13_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_13_28_2  (
            .in0(_gnd_net_),
            .in1(N__34676),
            .in2(N__34655),
            .in3(N__34637),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_13_28_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_13_28_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_13_28_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_13_28_3  (
            .in0(_gnd_net_),
            .in1(N__34634),
            .in2(N__34616),
            .in3(N__34595),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_13_28_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_13_28_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_13_28_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_13_28_4  (
            .in0(_gnd_net_),
            .in1(N__34592),
            .in2(N__34574),
            .in3(N__34559),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_13_28_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_13_28_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_13_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_13_28_5  (
            .in0(_gnd_net_),
            .in1(N__34556),
            .in2(N__34541),
            .in3(N__34520),
            .lcout(\pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_13_28_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_13_28_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_13_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_13_28_6  (
            .in0(_gnd_net_),
            .in1(N__34517),
            .in2(N__34499),
            .in3(N__34478),
            .lcout(\pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_13_28_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_13_28_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_13_28_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_13_28_7  (
            .in0(_gnd_net_),
            .in1(N__34994),
            .in2(N__34976),
            .in3(N__34958),
            .lcout(\pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_13_29_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_13_29_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_13_29_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_13_29_0  (
            .in0(_gnd_net_),
            .in1(N__34955),
            .in2(N__34934),
            .in3(N__34916),
            .lcout(\pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(bfn_13_29_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_13_29_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_13_29_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_13_29_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_13_29_1  (
            .in0(_gnd_net_),
            .in1(N__34913),
            .in2(N__34892),
            .in3(N__34874),
            .lcout(\pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_13_29_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_13_29_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_13_29_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_13_29_2  (
            .in0(_gnd_net_),
            .in1(N__34871),
            .in2(N__35322),
            .in3(N__34853),
            .lcout(\pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_13_29_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_13_29_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_13_29_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_13_29_3  (
            .in0(_gnd_net_),
            .in1(N__35311),
            .in2(N__34850),
            .in3(N__34829),
            .lcout(\pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_13_29_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_13_29_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_13_29_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_13_29_4  (
            .in0(_gnd_net_),
            .in1(N__34826),
            .in2(N__35323),
            .in3(N__34808),
            .lcout(\pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_13_29_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_13_29_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_13_29_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_13_29_5  (
            .in0(_gnd_net_),
            .in1(N__35315),
            .in2(N__34805),
            .in3(N__34787),
            .lcout(\pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_13_29_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_13_29_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_13_29_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_13_29_6  (
            .in0(_gnd_net_),
            .in1(N__34784),
            .in2(N__35324),
            .in3(N__34766),
            .lcout(\pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_13_29_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_13_29_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_13_29_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_13_29_7  (
            .in0(_gnd_net_),
            .in1(N__35319),
            .in2(N__35273),
            .in3(N__35255),
            .lcout(\pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_13_30_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_13_30_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_13_30_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_13_30_0  (
            .in0(N__38267),
            .in1(N__35252),
            .in2(_gnd_net_),
            .in3(N__35240),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_14_4_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_14_4_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_14_4_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_14_4_0  (
            .in0(_gnd_net_),
            .in1(N__35236),
            .in2(_gnd_net_),
            .in3(N__35201),
            .lcout(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_14_5_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_14_5_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_14_5_4 .LUT_INIT=16'b1010101000100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_14_5_4  (
            .in0(N__42392),
            .in1(N__42348),
            .in2(_gnd_net_),
            .in3(N__35041),
            .lcout(\phase_controller_inst1.stoper_hc.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_14_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_14_6_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_14_6_0 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_14_6_0  (
            .in0(N__35173),
            .in1(N__35138),
            .in2(N__35578),
            .in3(N__36120),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48782),
            .ce(),
            .sr(N__48128));
    defparam \phase_controller_inst1.stoper_hc.running_LC_14_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_LC_14_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.running_LC_14_6_3 .LUT_INIT=16'b1101010111110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_LC_14_6_3  (
            .in0(N__42356),
            .in1(N__35116),
            .in2(N__35045),
            .in3(N__35074),
            .lcout(\phase_controller_inst1.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48782),
            .ce(),
            .sr(N__48128));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_14_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_14_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_14_7_0  (
            .in0(_gnd_net_),
            .in1(N__38150),
            .in2(N__35030),
            .in3(N__35568),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_14_7_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_14_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_14_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_14_7_1  (
            .in0(_gnd_net_),
            .in1(N__35021),
            .in2(N__35009),
            .in3(N__35552),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_14_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_14_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_14_7_2  (
            .in0(_gnd_net_),
            .in1(N__35000),
            .in2(N__41327),
            .in3(N__35525),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_14_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_14_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_14_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_14_7_3  (
            .in0(_gnd_net_),
            .in1(N__38351),
            .in2(N__35393),
            .in3(N__35507),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_14_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_14_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_14_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_14_7_4  (
            .in0(_gnd_net_),
            .in1(N__38345),
            .in2(N__35384),
            .in3(N__35828),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_14_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_14_7_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_14_7_5  (
            .in0(N__35807),
            .in1(N__35375),
            .in2(N__38339),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_14_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_14_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_14_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_14_7_6  (
            .in0(_gnd_net_),
            .in1(N__35369),
            .in2(N__38171),
            .in3(N__35789),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_14_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_14_7_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_14_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_14_7_7  (
            .in0(_gnd_net_),
            .in1(N__38156),
            .in2(N__35363),
            .in3(N__35771),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_14_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_14_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(N__38162),
            .in2(N__35354),
            .in3(N__35753),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_14_8_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_14_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_14_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_14_8_1  (
            .in0(_gnd_net_),
            .in1(N__38435),
            .in2(N__35345),
            .in3(N__35735),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_14_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_14_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_14_8_2  (
            .in0(_gnd_net_),
            .in1(N__38618),
            .in2(N__35333),
            .in3(N__35717),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_14_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_14_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_14_8_3  (
            .in0(_gnd_net_),
            .in1(N__38630),
            .in2(N__35492),
            .in3(N__35699),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_14_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_14_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_14_8_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_14_8_4  (
            .in0(N__35939),
            .in1(N__35483),
            .in2(N__35468),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_14_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_14_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_14_8_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_14_8_5  (
            .in0(N__35921),
            .in1(N__35459),
            .in2(N__35447),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_14_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_14_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_14_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_14_8_6  (
            .in0(_gnd_net_),
            .in1(N__35438),
            .in2(N__35426),
            .in3(N__35903),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_14_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_14_8_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_14_8_7  (
            .in0(_gnd_net_),
            .in1(N__35417),
            .in2(N__35408),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_14_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_14_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_14_9_0  (
            .in0(_gnd_net_),
            .in1(N__38069),
            .in2(N__38144),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_9_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_14_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_14_9_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_14_9_1  (
            .in0(_gnd_net_),
            .in1(N__38516),
            .in2(N__38468),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_14_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_14_9_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_14_9_2  (
            .in0(_gnd_net_),
            .in1(N__38369),
            .in2(N__38423),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_14_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_14_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_14_9_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_14_9_3  (
            .in0(_gnd_net_),
            .in1(N__38276),
            .in2(N__38330),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_14_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_14_9_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_14_9_4  (
            .in0(_gnd_net_),
            .in1(N__41960),
            .in2(N__42038),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_14_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_14_9_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_14_9_5  (
            .in0(_gnd_net_),
            .in1(N__35681),
            .in2(N__35669),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_14_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_14_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_14_9_6  (
            .in0(_gnd_net_),
            .in1(N__35654),
            .in2(N__35642),
            .in3(N__35609),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_14_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_14_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_14_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35606),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_10_0  (
            .in0(_gnd_net_),
            .in1(N__35585),
            .in2(N__35579),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_10_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_14_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_14_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_14_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_14_10_1  (
            .in0(N__36169),
            .in1(N__35551),
            .in2(_gnd_net_),
            .in3(N__35537),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__48738),
            .ce(),
            .sr(N__48153));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_14_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_14_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_14_10_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_14_10_2  (
            .in0(N__36173),
            .in1(N__35524),
            .in2(N__35534),
            .in3(N__35510),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__48738),
            .ce(),
            .sr(N__48153));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_10_3  (
            .in0(N__36170),
            .in1(N__35506),
            .in2(_gnd_net_),
            .in3(N__35831),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__48738),
            .ce(),
            .sr(N__48153));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_14_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_14_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_14_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_14_10_4  (
            .in0(N__36174),
            .in1(N__35824),
            .in2(_gnd_net_),
            .in3(N__35810),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__48738),
            .ce(),
            .sr(N__48153));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_14_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_14_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_14_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_14_10_5  (
            .in0(N__36171),
            .in1(N__35806),
            .in2(_gnd_net_),
            .in3(N__35792),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__48738),
            .ce(),
            .sr(N__48153));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_14_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_14_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_14_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_14_10_6  (
            .in0(N__36175),
            .in1(N__35788),
            .in2(_gnd_net_),
            .in3(N__35774),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__48738),
            .ce(),
            .sr(N__48153));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_10_7  (
            .in0(N__36172),
            .in1(N__35770),
            .in2(_gnd_net_),
            .in3(N__35756),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__48738),
            .ce(),
            .sr(N__48153));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_11_0  (
            .in0(N__36124),
            .in1(N__35752),
            .in2(_gnd_net_),
            .in3(N__35738),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_14_11_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__48728),
            .ce(),
            .sr(N__48161));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_14_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_14_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_14_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_14_11_1  (
            .in0(N__36183),
            .in1(N__35734),
            .in2(_gnd_net_),
            .in3(N__35720),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__48728),
            .ce(),
            .sr(N__48161));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_14_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_14_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_14_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_14_11_2  (
            .in0(N__36121),
            .in1(N__35716),
            .in2(_gnd_net_),
            .in3(N__35702),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__48728),
            .ce(),
            .sr(N__48161));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_11_3  (
            .in0(N__36184),
            .in1(N__35698),
            .in2(_gnd_net_),
            .in3(N__35684),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__48728),
            .ce(),
            .sr(N__48161));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_11_4  (
            .in0(N__36122),
            .in1(N__35938),
            .in2(_gnd_net_),
            .in3(N__35924),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__48728),
            .ce(),
            .sr(N__48161));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_11_5  (
            .in0(N__36185),
            .in1(N__35920),
            .in2(_gnd_net_),
            .in3(N__35906),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__48728),
            .ce(),
            .sr(N__48161));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_11_6  (
            .in0(N__36123),
            .in1(N__35902),
            .in2(_gnd_net_),
            .in3(N__35888),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__48728),
            .ce(),
            .sr(N__48161));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_11_7  (
            .in0(N__36186),
            .in1(N__35884),
            .in2(_gnd_net_),
            .in3(N__35867),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__48728),
            .ce(),
            .sr(N__48161));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_12_0  (
            .in0(N__36187),
            .in1(N__35864),
            .in2(_gnd_net_),
            .in3(N__35846),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_14_12_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__48719),
            .ce(),
            .sr(N__48169));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_12_1  (
            .in0(N__36191),
            .in1(N__38083),
            .in2(_gnd_net_),
            .in3(N__35843),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__48719),
            .ce(),
            .sr(N__48169));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_14_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_14_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_14_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_14_12_2  (
            .in0(N__36188),
            .in1(N__38128),
            .in2(_gnd_net_),
            .in3(N__35840),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(N__48719),
            .ce(),
            .sr(N__48169));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_14_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_14_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_14_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_14_12_3  (
            .in0(N__36192),
            .in1(N__38503),
            .in2(_gnd_net_),
            .in3(N__35837),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(N__48719),
            .ce(),
            .sr(N__48169));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_14_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_14_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_14_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_14_12_4  (
            .in0(N__36189),
            .in1(N__38485),
            .in2(_gnd_net_),
            .in3(N__35834),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ),
            .clk(N__48719),
            .ce(),
            .sr(N__48169));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_14_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_14_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_14_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_14_12_5  (
            .in0(N__36193),
            .in1(N__38389),
            .in2(_gnd_net_),
            .in3(N__36002),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ),
            .clk(N__48719),
            .ce(),
            .sr(N__48169));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_14_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_14_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_14_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_14_12_6  (
            .in0(N__36190),
            .in1(N__38408),
            .in2(_gnd_net_),
            .in3(N__35999),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ),
            .clk(N__48719),
            .ce(),
            .sr(N__48169));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_14_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_14_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_14_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_14_12_7  (
            .in0(N__36194),
            .in1(N__38290),
            .in2(_gnd_net_),
            .in3(N__35996),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ),
            .clk(N__48719),
            .ce(),
            .sr(N__48169));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_14_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_14_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_14_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_14_13_0  (
            .in0(N__36176),
            .in1(N__38314),
            .in2(_gnd_net_),
            .in3(N__35993),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_14_13_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ),
            .clk(N__48709),
            .ce(),
            .sr(N__48178));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_14_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_14_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_14_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_14_13_1  (
            .in0(N__36180),
            .in1(N__41986),
            .in2(_gnd_net_),
            .in3(N__35990),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ),
            .clk(N__48709),
            .ce(),
            .sr(N__48178));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_14_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_14_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_14_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_14_13_2  (
            .in0(N__36177),
            .in1(N__42019),
            .in2(_gnd_net_),
            .in3(N__35987),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ),
            .clk(N__48709),
            .ce(),
            .sr(N__48178));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_14_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_14_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_14_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_14_13_3  (
            .in0(N__36181),
            .in1(N__35983),
            .in2(_gnd_net_),
            .in3(N__35966),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ),
            .clk(N__48709),
            .ce(),
            .sr(N__48178));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_14_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_14_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_14_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_14_13_4  (
            .in0(N__36178),
            .in1(N__35962),
            .in2(_gnd_net_),
            .in3(N__35942),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ),
            .clk(N__48709),
            .ce(),
            .sr(N__48178));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_14_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_14_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_14_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_14_13_5  (
            .in0(N__36182),
            .in1(N__36215),
            .in2(_gnd_net_),
            .in3(N__36197),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ),
            .clk(N__48709),
            .ce(),
            .sr(N__48178));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_14_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_14_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_14_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_14_13_6  (
            .in0(N__36179),
            .in1(N__36045),
            .in2(_gnd_net_),
            .in3(N__36050),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48709),
            .ce(),
            .sr(N__48178));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_14_14_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_14_14_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_14_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_14_14_0  (
            .in0(N__36717),
            .in1(N__38562),
            .in2(_gnd_net_),
            .in3(N__36023),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__48700),
            .ce(N__43940),
            .sr(N__48188));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_14_14_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_14_14_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_14_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_14_14_1  (
            .in0(N__36709),
            .in1(N__38535),
            .in2(_gnd_net_),
            .in3(N__36020),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__48700),
            .ce(N__43940),
            .sr(N__48188));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_14_14_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_14_14_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_14_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_14_14_2  (
            .in0(N__36718),
            .in1(N__38833),
            .in2(_gnd_net_),
            .in3(N__36017),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__48700),
            .ce(N__43940),
            .sr(N__48188));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_14_14_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_14_14_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_14_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_14_14_3  (
            .in0(N__36710),
            .in1(N__38809),
            .in2(_gnd_net_),
            .in3(N__36014),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__48700),
            .ce(N__43940),
            .sr(N__48188));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_14_14_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_14_14_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_14_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_14_14_4  (
            .in0(N__36719),
            .in1(N__38785),
            .in2(_gnd_net_),
            .in3(N__36011),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__48700),
            .ce(N__43940),
            .sr(N__48188));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_14_14_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_14_14_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_14_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_14_14_5  (
            .in0(N__36711),
            .in1(N__38761),
            .in2(_gnd_net_),
            .in3(N__36008),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__48700),
            .ce(N__43940),
            .sr(N__48188));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_14_14_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_14_14_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_14_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_14_14_6  (
            .in0(N__36720),
            .in1(N__38737),
            .in2(_gnd_net_),
            .in3(N__36005),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__48700),
            .ce(N__43940),
            .sr(N__48188));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_14_14_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_14_14_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_14_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_14_14_7  (
            .in0(N__36712),
            .in1(N__38713),
            .in2(_gnd_net_),
            .in3(N__36242),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__48700),
            .ce(N__43940),
            .sr(N__48188));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_14_15_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_14_15_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_14_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_14_15_0  (
            .in0(N__36716),
            .in1(N__38689),
            .in2(_gnd_net_),
            .in3(N__36239),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__48692),
            .ce(N__43939),
            .sr(N__48197));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_14_15_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_14_15_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_14_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_14_15_1  (
            .in0(N__36724),
            .in1(N__38665),
            .in2(_gnd_net_),
            .in3(N__36236),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__48692),
            .ce(N__43939),
            .sr(N__48197));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_14_15_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_14_15_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_14_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_14_15_2  (
            .in0(N__36713),
            .in1(N__39023),
            .in2(_gnd_net_),
            .in3(N__36233),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__48692),
            .ce(N__43939),
            .sr(N__48197));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_14_15_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_14_15_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_14_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_14_15_3  (
            .in0(N__36721),
            .in1(N__39001),
            .in2(_gnd_net_),
            .in3(N__36230),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__48692),
            .ce(N__43939),
            .sr(N__48197));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_14_15_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_14_15_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_14_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_14_15_4  (
            .in0(N__36714),
            .in1(N__38979),
            .in2(_gnd_net_),
            .in3(N__36227),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__48692),
            .ce(N__43939),
            .sr(N__48197));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_14_15_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_14_15_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_14_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_14_15_5  (
            .in0(N__36722),
            .in1(N__38953),
            .in2(_gnd_net_),
            .in3(N__36224),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__48692),
            .ce(N__43939),
            .sr(N__48197));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_14_15_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_14_15_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_14_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_14_15_6  (
            .in0(N__36715),
            .in1(N__38929),
            .in2(_gnd_net_),
            .in3(N__36221),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__48692),
            .ce(N__43939),
            .sr(N__48197));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_14_15_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_14_15_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_14_15_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_14_15_7  (
            .in0(N__36723),
            .in1(N__38905),
            .in2(_gnd_net_),
            .in3(N__36218),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__48692),
            .ce(N__43939),
            .sr(N__48197));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_14_16_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_14_16_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_14_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_14_16_0  (
            .in0(N__36703),
            .in1(N__38881),
            .in2(_gnd_net_),
            .in3(N__36269),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__48686),
            .ce(N__43938),
            .sr(N__48205));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_14_16_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_14_16_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_14_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_14_16_1  (
            .in0(N__36725),
            .in1(N__38857),
            .in2(_gnd_net_),
            .in3(N__36266),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__48686),
            .ce(N__43938),
            .sr(N__48205));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_14_16_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_14_16_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_14_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_14_16_2  (
            .in0(N__36704),
            .in1(N__39244),
            .in2(_gnd_net_),
            .in3(N__36263),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__48686),
            .ce(N__43938),
            .sr(N__48205));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_14_16_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_14_16_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_14_16_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_14_16_3  (
            .in0(N__36726),
            .in1(N__39220),
            .in2(_gnd_net_),
            .in3(N__36260),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__48686),
            .ce(N__43938),
            .sr(N__48205));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_14_16_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_14_16_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_14_16_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_14_16_4  (
            .in0(N__36705),
            .in1(N__39196),
            .in2(_gnd_net_),
            .in3(N__36257),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__48686),
            .ce(N__43938),
            .sr(N__48205));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_14_16_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_14_16_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_14_16_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_14_16_5  (
            .in0(N__36727),
            .in1(N__39172),
            .in2(_gnd_net_),
            .in3(N__36254),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__48686),
            .ce(N__43938),
            .sr(N__48205));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_14_16_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_14_16_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_14_16_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_14_16_6  (
            .in0(N__36706),
            .in1(N__39148),
            .in2(_gnd_net_),
            .in3(N__36251),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__48686),
            .ce(N__43938),
            .sr(N__48205));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_14_16_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_14_16_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_14_16_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_14_16_7  (
            .in0(N__36728),
            .in1(N__39124),
            .in2(_gnd_net_),
            .in3(N__36248),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__48686),
            .ce(N__43938),
            .sr(N__48205));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_14_17_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_14_17_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_14_17_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_14_17_0  (
            .in0(N__36699),
            .in1(N__39100),
            .in2(_gnd_net_),
            .in3(N__36245),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__48682),
            .ce(N__43934),
            .sr(N__48212));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_14_17_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_14_17_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_14_17_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_14_17_1  (
            .in0(N__36707),
            .in1(N__39076),
            .in2(_gnd_net_),
            .in3(N__36743),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__48682),
            .ce(N__43934),
            .sr(N__48212));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_14_17_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_14_17_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_14_17_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_14_17_2  (
            .in0(N__36700),
            .in1(N__39056),
            .in2(_gnd_net_),
            .in3(N__36740),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__48682),
            .ce(N__43934),
            .sr(N__48212));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_14_17_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_14_17_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_14_17_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_14_17_3  (
            .in0(N__36708),
            .in1(N__39418),
            .in2(_gnd_net_),
            .in3(N__36737),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__48682),
            .ce(N__43934),
            .sr(N__48212));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_14_17_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_14_17_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_14_17_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_14_17_4  (
            .in0(N__36701),
            .in1(N__39040),
            .in2(_gnd_net_),
            .in3(N__36734),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__48682),
            .ce(N__43934),
            .sr(N__48212));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_14_17_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_14_17_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_14_17_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_14_17_5  (
            .in0(N__39434),
            .in1(N__36702),
            .in2(_gnd_net_),
            .in3(N__36731),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48682),
            .ce(N__43934),
            .sr(N__48212));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_14_17_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_14_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_14_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43985),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_14_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_14_18_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(N__42344),
            .in2(_gnd_net_),
            .in3(N__42380),
            .lcout(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_14_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_14_18_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_0_LC_14_18_7  (
            .in0(_gnd_net_),
            .in1(N__39294),
            .in2(_gnd_net_),
            .in3(N__36954),
            .lcout(\phase_controller_inst1.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_14_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_14_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_14_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_3_LC_14_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36323),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48673),
            .ce(),
            .sr(N__48225));
    defparam \phase_controller_inst1.state_3_LC_14_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_14_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_14_19_4 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \phase_controller_inst1.state_3_LC_14_19_4  (
            .in0(N__39307),
            .in1(N__44564),
            .in2(N__36959),
            .in3(N__36293),
            .lcout(state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48673),
            .ce(),
            .sr(N__48225));
    defparam \phase_controller_inst1.state_2_LC_14_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_14_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_14_19_7 .LUT_INIT=16'b1010111000001100;
    LogicCell40 \phase_controller_inst1.state_2_LC_14_19_7  (
            .in0(N__36958),
            .in1(N__44631),
            .in2(N__42710),
            .in3(N__39306),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48673),
            .ce(),
            .sr(N__48225));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_14_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_14_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_14_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_14_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36935),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48666),
            .ce(),
            .sr(N__48229));
    defparam \current_shift_inst.stop_timer_s1_LC_14_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_LC_14_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.stop_timer_s1_LC_14_21_0 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \current_shift_inst.stop_timer_s1_LC_14_21_0  (
            .in0(N__39311),
            .in1(N__39333),
            .in2(N__36872),
            .in3(N__39352),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48662),
            .ce(),
            .sr(N__48234));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_14_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_14_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_14_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_14_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36905),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48662),
            .ce(),
            .sr(N__48234));
    defparam \current_shift_inst.timer_s1.running_LC_14_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_14_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_14_21_3 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_14_21_3  (
            .in0(N__39334),
            .in1(N__36868),
            .in2(_gnd_net_),
            .in3(N__36848),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48662),
            .ce(),
            .sr(N__48234));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_14_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_14_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_14_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_14_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36829),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48659),
            .ce(),
            .sr(N__48239));
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_14_25_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_14_25_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_14_25_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_14_25_0  (
            .in0(_gnd_net_),
            .in1(N__36785),
            .in2(_gnd_net_),
            .in3(N__36803),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_0 ),
            .ltout(),
            .carryin(bfn_14_25_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_14_25_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_14_25_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_14_25_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_14_25_1  (
            .in0(_gnd_net_),
            .in1(N__36761),
            .in2(_gnd_net_),
            .in3(N__36779),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_0 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_14_25_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_14_25_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_14_25_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_14_25_2  (
            .in0(_gnd_net_),
            .in1(N__37127),
            .in2(_gnd_net_),
            .in3(N__36755),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_1 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_14_25_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_14_25_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_14_25_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_14_25_3  (
            .in0(_gnd_net_),
            .in1(N__37103),
            .in2(_gnd_net_),
            .in3(N__37121),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_2 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_14_25_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_14_25_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_14_25_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_14_25_4  (
            .in0(_gnd_net_),
            .in1(N__37079),
            .in2(_gnd_net_),
            .in3(N__37097),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_3 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_14_25_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_14_25_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_14_25_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_14_25_5  (
            .in0(_gnd_net_),
            .in1(N__37055),
            .in2(_gnd_net_),
            .in3(N__37073),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_4 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_14_25_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_14_25_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_14_25_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_14_25_6  (
            .in0(_gnd_net_),
            .in1(N__37031),
            .in2(_gnd_net_),
            .in3(N__37049),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_5 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_14_25_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_14_25_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_14_25_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_14_25_7  (
            .in0(_gnd_net_),
            .in1(N__37013),
            .in2(_gnd_net_),
            .in3(N__37025),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_6 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_14_26_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_14_26_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_14_26_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_14_26_0  (
            .in0(_gnd_net_),
            .in1(N__36989),
            .in2(_gnd_net_),
            .in3(N__37007),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_8 ),
            .ltout(),
            .carryin(bfn_14_26_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_14_26_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_14_26_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_14_26_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_14_26_1  (
            .in0(_gnd_net_),
            .in1(N__36965),
            .in2(_gnd_net_),
            .in3(N__36983),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_8 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_14_26_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_14_26_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_14_26_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_14_26_2  (
            .in0(_gnd_net_),
            .in1(N__44395),
            .in2(_gnd_net_),
            .in3(N__37313),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_9 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_14_26_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_14_26_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_14_26_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_14_26_3  (
            .in0(N__37295),
            .in1(N__37397),
            .in2(_gnd_net_),
            .in3(N__37214),
            .lcout(\pwm_generator_inst.un19_threshold_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_10 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_14_26_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_14_26_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_14_26_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_14_26_4  (
            .in0(_gnd_net_),
            .in1(N__37413),
            .in2(_gnd_net_),
            .in3(N__37205),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_11 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_14_26_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_14_26_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_14_26_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_14_26_5  (
            .in0(_gnd_net_),
            .in1(N__40749),
            .in2(_gnd_net_),
            .in3(N__37196),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_12 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_14_26_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_14_26_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_14_26_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_14_26_6  (
            .in0(_gnd_net_),
            .in1(N__41367),
            .in2(_gnd_net_),
            .in3(N__37187),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_13 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_14_26_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_14_26_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_14_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_14_26_7  (
            .in0(_gnd_net_),
            .in1(N__37434),
            .in2(_gnd_net_),
            .in3(N__37178),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_14 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_14_27_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_14_27_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_14_27_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_14_27_0  (
            .in0(_gnd_net_),
            .in1(N__37170),
            .in2(_gnd_net_),
            .in3(N__37145),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_14_27_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_14_27_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_14_27_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_14_27_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_14_27_1  (
            .in0(_gnd_net_),
            .in1(N__37452),
            .in2(_gnd_net_),
            .in3(N__37136),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_16 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_14_27_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_14_27_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_14_27_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_14_27_2  (
            .in0(_gnd_net_),
            .in1(N__37467),
            .in2(_gnd_net_),
            .in3(N__37487),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_17 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_14_27_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_14_27_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_14_27_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_14_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37484),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_14_27_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_14_27_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_14_27_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_14_27_4  (
            .in0(_gnd_net_),
            .in1(N__37534),
            .in2(_gnd_net_),
            .in3(N__37468),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_14_27_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_14_27_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_14_27_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_14_27_5  (
            .in0(_gnd_net_),
            .in1(N__37927),
            .in2(_gnd_net_),
            .in3(N__37453),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_14_27_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_14_27_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_14_27_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_14_27_6  (
            .in0(_gnd_net_),
            .in1(N__37978),
            .in2(_gnd_net_),
            .in3(N__37438),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_14_27_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_14_27_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_14_27_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_14_27_7  (
            .in0(_gnd_net_),
            .in1(N__37354),
            .in2(_gnd_net_),
            .in3(N__37417),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_14_28_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_14_28_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_14_28_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_LC_14_28_0  (
            .in0(_gnd_net_),
            .in1(N__37393),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_28_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_14_28_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_14_28_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_14_28_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_14_28_1  (
            .in0(_gnd_net_),
            .in1(N__37370),
            .in2(_gnd_net_),
            .in3(N__37343),
            .lcout(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_14_28_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_14_28_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_14_28_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_14_28_2  (
            .in0(_gnd_net_),
            .in1(N__37340),
            .in2(_gnd_net_),
            .in3(N__37322),
            .lcout(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_14_28_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_14_28_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_14_28_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_14_28_3  (
            .in0(_gnd_net_),
            .in1(N__38009),
            .in2(_gnd_net_),
            .in3(N__37994),
            .lcout(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_14_28_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_14_28_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_14_28_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_14_28_4  (
            .in0(_gnd_net_),
            .in1(N__37991),
            .in2(_gnd_net_),
            .in3(N__37967),
            .lcout(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_14_28_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_14_28_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_14_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_14_28_5  (
            .in0(_gnd_net_),
            .in1(N__37632),
            .in2(N__37964),
            .in3(N__37937),
            .lcout(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_14_28_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_14_28_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_14_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_14_28_6  (
            .in0(_gnd_net_),
            .in1(N__37934),
            .in2(N__37716),
            .in3(N__37916),
            .lcout(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_14_28_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_14_28_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_14_28_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_14_28_7  (
            .in0(_gnd_net_),
            .in1(N__37636),
            .in2(N__37547),
            .in3(N__37523),
            .lcout(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_14_29_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_14_29_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_14_29_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_14_29_0  (
            .in0(_gnd_net_),
            .in1(N__37520),
            .in2(_gnd_net_),
            .in3(N__37502),
            .lcout(\pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ),
            .ltout(),
            .carryin(bfn_14_29_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_14_29_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_14_29_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_14_29_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_9_c_LC_14_29_1  (
            .in0(_gnd_net_),
            .in1(N__37499),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_14_29_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_14_29_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_14_29_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_10_c_LC_14_29_2  (
            .in0(_gnd_net_),
            .in1(N__37493),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_14_29_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_14_29_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_14_29_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_11_c_LC_14_29_3  (
            .in0(_gnd_net_),
            .in1(N__38063),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_14_29_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_14_29_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_14_29_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_12_c_LC_14_29_4  (
            .in0(_gnd_net_),
            .in1(N__38057),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_14_29_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_14_29_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_14_29_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_13_c_LC_14_29_5  (
            .in0(_gnd_net_),
            .in1(N__38051),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_14_29_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_14_29_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_14_29_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_14_c_LC_14_29_6  (
            .in0(_gnd_net_),
            .in1(N__38045),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_14_29_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_14_29_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_14_29_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_15_c_LC_14_29_7  (
            .in0(_gnd_net_),
            .in1(N__38039),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_14_30_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_14_30_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_14_30_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_16_c_LC_14_30_0  (
            .in0(_gnd_net_),
            .in1(N__38033),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_30_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_14_30_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_14_30_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_14_30_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_17_c_LC_14_30_1  (
            .in0(_gnd_net_),
            .in1(N__38027),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_14_30_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_14_30_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_14_30_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_18_c_LC_14_30_2  (
            .in0(_gnd_net_),
            .in1(N__38021),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_14_30_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_14_30_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_14_30_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_c_LC_14_30_3  (
            .in0(_gnd_net_),
            .in1(N__38015),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_14_30_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_14_30_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_14_30_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_14_30_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38270),
            .lcout(\pwm_generator_inst.un3_threshold_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_15_6_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_15_6_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_15_6_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_15_6_0  (
            .in0(N__38196),
            .in1(N__38261),
            .in2(_gnd_net_),
            .in3(N__41880),
            .lcout(elapsed_time_ns_1_RNI25DN9_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_15_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_15_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_15_7_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_7_LC_15_7_0  (
            .in0(N__47062),
            .in1(N__44882),
            .in2(_gnd_net_),
            .in3(N__44853),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48783),
            .ce(N__46107),
            .sr(N__48129));
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_15_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_15_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_15_7_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_9_LC_15_7_1  (
            .in0(N__44372),
            .in1(N__44350),
            .in2(_gnd_net_),
            .in3(N__47064),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48783),
            .ce(N__46107),
            .sr(N__48129));
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_15_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_15_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_15_7_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_8_LC_15_7_2  (
            .in0(N__47063),
            .in1(N__44937),
            .in2(_gnd_net_),
            .in3(N__44920),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48783),
            .ce(N__46107),
            .sr(N__48129));
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_15_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_15_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_15_7_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_1_LC_15_7_4  (
            .in0(N__47061),
            .in1(N__43173),
            .in2(_gnd_net_),
            .in3(N__43157),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48783),
            .ce(N__46107),
            .sr(N__48129));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_15_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_15_8_0 .LUT_INIT=16'b0101110100000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_15_8_0  (
            .in0(N__38135),
            .in1(N__41351),
            .in2(N__38093),
            .in3(N__38113),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_15_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_15_8_1 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_15_8_1  (
            .in0(N__41350),
            .in1(N__38134),
            .in2(N__38114),
            .in3(N__38092),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_15_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_15_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_15_8_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_4_LC_15_8_4  (
            .in0(N__47058),
            .in1(N__43498),
            .in2(_gnd_net_),
            .in3(N__43473),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48771),
            .ce(N__46108),
            .sr(N__48133));
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_15_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_15_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_15_8_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_5_LC_15_8_5  (
            .in0(N__45004),
            .in1(N__44964),
            .in2(_gnd_net_),
            .in3(N__47060),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48771),
            .ce(N__46108),
            .sr(N__48133));
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_15_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_15_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_15_8_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_6_LC_15_8_6  (
            .in0(N__47059),
            .in1(N__44302),
            .in2(_gnd_net_),
            .in3(N__44253),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48771),
            .ce(N__46108),
            .sr(N__48133));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_15_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_15_9_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_15_9_0  (
            .in0(N__38321),
            .in1(N__38296),
            .in2(N__41342),
            .in3(N__38606),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_15_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_15_9_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_15_9_1  (
            .in0(N__38605),
            .in1(N__38320),
            .in2(N__38300),
            .in3(N__41338),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_15_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_15_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_15_9_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_27_LC_15_9_6  (
            .in0(N__46935),
            .in1(N__43868),
            .in2(_gnd_net_),
            .in3(N__43824),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48763),
            .ce(N__46111),
            .sr(N__48139));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_15_10_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_15_10_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_15_10_0  (
            .in0(N__43472),
            .in1(N__43580),
            .in2(N__43559),
            .in3(N__43145),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_15_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_15_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_15_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_15_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38573),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48750),
            .ce(N__44117),
            .sr(N__48144));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_15_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_15_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_15_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_15_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38546),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48750),
            .ce(N__44117),
            .sr(N__48144));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_15_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_15_10_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_15_10_5  (
            .in0(N__43581),
            .in1(N__43618),
            .in2(_gnd_net_),
            .in3(N__46841),
            .lcout(elapsed_time_ns_1_RNIED91B_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_15_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_15_11_0 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_15_11_0  (
            .in0(N__38444),
            .in1(N__38453),
            .in2(N__38504),
            .in3(N__38484),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_15_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_15_11_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_15_11_1  (
            .in0(N__38452),
            .in1(N__38502),
            .in2(N__38486),
            .in3(N__38443),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_15_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_15_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_15_11_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_20_LC_15_11_2  (
            .in0(N__46932),
            .in1(N__43274),
            .in2(_gnd_net_),
            .in3(N__43245),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48739),
            .ce(N__46114),
            .sr(N__48154));
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_15_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_15_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_15_11_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_21_LC_15_11_3  (
            .in0(N__42552),
            .in1(N__42487),
            .in2(_gnd_net_),
            .in3(N__46934),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48739),
            .ce(N__46114),
            .sr(N__48154));
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_15_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_15_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_15_11_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_10_LC_15_11_7  (
            .in0(N__42104),
            .in1(N__42116),
            .in2(_gnd_net_),
            .in3(N__46933),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48739),
            .ce(N__46114),
            .sr(N__48154));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_15_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_15_12_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_15_12_0  (
            .in0(N__38385),
            .in1(N__38406),
            .in2(N__38645),
            .in3(N__38360),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_15_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_15_12_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_15_12_1  (
            .in0(N__38359),
            .in1(N__38407),
            .in2(N__38390),
            .in3(N__38641),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_15_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_15_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_15_12_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_22_LC_15_12_2  (
            .in0(N__47231),
            .in1(N__47209),
            .in2(_gnd_net_),
            .in3(N__47144),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48729),
            .ce(N__46116),
            .sr(N__48162));
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_15_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_15_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_15_12_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_23_LC_15_12_3  (
            .in0(N__47348),
            .in1(N__47319),
            .in2(_gnd_net_),
            .in3(N__47110),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48729),
            .ce(N__46116),
            .sr(N__48162));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_15_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_15_12_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_15_12_4  (
            .in0(N__42071),
            .in1(N__42049),
            .in2(_gnd_net_),
            .in3(N__47141),
            .lcout(elapsed_time_ns_1_RNIV8OBB_0_12),
            .ltout(elapsed_time_ns_1_RNIV8OBB_0_12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_15_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_15_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_15_12_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_12_LC_15_12_5  (
            .in0(_gnd_net_),
            .in1(N__47111),
            .in2(N__38633),
            .in3(N__42072),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48729),
            .ce(N__46116),
            .sr(N__48162));
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_15_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_15_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_15_12_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_11_LC_15_12_6  (
            .in0(N__45996),
            .in1(N__45974),
            .in2(_gnd_net_),
            .in3(N__47143),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48729),
            .ce(N__46116),
            .sr(N__48162));
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_15_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_15_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_15_12_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_24_LC_15_12_7  (
            .in0(N__47142),
            .in1(N__45540),
            .in2(_gnd_net_),
            .in3(N__45522),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48729),
            .ce(N__46116),
            .sr(N__48162));
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_15_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_15_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_15_13_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_13_LC_15_13_0  (
            .in0(N__42193),
            .in1(N__38591),
            .in2(_gnd_net_),
            .in3(N__47109),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48720),
            .ce(N__46677),
            .sr(N__48170));
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_15_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_15_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_15_13_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_16_LC_15_13_1  (
            .in0(N__47107),
            .in1(N__42169),
            .in2(_gnd_net_),
            .in3(N__42258),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48720),
            .ce(N__46677),
            .sr(N__48170));
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_15_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_15_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_15_13_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_17_LC_15_13_3  (
            .in0(N__47108),
            .in1(N__42216),
            .in2(_gnd_net_),
            .in3(N__42523),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48720),
            .ce(N__46677),
            .sr(N__48170));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_15_14_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_15_14_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_15_14_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(N__38832),
            .in2(N__38569),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_15_14_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__48710),
            .ce(N__44112),
            .sr(N__48179));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_15_14_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_15_14_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_15_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(N__38808),
            .in2(N__38542),
            .in3(N__38519),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__48710),
            .ce(N__44112),
            .sr(N__48179));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_15_14_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_15_14_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_15_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_15_14_2  (
            .in0(_gnd_net_),
            .in1(N__38784),
            .in2(N__38837),
            .in3(N__38816),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__48710),
            .ce(N__44112),
            .sr(N__48179));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_15_14_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_15_14_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_15_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(N__38760),
            .in2(N__38813),
            .in3(N__38792),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__48710),
            .ce(N__44112),
            .sr(N__48179));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_15_14_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_15_14_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_15_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_15_14_4  (
            .in0(_gnd_net_),
            .in1(N__38736),
            .in2(N__38789),
            .in3(N__38768),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__48710),
            .ce(N__44112),
            .sr(N__48179));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_15_14_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_15_14_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_15_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_15_14_5  (
            .in0(_gnd_net_),
            .in1(N__38712),
            .in2(N__38765),
            .in3(N__38744),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__48710),
            .ce(N__44112),
            .sr(N__48179));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_15_14_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_15_14_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_15_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(N__38688),
            .in2(N__38741),
            .in3(N__38720),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__48710),
            .ce(N__44112),
            .sr(N__48179));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_15_14_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_15_14_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_15_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_15_14_7  (
            .in0(_gnd_net_),
            .in1(N__38664),
            .in2(N__38717),
            .in3(N__38696),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__48710),
            .ce(N__44112),
            .sr(N__48179));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_15_15_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_15_15_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_15_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_15_15_0  (
            .in0(_gnd_net_),
            .in1(N__39021),
            .in2(N__38693),
            .in3(N__38672),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_15_15_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__48701),
            .ce(N__44116),
            .sr(N__48189));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_15_15_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_15_15_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_15_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_15_15_1  (
            .in0(_gnd_net_),
            .in1(N__39000),
            .in2(N__38669),
            .in3(N__38648),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__48701),
            .ce(N__44116),
            .sr(N__48189));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_15_15_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_15_15_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_15_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_15_15_2  (
            .in0(_gnd_net_),
            .in1(N__39022),
            .in2(N__38980),
            .in3(N__39008),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__48701),
            .ce(N__44116),
            .sr(N__48189));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_15_15_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_15_15_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_15_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_15_15_3  (
            .in0(_gnd_net_),
            .in1(N__38952),
            .in2(N__39005),
            .in3(N__38984),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__48701),
            .ce(N__44116),
            .sr(N__48189));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_15_15_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_15_15_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_15_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_15_15_4  (
            .in0(_gnd_net_),
            .in1(N__38928),
            .in2(N__38981),
            .in3(N__38960),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__48701),
            .ce(N__44116),
            .sr(N__48189));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_15_15_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_15_15_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_15_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_15_15_5  (
            .in0(_gnd_net_),
            .in1(N__38904),
            .in2(N__38957),
            .in3(N__38936),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__48701),
            .ce(N__44116),
            .sr(N__48189));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_15_15_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_15_15_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_15_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_15_15_6  (
            .in0(_gnd_net_),
            .in1(N__38880),
            .in2(N__38933),
            .in3(N__38912),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__48701),
            .ce(N__44116),
            .sr(N__48189));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_15_15_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_15_15_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_15_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_15_15_7  (
            .in0(_gnd_net_),
            .in1(N__38856),
            .in2(N__38909),
            .in3(N__38888),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__48701),
            .ce(N__44116),
            .sr(N__48189));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_15_16_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_15_16_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_15_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_15_16_0  (
            .in0(_gnd_net_),
            .in1(N__39243),
            .in2(N__38885),
            .in3(N__38864),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_15_16_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__48693),
            .ce(N__44108),
            .sr(N__48198));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_15_16_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_15_16_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_15_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_15_16_1  (
            .in0(_gnd_net_),
            .in1(N__39219),
            .in2(N__38861),
            .in3(N__38840),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__48693),
            .ce(N__44108),
            .sr(N__48198));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_15_16_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_15_16_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_15_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_15_16_2  (
            .in0(_gnd_net_),
            .in1(N__39195),
            .in2(N__39248),
            .in3(N__39227),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__48693),
            .ce(N__44108),
            .sr(N__48198));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_15_16_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_15_16_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_15_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_15_16_3  (
            .in0(_gnd_net_),
            .in1(N__39171),
            .in2(N__39224),
            .in3(N__39203),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__48693),
            .ce(N__44108),
            .sr(N__48198));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_15_16_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_15_16_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_15_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_15_16_4  (
            .in0(_gnd_net_),
            .in1(N__39147),
            .in2(N__39200),
            .in3(N__39179),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__48693),
            .ce(N__44108),
            .sr(N__48198));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_15_16_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_15_16_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_15_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_15_16_5  (
            .in0(_gnd_net_),
            .in1(N__39123),
            .in2(N__39176),
            .in3(N__39155),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__48693),
            .ce(N__44108),
            .sr(N__48198));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_15_16_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_15_16_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_15_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_15_16_6  (
            .in0(_gnd_net_),
            .in1(N__39099),
            .in2(N__39152),
            .in3(N__39131),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__48693),
            .ce(N__44108),
            .sr(N__48198));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_15_16_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_15_16_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_15_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_15_16_7  (
            .in0(_gnd_net_),
            .in1(N__39075),
            .in2(N__39128),
            .in3(N__39107),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__48693),
            .ce(N__44108),
            .sr(N__48198));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_15_17_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_15_17_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_15_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_15_17_0  (
            .in0(_gnd_net_),
            .in1(N__39054),
            .in2(N__39104),
            .in3(N__39083),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_15_17_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__48687),
            .ce(N__44095),
            .sr(N__48206));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_15_17_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_15_17_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_15_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(N__39417),
            .in2(N__39080),
            .in3(N__39059),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__48687),
            .ce(N__44095),
            .sr(N__48206));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_15_17_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_15_17_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_15_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_15_17_2  (
            .in0(_gnd_net_),
            .in1(N__39055),
            .in2(N__39041),
            .in3(N__39026),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__48687),
            .ce(N__44095),
            .sr(N__48206));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_15_17_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_15_17_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_15_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(N__39433),
            .in2(N__39422),
            .in3(N__39401),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__48687),
            .ce(N__44095),
            .sr(N__48206));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_15_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_15_17_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_15_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39398),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48687),
            .ce(N__44095),
            .sr(N__48206));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_15_18_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_15_18_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_15_18_2 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_15_18_2  (
            .in0(N__43999),
            .in1(N__43964),
            .in2(_gnd_net_),
            .in3(N__44018),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48683),
            .ce(),
            .sr(N__48213));
    defparam \phase_controller_inst1.start_timer_hc_LC_15_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_15_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_15_18_6 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_15_18_6  (
            .in0(N__42967),
            .in1(N__42668),
            .in2(N__42388),
            .in3(N__39395),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48683),
            .ce(),
            .sr(N__48213));
    defparam \delay_measurement_inst.start_timer_tr_LC_15_19_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_15_19_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_tr_LC_15_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_15_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43965),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42721),
            .ce(),
            .sr(N__48219));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_15_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_15_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_15_20_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_15_20_2  (
            .in0(_gnd_net_),
            .in1(N__39388),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48674),
            .ce(),
            .sr(N__48226));
    defparam \phase_controller_inst1.S1_LC_15_21_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_15_21_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_15_21_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.S1_LC_15_21_1  (
            .in0(N__39309),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48667),
            .ce(),
            .sr(N__48230));
    defparam \current_shift_inst.start_timer_s1_LC_15_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_15_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.start_timer_s1_LC_15_21_2 .LUT_INIT=16'b1011101101000100;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_15_21_2  (
            .in0(N__39351),
            .in1(N__39308),
            .in2(_gnd_net_),
            .in3(N__39332),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48667),
            .ce(),
            .sr(N__48230));
    defparam \phase_controller_inst1.T01_LC_15_22_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.T01_LC_15_22_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T01_LC_15_22_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \phase_controller_inst1.T01_LC_15_22_5  (
            .in0(_gnd_net_),
            .in1(N__39259),
            .in2(_gnd_net_),
            .in3(N__39310),
            .lcout(T01_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48663),
            .ce(),
            .sr(N__48235));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_15_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_15_23_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_15_23_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_15_23_0  (
            .in0(_gnd_net_),
            .in1(N__39892),
            .in2(N__39878),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_23_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_15_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_15_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_15_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_15_23_1  (
            .in0(_gnd_net_),
            .in1(N__39809),
            .in2(N__39800),
            .in3(N__39773),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .clk(N__48660),
            .ce(),
            .sr(N__48240));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_15_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_15_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_15_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_15_23_2  (
            .in0(_gnd_net_),
            .in1(N__39770),
            .in2(N__39758),
            .in3(N__39710),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .clk(N__48660),
            .ce(),
            .sr(N__48240));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_15_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_15_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_15_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_15_23_3  (
            .in0(_gnd_net_),
            .in1(N__39707),
            .in2(N__39695),
            .in3(N__39650),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__48660),
            .ce(),
            .sr(N__48240));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_15_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_15_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_15_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_15_23_4  (
            .in0(_gnd_net_),
            .in1(N__39646),
            .in2(N__39605),
            .in3(N__39593),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__48660),
            .ce(),
            .sr(N__48240));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_15_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_15_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_15_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_15_23_5  (
            .in0(_gnd_net_),
            .in1(N__39590),
            .in2(N__39580),
            .in3(N__39542),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__48660),
            .ce(),
            .sr(N__48240));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_15_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_15_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_15_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_15_23_6  (
            .in0(_gnd_net_),
            .in1(N__39539),
            .in2(N__39530),
            .in3(N__39488),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__48660),
            .ce(),
            .sr(N__48240));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_15_23_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_15_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_15_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_15_23_7  (
            .in0(_gnd_net_),
            .in1(N__39485),
            .in2(N__39476),
            .in3(N__39437),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__48660),
            .ce(),
            .sr(N__48240));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_15_24_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_15_24_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_15_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_15_24_0  (
            .in0(_gnd_net_),
            .in1(N__40343),
            .in2(N__40334),
            .in3(N__40283),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(bfn_15_24_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__48657),
            .ce(),
            .sr(N__48245));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_15_24_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_15_24_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_15_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_15_24_1  (
            .in0(_gnd_net_),
            .in1(N__40280),
            .in2(N__40271),
            .in3(N__40217),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__48657),
            .ce(),
            .sr(N__48245));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_15_24_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_15_24_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_15_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_15_24_2  (
            .in0(_gnd_net_),
            .in1(N__40214),
            .in2(N__40202),
            .in3(N__40151),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__48657),
            .ce(),
            .sr(N__48245));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_15_24_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_15_24_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_15_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_15_24_3  (
            .in0(_gnd_net_),
            .in1(N__40148),
            .in2(N__40136),
            .in3(N__40085),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__48657),
            .ce(),
            .sr(N__48245));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_15_24_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_15_24_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_15_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_15_24_4  (
            .in0(_gnd_net_),
            .in1(N__40082),
            .in2(N__40043),
            .in3(N__40031),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__48657),
            .ce(),
            .sr(N__48245));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_15_24_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_15_24_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_15_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_15_24_5  (
            .in0(_gnd_net_),
            .in1(N__40833),
            .in2(N__40028),
            .in3(N__39986),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__48657),
            .ce(),
            .sr(N__48245));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_15_24_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_15_24_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_15_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_15_24_6  (
            .in0(_gnd_net_),
            .in1(N__39983),
            .in2(N__40867),
            .in3(N__39941),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__48657),
            .ce(),
            .sr(N__48245));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_15_24_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_15_24_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_15_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_15_24_7  (
            .in0(_gnd_net_),
            .in1(N__40837),
            .in2(N__39938),
            .in3(N__39896),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__48657),
            .ce(),
            .sr(N__48245));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_15_25_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_15_25_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_15_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_15_25_0  (
            .in0(_gnd_net_),
            .in1(N__40838),
            .in2(N__40736),
            .in3(N__40676),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(bfn_15_25_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__48654),
            .ce(),
            .sr(N__48253));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_15_25_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_15_25_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_15_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_15_25_1  (
            .in0(_gnd_net_),
            .in1(N__40673),
            .in2(N__40868),
            .in3(N__40628),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__48654),
            .ce(),
            .sr(N__48253));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_15_25_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_15_25_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_15_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_15_25_2  (
            .in0(_gnd_net_),
            .in1(N__40842),
            .in2(N__40625),
            .in3(N__40580),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__48654),
            .ce(),
            .sr(N__48253));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_15_25_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_15_25_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_15_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_15_25_3  (
            .in0(_gnd_net_),
            .in1(N__40577),
            .in2(N__40869),
            .in3(N__40532),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__48654),
            .ce(),
            .sr(N__48253));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_15_25_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_15_25_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_15_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_15_25_4  (
            .in0(_gnd_net_),
            .in1(N__40846),
            .in2(N__40528),
            .in3(N__40487),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__48654),
            .ce(),
            .sr(N__48253));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_15_25_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_15_25_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_15_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_15_25_5  (
            .in0(_gnd_net_),
            .in1(N__40484),
            .in2(N__40870),
            .in3(N__40439),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__48654),
            .ce(),
            .sr(N__48253));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_15_25_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_15_25_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_15_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_15_25_6  (
            .in0(_gnd_net_),
            .in1(N__40850),
            .in2(N__40436),
            .in3(N__40391),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__48654),
            .ce(),
            .sr(N__48253));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_15_25_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_15_25_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_15_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_15_25_7  (
            .in0(_gnd_net_),
            .in1(N__40388),
            .in2(N__40871),
            .in3(N__40346),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__48654),
            .ce(),
            .sr(N__48253));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_15_26_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_15_26_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_15_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_15_26_0  (
            .in0(_gnd_net_),
            .in1(N__40854),
            .in2(N__41315),
            .in3(N__41273),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(bfn_15_26_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__48651),
            .ce(),
            .sr(N__48260));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_15_26_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_15_26_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_15_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_15_26_1  (
            .in0(_gnd_net_),
            .in1(N__41269),
            .in2(N__40872),
            .in3(N__41234),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__48651),
            .ce(),
            .sr(N__48260));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_15_26_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_15_26_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_15_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_15_26_2  (
            .in0(_gnd_net_),
            .in1(N__40858),
            .in2(N__41231),
            .in3(N__41183),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__48651),
            .ce(),
            .sr(N__48260));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_15_26_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_15_26_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_15_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_15_26_3  (
            .in0(_gnd_net_),
            .in1(N__41180),
            .in2(N__40873),
            .in3(N__41144),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__48651),
            .ce(),
            .sr(N__48260));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_15_26_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_15_26_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_15_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_15_26_4  (
            .in0(_gnd_net_),
            .in1(N__40862),
            .in2(N__41141),
            .in3(N__41099),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__48651),
            .ce(),
            .sr(N__48260));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_15_26_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_15_26_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_15_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_15_26_5  (
            .in0(_gnd_net_),
            .in1(N__41096),
            .in2(N__40874),
            .in3(N__41054),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__48651),
            .ce(),
            .sr(N__48260));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_15_26_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_15_26_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_15_26_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_15_26_6  (
            .in0(N__41051),
            .in1(N__40866),
            .in2(_gnd_net_),
            .in3(N__40781),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48651),
            .ce(),
            .sr(N__48260));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_15_27_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_15_27_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_15_27_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_15_27_2  (
            .in0(N__40759),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40774),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_15_27_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_15_27_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_15_27_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_15_27_5  (
            .in0(N__41371),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41386),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_16_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_16_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_16_7_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_18_LC_16_7_1  (
            .in0(N__43317),
            .in1(N__43337),
            .in2(_gnd_net_),
            .in3(N__47056),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48789),
            .ce(N__46109),
            .sr(N__48123));
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_16_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_16_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_16_7_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_25_LC_16_7_2  (
            .in0(N__47055),
            .in1(N__45072),
            .in2(_gnd_net_),
            .in3(N__45056),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48789),
            .ce(N__46109),
            .sr(N__48123));
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_16_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_16_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_16_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_3_LC_16_7_7  (
            .in0(N__43520),
            .in1(N__43565),
            .in2(_gnd_net_),
            .in3(N__47057),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48789),
            .ce(N__46109),
            .sr(N__48123));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_16_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_16_8_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_16_8_0  (
            .in0(N__43177),
            .in1(N__43155),
            .in2(_gnd_net_),
            .in3(N__47052),
            .lcout(elapsed_time_ns_1_RNIDC91B_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_16_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_16_8_1 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_16_8_1  (
            .in0(N__44056),
            .in1(N__42907),
            .in2(_gnd_net_),
            .in3(N__46228),
            .lcout(\phase_controller_inst1.stoper_tr.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_16_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_16_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_16_8_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_16_8_3  (
            .in0(N__47054),
            .in1(N__44298),
            .in2(_gnd_net_),
            .in3(N__44257),
            .lcout(elapsed_time_ns_1_RNIIH91B_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_16_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_16_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_16_8_6  (
            .in0(N__44941),
            .in1(N__44919),
            .in2(_gnd_net_),
            .in3(N__47051),
            .lcout(elapsed_time_ns_1_RNIKJ91B_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_16_8_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_16_8_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_16_8_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_16_8_7  (
            .in0(N__47053),
            .in1(N__43272),
            .in2(_gnd_net_),
            .in3(N__43249),
            .lcout(elapsed_time_ns_1_RNIU8PBB_0_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_16_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_16_9_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_16_9_1  (
            .in0(N__43519),
            .in1(N__43560),
            .in2(_gnd_net_),
            .in3(N__46927),
            .lcout(elapsed_time_ns_1_RNIFE91B_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_16_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_16_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_16_9_2 .LUT_INIT=16'b0100110101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_16_9_2  (
            .in0(N__42025),
            .in1(N__41972),
            .in2(N__42005),
            .in3(N__46130),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_16_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_16_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_16_9_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_16_9_3  (
            .in0(N__43874),
            .in1(N__43828),
            .in2(_gnd_net_),
            .in3(N__46926),
            .lcout(elapsed_time_ns_1_RNI5GPBB_0_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_16_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_16_9_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_16_9_4  (
            .in0(N__46928),
            .in1(N__45003),
            .in2(_gnd_net_),
            .in3(N__44965),
            .lcout(elapsed_time_ns_1_RNIHG91B_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_16_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_16_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_16_9_5 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_16_9_5  (
            .in0(N__46129),
            .in1(N__42026),
            .in2(N__42004),
            .in3(N__41971),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_16_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_16_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_16_9_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_16_9_6  (
            .in0(N__46925),
            .in1(N__44877),
            .in2(_gnd_net_),
            .in3(N__44854),
            .lcout(elapsed_time_ns_1_RNIJI91B_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_16_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_16_9_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_16_9_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_16_9_7  (
            .in0(N__43499),
            .in1(N__43480),
            .in2(_gnd_net_),
            .in3(N__46929),
            .lcout(elapsed_time_ns_1_RNIGF91B_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_16_10_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_16_10_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_16_10_0  (
            .in0(N__43869),
            .in1(N__44231),
            .in2(_gnd_net_),
            .in3(N__41951),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_16_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_16_10_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_16_10_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_16_10_2  (
            .in0(N__41415),
            .in1(N__41944),
            .in2(_gnd_net_),
            .in3(N__41888),
            .lcout(elapsed_time_ns_1_RNIV1DN9_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_16_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_16_10_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_16_10_3  (
            .in0(_gnd_net_),
            .in1(N__44915),
            .in2(_gnd_net_),
            .in3(N__44849),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_16_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_16_10_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_16_10_4  (
            .in0(N__42122),
            .in1(N__44297),
            .in2(N__42137),
            .in3(N__45002),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_16_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_16_10_5 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_16_10_5  (
            .in0(N__46394),
            .in1(N__42566),
            .in2(N__42134),
            .in3(N__42131),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_16_10_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_16_10_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_16_10_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_16_10_6  (
            .in0(N__43405),
            .in1(_gnd_net_),
            .in2(N__42125),
            .in3(N__43384),
            .lcout(elapsed_time_ns_1_RNI2COBB_0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_16_11_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_16_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_16_11_0  (
            .in0(N__45976),
            .in1(N__42101),
            .in2(N__42077),
            .in3(N__44345),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_16_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_16_11_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_16_11_2  (
            .in0(N__46930),
            .in1(N__42115),
            .in2(_gnd_net_),
            .in3(N__42102),
            .lcout(elapsed_time_ns_1_RNIT6OBB_0_10),
            .ltout(elapsed_time_ns_1_RNIT6OBB_0_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_16_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_16_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_16_11_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_10_LC_16_11_3  (
            .in0(N__42103),
            .in1(_gnd_net_),
            .in2(N__42080),
            .in3(N__46931),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48751),
            .ce(N__46699),
            .sr(N__48145));
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_16_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_16_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_16_11_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_12_LC_16_11_7  (
            .in0(N__46936),
            .in1(N__42076),
            .in2(_gnd_net_),
            .in3(N__42050),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48751),
            .ce(N__46699),
            .sr(N__48145));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_16_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_16_12_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_16_12_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_16_12_0  (
            .in0(N__46975),
            .in1(N__45550),
            .in2(_gnd_net_),
            .in3(N__45523),
            .lcout(elapsed_time_ns_1_RNI2DPBB_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_16_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_16_12_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_16_12_2  (
            .in0(N__46974),
            .in1(N__42553),
            .in2(_gnd_net_),
            .in3(N__42488),
            .lcout(elapsed_time_ns_1_RNIV9PBB_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIIMJC3_28_LC_16_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIIMJC3_28_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIIMJC3_28_LC_16_12_4 .LUT_INIT=16'b1111101100111011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIIMJC3_28_LC_16_12_4  (
            .in0(N__45829),
            .in1(N__46246),
            .in2(N__45695),
            .in3(N__45632),
            .lcout(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_16_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_16_12_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_16_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42287),
            .in3(N__46190),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_16_12_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_16_12_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_16_12_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_16_12_6  (
            .in0(N__46976),
            .in1(N__46000),
            .in2(_gnd_net_),
            .in3(N__45975),
            .lcout(elapsed_time_ns_1_RNIU7OBB_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4_28_LC_16_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4_28_LC_16_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4_28_LC_16_12_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4_28_LC_16_12_7  (
            .in0(_gnd_net_),
            .in1(N__46191),
            .in2(_gnd_net_),
            .in3(N__42277),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_16_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_16_13_0 .LUT_INIT=16'b0010111100000010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_16_13_0  (
            .in0(N__42242),
            .in1(N__43789),
            .in2(N__43772),
            .in3(N__42233),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_16_13_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_16_13_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_16_13_1  (
            .in0(N__47083),
            .in1(N__42262),
            .in2(_gnd_net_),
            .in3(N__42165),
            .lcout(elapsed_time_ns_1_RNI3DOBB_0_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_16_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_16_13_4 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_16_13_4  (
            .in0(N__42241),
            .in1(N__43788),
            .in2(N__43771),
            .in3(N__42232),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_16_13_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_16_13_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_16_13_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_16_13_7  (
            .in0(N__47084),
            .in1(N__42220),
            .in2(_gnd_net_),
            .in3(N__42522),
            .lcout(elapsed_time_ns_1_RNI4EOBB_0_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_16_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_16_14_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_16_14_0  (
            .in0(N__42192),
            .in1(N__43358),
            .in2(N__42164),
            .in3(N__46319),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_16_14_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_16_14_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_16_14_1  (
            .in0(N__42533),
            .in1(N__42455),
            .in2(N__42569),
            .in3(N__42494),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_16_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_16_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_16_14_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_21_LC_16_14_6  (
            .in0(N__42554),
            .in1(N__42486),
            .in2(_gnd_net_),
            .in3(N__47082),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48721),
            .ce(N__46614),
            .sr(N__48171));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_16_15_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_16_15_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_16_15_1  (
            .in0(N__42418),
            .in1(_gnd_net_),
            .in2(N__47145),
            .in3(N__42445),
            .lcout(elapsed_time_ns_1_RNI7IPBB_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_16_15_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_16_15_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_16_15_2  (
            .in0(N__45029),
            .in1(N__42417),
            .in2(N__45785),
            .in3(N__46044),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_16_15_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_16_15_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_16_15_5  (
            .in0(N__44766),
            .in1(N__43299),
            .in2(N__43232),
            .in3(N__42512),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_16_15_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_16_15_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_16_15_7  (
            .in0(N__47298),
            .in1(N__45507),
            .in2(N__47195),
            .in3(N__42473),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_16_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_16_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_16_16_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_29_LC_16_16_3  (
            .in0(N__47081),
            .in1(N__42441),
            .in2(_gnd_net_),
            .in3(N__42413),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48702),
            .ce(N__46676),
            .sr(N__48190));
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_16_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_16_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_16_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_LC_16_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42384),
            .lcout(\phase_controller_inst1.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48694),
            .ce(),
            .sr(N__48199));
    defparam \phase_controller_inst1.start_timer_tr_LC_16_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_16_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_16_17_7 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_16_17_7  (
            .in0(N__42962),
            .in1(N__42677),
            .in2(N__44055),
            .in3(N__44563),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48694),
            .ce(),
            .sr(N__48199));
    defparam \delay_measurement_inst.stop_timer_tr_LC_16_18_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_16_18_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_tr_LC_16_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_16_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43966),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42722),
            .ce(),
            .sr(N__48207));
    defparam \phase_controller_inst1.state_RNIE87F_2_LC_16_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNIE87F_2_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNIE87F_2_LC_16_19_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.state_RNIE87F_2_LC_16_19_0  (
            .in0(N__44627),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42709),
            .lcout(\phase_controller_inst1.state_RNIE87FZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_16_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_16_19_4 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_RNO_0_LC_16_19_4  (
            .in0(N__42633),
            .in1(N__42708),
            .in2(N__44632),
            .in3(N__43057),
            .lcout(\phase_controller_inst1.start_timer_tr_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_1_LC_16_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_16_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_16_20_0 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \phase_controller_inst1.state_1_LC_16_20_0  (
            .in0(N__42634),
            .in1(N__43067),
            .in2(_gnd_net_),
            .in3(N__42667),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48678),
            .ce(),
            .sr(N__48220));
    defparam \phase_controller_inst1.T45_LC_16_22_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.T45_LC_16_22_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T45_LC_16_22_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \phase_controller_inst1.T45_LC_16_22_1  (
            .in0(_gnd_net_),
            .in1(N__42652),
            .in2(_gnd_net_),
            .in3(N__44578),
            .lcout(T45_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48668),
            .ce(),
            .sr(N__48231));
    defparam \phase_controller_inst1.state_0_LC_16_22_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_16_22_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_16_22_7 .LUT_INIT=16'b1111010001000100;
    LogicCell40 \phase_controller_inst1.state_0_LC_16_22_7  (
            .in0(N__46163),
            .in1(N__44579),
            .in2(N__42641),
            .in3(N__43069),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48668),
            .ce(),
            .sr(N__48231));
    defparam \phase_controller_inst1.T23_LC_16_23_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.T23_LC_16_23_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T23_LC_16_23_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \phase_controller_inst1.T23_LC_16_23_6  (
            .in0(_gnd_net_),
            .in1(N__42586),
            .in2(_gnd_net_),
            .in3(N__43068),
            .lcout(T23_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48664),
            .ce(),
            .sr(N__48236));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_16_24_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_16_24_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_16_24_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_16_24_0  (
            .in0(N__42869),
            .in1(N__42575),
            .in2(N__43103),
            .in3(N__42881),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_16_24_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_16_24_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_16_24_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_16_24_2  (
            .in0(N__42824),
            .in1(N__42860),
            .in2(N__42812),
            .in3(N__42851),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_16_24_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_16_24_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_16_24_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_16_24_3  (
            .in0(N__42890),
            .in1(N__42842),
            .in2(N__42797),
            .in3(N__42833),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_16_24_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_16_24_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_16_24_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_16_24_4  (
            .in0(_gnd_net_),
            .in1(N__42889),
            .in2(_gnd_net_),
            .in3(N__42880),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_16_24_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_16_24_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_16_24_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_16_24_5  (
            .in0(N__42773),
            .in1(N__42779),
            .in2(N__42872),
            .in3(N__42868),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_16_24_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_16_24_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_16_24_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_16_24_6  (
            .in0(N__44455),
            .in1(N__42859),
            .in2(N__44476),
            .in3(N__42850),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_16_24_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_16_24_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_16_24_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_16_24_7  (
            .in0(_gnd_net_),
            .in1(N__42841),
            .in2(_gnd_net_),
            .in3(N__42832),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_16_25_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_16_25_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_16_25_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_16_25_0  (
            .in0(N__42823),
            .in1(N__42808),
            .in2(N__42755),
            .in3(N__42790),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_16_25_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_16_25_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_16_25_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_16_25_1  (
            .in0(N__42740),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42730),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_16_25_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_16_25_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_16_25_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_16_25_2  (
            .in0(N__42772),
            .in1(N__43093),
            .in2(N__42758),
            .in3(N__42754),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_16_25_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_16_25_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_16_25_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_16_25_3  (
            .in0(N__42739),
            .in1(N__43123),
            .in2(N__43115),
            .in3(N__42731),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_16_25_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_16_25_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_16_25_4 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_16_25_4  (
            .in0(N__43124),
            .in1(N__43111),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_16_25_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_16_25_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_16_25_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_16_25_6  (
            .in0(N__44491),
            .in1(N__44509),
            .in2(N__43094),
            .in3(N__43079),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.S2_LC_16_30_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_16_30_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_16_30_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_16_30_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43073),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48647),
            .ce(),
            .sr(N__48272));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_17_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_17_7_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_17_7_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_17_7_3  (
            .in0(N__45076),
            .in1(N__45048),
            .in2(_gnd_net_),
            .in3(N__47065),
            .lcout(elapsed_time_ns_1_RNI3EPBB_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_17_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_17_7_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_17_7_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_17_7_6  (
            .in0(N__47066),
            .in1(N__44371),
            .in2(_gnd_net_),
            .in3(N__44349),
            .lcout(elapsed_time_ns_1_RNILK91B_0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_17_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_17_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_17_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_LC_17_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44057),
            .lcout(\phase_controller_inst1.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48790),
            .ce(),
            .sr(N__48124));
    defparam \phase_controller_inst1.state_4_LC_17_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_17_8_6 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_17_8_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.state_4_LC_17_8_6  (
            .in0(_gnd_net_),
            .in1(N__42999),
            .in2(_gnd_net_),
            .in3(N__42929),
            .lcout(phase_controller_inst1_state_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48790),
            .ce(),
            .sr(N__48124));
    defparam \phase_controller_inst1.stoper_tr.running_LC_17_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_LC_17_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.running_LC_17_8_7 .LUT_INIT=16'b1101010111110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_LC_17_8_7  (
            .in0(N__46238),
            .in1(N__46271),
            .in2(N__42908),
            .in3(N__46189),
            .lcout(\phase_controller_inst1.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48790),
            .ce(),
            .sr(N__48124));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_17_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_17_9_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_17_9_0  (
            .in0(N__43747),
            .in1(N__43723),
            .in2(N__44750),
            .in3(N__43283),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_17_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_17_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_17_9_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_17_9_1  (
            .in0(N__43282),
            .in1(N__43748),
            .in2(N__43727),
            .in3(N__44746),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_17_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_17_9_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_17_9_2  (
            .in0(N__44809),
            .in1(N__44788),
            .in2(_gnd_net_),
            .in3(N__46921),
            .lcout(elapsed_time_ns_1_RNI6GOBB_0_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_17_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_17_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_17_9_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_15_LC_17_9_4  (
            .in0(N__43401),
            .in1(N__43385),
            .in2(_gnd_net_),
            .in3(N__46924),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48784),
            .ce(N__46706),
            .sr(N__48130));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_17_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_17_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_17_9_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_17_9_6  (
            .in0(N__43318),
            .in1(N__43333),
            .in2(_gnd_net_),
            .in3(N__46922),
            .lcout(elapsed_time_ns_1_RNI5FOBB_0_18),
            .ltout(elapsed_time_ns_1_RNI5FOBB_0_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_17_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_17_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_17_9_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_18_LC_17_9_7  (
            .in0(N__46923),
            .in1(_gnd_net_),
            .in2(N__43322),
            .in3(N__43319),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48784),
            .ce(N__46706),
            .sr(N__48130));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_17_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_17_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_17_10_0 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_17_10_0  (
            .in0(N__43703),
            .in1(N__43192),
            .in2(N__43682),
            .in3(N__43205),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_17_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_17_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_17_10_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_20_LC_17_10_2  (
            .in0(N__43273),
            .in1(N__43250),
            .in2(_gnd_net_),
            .in3(N__46993),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48772),
            .ce(N__46675),
            .sr(N__48134));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_17_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_17_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_17_10_3 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_17_10_3  (
            .in0(N__43204),
            .in1(N__43681),
            .in2(N__43196),
            .in3(N__43702),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_17_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_17_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_17_10_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_1_LC_17_10_4  (
            .in0(N__43178),
            .in1(N__43156),
            .in2(_gnd_net_),
            .in3(N__46992),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48772),
            .ce(N__46675),
            .sr(N__48134));
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_17_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_17_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_17_10_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_2_LC_17_10_5  (
            .in0(N__46990),
            .in1(N__43617),
            .in2(_gnd_net_),
            .in3(N__43588),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48772),
            .ce(N__46675),
            .sr(N__48134));
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_17_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_17_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_17_10_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_3_LC_17_10_6  (
            .in0(N__43564),
            .in1(N__43518),
            .in2(_gnd_net_),
            .in3(N__46994),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48772),
            .ce(N__46675),
            .sr(N__48134));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_17_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_17_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_17_10_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_LC_17_10_7  (
            .in0(N__46991),
            .in1(N__43497),
            .in2(_gnd_net_),
            .in3(N__43481),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48772),
            .ce(N__46675),
            .sr(N__48134));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_17_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_17_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_17_11_0  (
            .in0(_gnd_net_),
            .in1(N__43442),
            .in2(N__44738),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_17_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_17_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_17_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_17_11_1  (
            .in0(N__46694),
            .in1(N__44687),
            .in2(_gnd_net_),
            .in3(N__43436),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__48764),
            .ce(),
            .sr(N__48140));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_17_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_17_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_17_11_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_17_11_2  (
            .in0(N__46601),
            .in1(N__44651),
            .in2(N__43433),
            .in3(N__43421),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__48764),
            .ce(),
            .sr(N__48140));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_17_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_17_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_17_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_17_11_3  (
            .in0(N__46695),
            .in1(N__45284),
            .in2(_gnd_net_),
            .in3(N__43418),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__48764),
            .ce(),
            .sr(N__48140));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_17_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_17_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_17_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_17_11_4  (
            .in0(N__46602),
            .in1(N__45266),
            .in2(_gnd_net_),
            .in3(N__43415),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__48764),
            .ce(),
            .sr(N__48140));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_17_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_17_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_17_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_17_11_5  (
            .in0(N__46696),
            .in1(N__45230),
            .in2(_gnd_net_),
            .in3(N__43412),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__48764),
            .ce(),
            .sr(N__48140));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_17_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_17_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_17_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_17_11_6  (
            .in0(N__46603),
            .in1(N__45203),
            .in2(_gnd_net_),
            .in3(N__43649),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__48764),
            .ce(),
            .sr(N__48140));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_17_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_17_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_17_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_17_11_7  (
            .in0(N__46697),
            .in1(N__45176),
            .in2(_gnd_net_),
            .in3(N__43646),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__48764),
            .ce(),
            .sr(N__48140));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_17_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_17_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_17_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_17_12_0  (
            .in0(N__46594),
            .in1(N__45145),
            .in2(_gnd_net_),
            .in3(N__43643),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_17_12_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__48752),
            .ce(),
            .sr(N__48146));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_17_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_17_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_17_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_17_12_1  (
            .in0(N__46604),
            .in1(N__45122),
            .in2(_gnd_net_),
            .in3(N__43640),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__48752),
            .ce(),
            .sr(N__48146));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_17_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_17_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_17_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_17_12_2  (
            .in0(N__46591),
            .in1(N__45089),
            .in2(_gnd_net_),
            .in3(N__43637),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__48752),
            .ce(),
            .sr(N__48146));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_17_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_17_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_17_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_17_12_3  (
            .in0(N__46605),
            .in1(N__45476),
            .in2(_gnd_net_),
            .in3(N__43634),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__48752),
            .ce(),
            .sr(N__48146));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_17_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_17_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_17_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_17_12_4  (
            .in0(N__46592),
            .in1(N__45455),
            .in2(_gnd_net_),
            .in3(N__43631),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__48752),
            .ce(),
            .sr(N__48146));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_17_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_17_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_17_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_17_12_5  (
            .in0(N__46606),
            .in1(N__45422),
            .in2(_gnd_net_),
            .in3(N__43628),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__48752),
            .ce(),
            .sr(N__48146));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_17_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_17_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_17_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_17_12_6  (
            .in0(N__46593),
            .in1(N__45392),
            .in2(_gnd_net_),
            .in3(N__43625),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__48752),
            .ce(),
            .sr(N__48146));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_12_7  (
            .in0(N__46607),
            .in1(N__43790),
            .in2(_gnd_net_),
            .in3(N__43775),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__48752),
            .ce(),
            .sr(N__48146));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_13_0  (
            .in0(N__46678),
            .in1(N__43770),
            .in2(_gnd_net_),
            .in3(N__43751),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_17_13_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__48740),
            .ce(),
            .sr(N__48155));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_17_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_17_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_17_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_17_13_1  (
            .in0(N__46682),
            .in1(N__43746),
            .in2(_gnd_net_),
            .in3(N__43730),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__48740),
            .ce(),
            .sr(N__48155));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_17_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_17_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_17_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_17_13_2  (
            .in0(N__46679),
            .in1(N__43722),
            .in2(_gnd_net_),
            .in3(N__43706),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(N__48740),
            .ce(),
            .sr(N__48155));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_17_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_17_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_17_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_17_13_3  (
            .in0(N__46683),
            .in1(N__43701),
            .in2(_gnd_net_),
            .in3(N__43685),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(N__48740),
            .ce(),
            .sr(N__48155));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_17_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_17_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_17_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_17_13_4  (
            .in0(N__46680),
            .in1(N__43677),
            .in2(_gnd_net_),
            .in3(N__43661),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ),
            .clk(N__48740),
            .ce(),
            .sr(N__48155));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_17_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_17_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_17_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_17_13_5  (
            .in0(N__46684),
            .in1(N__47395),
            .in2(_gnd_net_),
            .in3(N__43658),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ),
            .clk(N__48740),
            .ce(),
            .sr(N__48155));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_17_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_17_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_17_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_17_13_6  (
            .in0(N__46681),
            .in1(N__47371),
            .in2(_gnd_net_),
            .in3(N__43655),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ),
            .clk(N__48740),
            .ce(),
            .sr(N__48155));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_17_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_17_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_17_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_17_13_7  (
            .in0(N__46685),
            .in1(N__45578),
            .in2(_gnd_net_),
            .in3(N__43652),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ),
            .clk(N__48740),
            .ce(),
            .sr(N__48155));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_17_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_17_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_17_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_17_14_0  (
            .in0(N__46661),
            .in1(N__45610),
            .in2(_gnd_net_),
            .in3(N__43895),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_17_14_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ),
            .clk(N__48730),
            .ce(),
            .sr(N__48163));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_17_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_17_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_17_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_17_14_1  (
            .in0(N__46608),
            .in1(N__45873),
            .in2(_gnd_net_),
            .in3(N__43892),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ),
            .clk(N__48730),
            .ce(),
            .sr(N__48163));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_17_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_17_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_17_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_17_14_2  (
            .in0(N__46662),
            .in1(N__45895),
            .in2(_gnd_net_),
            .in3(N__43889),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ),
            .clk(N__48730),
            .ce(),
            .sr(N__48163));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_17_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_17_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_17_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_17_14_3  (
            .in0(N__46609),
            .in1(N__44198),
            .in2(_gnd_net_),
            .in3(N__43886),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ),
            .clk(N__48730),
            .ce(),
            .sr(N__48163));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_17_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_17_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_17_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_17_14_4  (
            .in0(N__46663),
            .in1(N__44164),
            .in2(_gnd_net_),
            .in3(N__43883),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ),
            .clk(N__48730),
            .ce(),
            .sr(N__48163));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_17_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_17_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_17_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_17_14_5  (
            .in0(N__46610),
            .in1(N__45713),
            .in2(_gnd_net_),
            .in3(N__43880),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ),
            .clk(N__48730),
            .ce(),
            .sr(N__48163));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_17_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_17_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_17_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_17_14_6  (
            .in0(N__46664),
            .in1(N__45733),
            .in2(_gnd_net_),
            .in3(N__43877),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48730),
            .ce(),
            .sr(N__48163));
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_17_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_17_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_17_15_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_27_LC_17_15_1  (
            .in0(N__47089),
            .in1(N__43873),
            .in2(_gnd_net_),
            .in3(N__43832),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48722),
            .ce(N__46657),
            .sr(N__48172));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_17_15_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_17_15_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_17_15_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_17_15_2  (
            .in0(N__44233),
            .in1(N__43801),
            .in2(_gnd_net_),
            .in3(N__47088),
            .lcout(elapsed_time_ns_1_RNI6HPBB_0_28),
            .ltout(elapsed_time_ns_1_RNI6HPBB_0_28_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_17_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_17_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_17_15_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_28_LC_17_15_3  (
            .in0(N__47090),
            .in1(_gnd_net_),
            .in2(N__44237),
            .in3(N__44234),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48722),
            .ce(N__46657),
            .sr(N__48172));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_17_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_17_15_4 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_17_15_4  (
            .in0(N__44146),
            .in1(N__44163),
            .in2(N__44183),
            .in3(N__44197),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_17_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_17_15_5 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_17_15_5  (
            .in0(N__44196),
            .in1(N__44179),
            .in2(N__44165),
            .in3(N__44147),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_17_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_17_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_17_15_7 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_17_15_7  (
            .in0(N__45911),
            .in1(N__45891),
            .in2(N__45874),
            .in3(N__45850),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_17_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_17_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_17_16_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_31_LC_17_16_6  (
            .in0(N__46396),
            .in1(N__46354),
            .in2(_gnd_net_),
            .in3(N__47106),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48711),
            .ce(N__46118),
            .sr(N__48180));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_17_17_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_17_17_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_17_17_3  (
            .in0(_gnd_net_),
            .in1(N__44000),
            .in2(_gnd_net_),
            .in3(N__44016),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_200_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_17_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_17_17_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_17_17_6  (
            .in0(_gnd_net_),
            .in1(N__46242),
            .in2(_gnd_net_),
            .in3(N__44042),
            .lcout(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_17_18_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_17_18_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_17_18_6 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_17_18_6  (
            .in0(N__44017),
            .in1(N__43995),
            .in2(_gnd_net_),
            .in3(N__43970),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_201_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.T12_LC_17_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.T12_LC_17_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T12_LC_17_19_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \phase_controller_inst1.T12_LC_17_19_0  (
            .in0(_gnd_net_),
            .in1(N__44590),
            .in2(_gnd_net_),
            .in3(N__44633),
            .lcout(T12_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48688),
            .ce(),
            .sr(N__48208));
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_17_22_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_17_22_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_17_22_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNI7NN7_0_LC_17_22_3  (
            .in0(_gnd_net_),
            .in1(N__46159),
            .in2(_gnd_net_),
            .in3(N__44577),
            .lcout(\phase_controller_inst1.state_RNI7NN7Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_17_24_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_17_24_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_17_24_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_17_24_3  (
            .in0(N__44543),
            .in1(N__44537),
            .in2(N__44531),
            .in3(N__44522),
            .lcout(\current_shift_inst.PI_CTRL.N_159 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_17_25_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_17_25_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_17_25_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_17_25_3  (
            .in0(N__44516),
            .in1(N__44498),
            .in2(N__44480),
            .in3(N__44459),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_17_25_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_17_25_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_17_25_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_17_25_4  (
            .in0(N__44444),
            .in1(N__44438),
            .in2(N__44432),
            .in3(N__44429),
            .lcout(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_17_26_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_17_26_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_17_26_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_17_26_4  (
            .in0(_gnd_net_),
            .in1(N__44419),
            .in2(_gnd_net_),
            .in3(N__44394),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_18_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_18_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_18_7_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_9_LC_18_7_4  (
            .in0(N__44367),
            .in1(N__44351),
            .in2(_gnd_net_),
            .in3(N__47138),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48802),
            .ce(N__46702),
            .sr(N__48121));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_18_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_18_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_18_8_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_LC_18_8_2  (
            .in0(N__44303),
            .in1(N__44258),
            .in2(_gnd_net_),
            .in3(N__47137),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48798),
            .ce(N__46698),
            .sr(N__48122));
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_18_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_18_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_18_9_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_25_LC_18_9_1  (
            .in0(N__45077),
            .in1(N__45055),
            .in2(_gnd_net_),
            .in3(N__47135),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48791),
            .ce(N__46687),
            .sr(N__48125));
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_18_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_18_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_18_9_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_5_LC_18_9_4  (
            .in0(N__47132),
            .in1(N__45008),
            .in2(_gnd_net_),
            .in3(N__44966),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48791),
            .ce(N__46687),
            .sr(N__48125));
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_18_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_18_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_18_9_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_8_LC_18_9_5  (
            .in0(N__44945),
            .in1(N__44921),
            .in2(_gnd_net_),
            .in3(N__47136),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48791),
            .ce(N__46687),
            .sr(N__48125));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_18_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_18_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_18_9_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_LC_18_9_6  (
            .in0(N__47133),
            .in1(N__44878),
            .in2(_gnd_net_),
            .in3(N__44855),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48791),
            .ce(N__46687),
            .sr(N__48125));
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_18_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_18_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_18_9_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_19_LC_18_9_7  (
            .in0(N__44805),
            .in1(N__44789),
            .in2(_gnd_net_),
            .in3(N__47134),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48791),
            .ce(N__46687),
            .sr(N__48125));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_18_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_18_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_18_10_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_18_10_0  (
            .in0(N__44734),
            .in1(N__44702),
            .in2(N__44696),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_18_10_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_18_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_18_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_18_10_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_18_10_1  (
            .in0(N__44686),
            .in1(N__44666),
            .in2(N__44675),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_18_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_18_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_18_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_18_10_2  (
            .in0(_gnd_net_),
            .in1(N__44639),
            .in2(N__44660),
            .in3(N__44650),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_18_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_18_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_18_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_18_10_3  (
            .in0(_gnd_net_),
            .in1(N__45272),
            .in2(N__45293),
            .in3(N__45283),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_18_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_18_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_18_10_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_18_10_4  (
            .in0(N__45265),
            .in1(N__45245),
            .in2(N__45254),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_18_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_18_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_18_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_18_10_5  (
            .in0(_gnd_net_),
            .in1(N__45239),
            .in2(N__45218),
            .in3(N__45229),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_18_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_18_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_18_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_18_10_6  (
            .in0(_gnd_net_),
            .in1(N__45209),
            .in2(N__45191),
            .in3(N__45202),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_18_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_18_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_18_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_18_10_7  (
            .in0(_gnd_net_),
            .in1(N__45182),
            .in2(N__45164),
            .in3(N__45175),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_18_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_18_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_18_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_18_11_0  (
            .in0(_gnd_net_),
            .in1(N__45155),
            .in2(N__45131),
            .in3(N__45146),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_18_11_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_18_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_18_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_18_11_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_18_11_1  (
            .in0(N__45121),
            .in1(N__45110),
            .in2(N__45101),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_18_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_18_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_18_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_18_11_2  (
            .in0(_gnd_net_),
            .in1(N__45491),
            .in2(N__45944),
            .in3(N__45088),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_18_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_18_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_18_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_18_11_3  (
            .in0(_gnd_net_),
            .in1(N__45485),
            .in2(N__45464),
            .in3(N__45475),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_18_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_18_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_18_11_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_18_11_4  (
            .in0(N__45454),
            .in1(N__45443),
            .in2(N__45431),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_18_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_18_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_18_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_18_11_5  (
            .in0(_gnd_net_),
            .in1(N__45680),
            .in2(N__45410),
            .in3(N__45421),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_18_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_18_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_18_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_18_11_6  (
            .in0(_gnd_net_),
            .in1(N__45401),
            .in2(N__45380),
            .in3(N__45391),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_18_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_18_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_18_11_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_18_11_7  (
            .in0(_gnd_net_),
            .in1(N__45368),
            .in2(N__45356),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_18_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_18_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_18_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_18_12_0  (
            .in0(_gnd_net_),
            .in1(N__45341),
            .in2(N__45329),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_12_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_18_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_18_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_18_12_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_18_12_1  (
            .in0(_gnd_net_),
            .in1(N__45314),
            .in2(N__45305),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_18_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_18_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_18_12_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_18_12_2  (
            .in0(_gnd_net_),
            .in1(N__47357),
            .in2(N__45932),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_18_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_18_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_18_12_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_18_12_3  (
            .in0(_gnd_net_),
            .in1(N__45617),
            .in2(N__45563),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_18_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_18_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_18_12_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_18_12_4  (
            .in0(_gnd_net_),
            .in1(N__45836),
            .in2(N__45671),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_18_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_18_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_18_12_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_18_12_5  (
            .in0(_gnd_net_),
            .in1(N__45656),
            .in2(N__45647),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_18_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_18_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_18_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_18_12_6  (
            .in0(_gnd_net_),
            .in1(N__45755),
            .in2(N__45830),
            .in3(N__45623),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_18_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_18_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_18_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_18_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45620),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_18_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_18_13_0 .LUT_INIT=16'b0100111100000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_18_13_0  (
            .in0(N__45577),
            .in1(N__45920),
            .in2(N__45611),
            .in3(N__45592),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_18_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_18_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_18_13_1 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_18_13_1  (
            .in0(N__45919),
            .in1(N__45606),
            .in2(N__45593),
            .in3(N__45576),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_18_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_18_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_18_13_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_24_LC_18_13_5  (
            .in0(N__47130),
            .in1(N__45551),
            .in2(_gnd_net_),
            .in3(N__45527),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48753),
            .ce(N__46665),
            .sr(N__48147));
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_18_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_18_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_18_13_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_26_LC_18_13_6  (
            .in0(N__46028),
            .in1(N__46068),
            .in2(_gnd_net_),
            .in3(N__47131),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48753),
            .ce(N__46665),
            .sr(N__48147));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_18_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_18_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_18_13_7 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_18_13_7  (
            .in0(N__45907),
            .in1(N__45896),
            .in2(N__45875),
            .in3(N__45851),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_0_30_LC_18_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_0_30_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_0_30_LC_18_14_0 .LUT_INIT=16'b0000110010001110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_0_30_LC_18_14_0  (
            .in0(N__45745),
            .in1(N__45728),
            .in2(N__46414),
            .in3(N__45711),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_18_14_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_18_14_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_18_14_1  (
            .in0(N__45786),
            .in1(N__45802),
            .in2(_gnd_net_),
            .in3(N__47123),
            .lcout(elapsed_time_ns_1_RNIVAQBB_0_30),
            .ltout(elapsed_time_ns_1_RNIVAQBB_0_30_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_18_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_18_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_18_14_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_30_LC_18_14_2  (
            .in0(N__47124),
            .in1(_gnd_net_),
            .in2(N__45791),
            .in3(N__45787),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48741),
            .ce(N__46615),
            .sr(N__48156));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_18_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_18_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_18_14_3 .LUT_INIT=16'b1111001101110001;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_18_14_3  (
            .in0(N__45712),
            .in1(N__46413),
            .in2(N__45734),
            .in3(N__45746),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_30_LC_18_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_30_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_30_LC_18_14_6 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_30_LC_18_14_6  (
            .in0(N__45744),
            .in1(N__45729),
            .in2(N__46415),
            .in3(N__45710),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_df30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_18_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_18_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_18_15_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_14_LC_18_15_1  (
            .in0(N__46287),
            .in1(N__46335),
            .in2(_gnd_net_),
            .in3(N__47161),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48731),
            .ce(N__46589),
            .sr(N__48164));
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_18_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_18_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_18_15_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_31_LC_18_15_6  (
            .in0(N__47160),
            .in1(N__46397),
            .in2(_gnd_net_),
            .in3(N__46353),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48731),
            .ce(N__46589),
            .sr(N__48164));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_18_16_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_18_16_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_18_16_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_18_16_5  (
            .in0(N__46355),
            .in1(N__46395),
            .in2(_gnd_net_),
            .in3(N__47140),
            .lcout(elapsed_time_ns_1_RNI0CQBB_0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_18_16_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_18_16_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_18_16_6  (
            .in0(N__47139),
            .in1(N__46291),
            .in2(_gnd_net_),
            .in3(N__46336),
            .lcout(elapsed_time_ns_1_RNI1BOBB_0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_18_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_18_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_18_17_4 .LUT_INIT=16'b1101000011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_18_17_4  (
            .in0(N__46267),
            .in1(N__46149),
            .in2(N__46253),
            .in3(N__46201),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48712),
            .ce(),
            .sr(N__48181));
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_20_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_20_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_20_9_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_26_LC_20_9_5  (
            .in0(N__47163),
            .in1(N__46020),
            .in2(_gnd_net_),
            .in3(N__46076),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48803),
            .ce(N__46117),
            .sr(N__48126));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_20_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_20_10_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_20_10_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_20_10_4  (
            .in0(N__46024),
            .in1(N__46075),
            .in2(_gnd_net_),
            .in3(N__46977),
            .lcout(elapsed_time_ns_1_RNI4FPBB_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_20_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_20_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_20_11_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_11_LC_20_11_3  (
            .in0(N__47162),
            .in1(N__46004),
            .in2(_gnd_net_),
            .in3(N__45980),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48792),
            .ce(N__46700),
            .sr(N__48135));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_20_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_20_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_20_12_0 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_20_12_0  (
            .in0(N__47282),
            .in1(N__46715),
            .in2(N__47405),
            .in3(N__47380),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_20_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_20_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_20_12_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_20_12_1  (
            .in0(N__46714),
            .in1(N__47404),
            .in2(N__47381),
            .in3(N__47281),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_20_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_20_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_20_12_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_20_12_2  (
            .in0(N__47346),
            .in1(N__47323),
            .in2(_gnd_net_),
            .in3(N__47147),
            .lcout(elapsed_time_ns_1_RNI1CPBB_0_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_20_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_20_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_20_12_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_20_12_4  (
            .in0(N__47205),
            .in1(N__47230),
            .in2(_gnd_net_),
            .in3(N__47146),
            .lcout(elapsed_time_ns_1_RNI0BPBB_0_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_20_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_20_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_20_15_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_23_LC_20_15_6  (
            .in0(N__47347),
            .in1(N__47324),
            .in2(_gnd_net_),
            .in3(N__47165),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48754),
            .ce(N__46590),
            .sr(N__48165));
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_20_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_20_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_20_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_0_LC_20_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47270),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48713),
            .ce(),
            .sr(N__48200));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_20_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_20_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_20_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_20_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47240),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48695),
            .ce(),
            .sr(N__48214));
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_21_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_21_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_21_12_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_22_LC_21_12_1  (
            .in0(N__47226),
            .in1(N__47210),
            .in2(_gnd_net_),
            .in3(N__47164),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48793),
            .ce(N__46686),
            .sr(N__48148));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_22_23_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_22_23_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_22_23_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_22_23_2  (
            .in0(N__49177),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47691),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_22_23_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_22_23_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_22_23_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_22_23_5  (
            .in0(_gnd_net_),
            .in1(N__48900),
            .in2(_gnd_net_),
            .in3(N__49176),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_22_23_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_22_23_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_22_23_6 .LUT_INIT=16'b1010111110101011;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_LC_22_23_6  (
            .in0(N__47411),
            .in1(N__47573),
            .in2(N__49094),
            .in3(N__47780),
            .lcout(\pwm_generator_inst.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_22_24_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_22_24_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_22_24_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_22_24_1  (
            .in0(N__49234),
            .in1(N__47501),
            .in2(N__48907),
            .in3(N__47758),
            .lcout(\current_shift_inst.PI_CTRL.N_27 ),
            .ltout(\current_shift_inst.PI_CTRL.N_27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_22_24_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_22_24_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_22_24_2 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_22_24_2  (
            .in0(N__48962),
            .in1(N__47486),
            .in2(N__47495),
            .in3(N__48851),
            .lcout(\current_shift_inst.PI_CTRL.N_96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_22_24_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_22_24_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_22_24_5 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_22_24_5  (
            .in0(N__49233),
            .in1(N__47757),
            .in2(N__47705),
            .in3(N__47492),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_22_24_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_22_24_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_22_24_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_22_24_7  (
            .in0(_gnd_net_),
            .in1(N__49116),
            .in2(_gnd_net_),
            .in3(N__47605),
            .lcout(\current_shift_inst.PI_CTRL.N_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_23_23_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_23_23_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_23_23_0 .LUT_INIT=16'b0000000010101110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_23_23_0  (
            .in0(N__49300),
            .in1(N__47620),
            .in2(N__49066),
            .in3(N__47609),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_23_23_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_23_23_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_23_23_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_23_23_1  (
            .in0(N__47665),
            .in1(N__48827),
            .in2(N__49208),
            .in3(N__47722),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_23_23_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_23_23_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_23_23_2 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_LC_23_23_2  (
            .in0(N__49160),
            .in1(N__47572),
            .in2(N__47480),
            .in3(N__49087),
            .lcout(\pwm_generator_inst.N_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_23_23_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_23_23_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_23_23_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_23_23_5  (
            .in0(_gnd_net_),
            .in1(N__47721),
            .in2(_gnd_net_),
            .in3(N__49159),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_23_23_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_23_23_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_23_23_6 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_3_LC_23_23_6  (
            .in0(N__48826),
            .in1(N__47664),
            .in2(N__47414),
            .in3(N__49203),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_23_23_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_23_23_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_23_23_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pwm_generator_inst.un1_duty_inputlto2_LC_23_23_7  (
            .in0(N__47635),
            .in1(N__49345),
            .in2(_gnd_net_),
            .in3(N__49252),
            .lcout(\pwm_generator_inst.un1_duty_inputlt3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_23_24_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_23_24_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_23_24_1 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_23_24_1  (
            .in0(N__48959),
            .in1(N__49125),
            .in2(_gnd_net_),
            .in3(N__47772),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_23_24_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_23_24_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_23_24_3 .LUT_INIT=16'b0101000101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_23_24_3  (
            .in0(N__48961),
            .in1(N__47774),
            .in2(N__49065),
            .in3(N__49126),
            .lcout(\current_shift_inst.PI_CTRL.N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_23_24_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_23_24_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_23_24_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_23_24_4  (
            .in0(N__47773),
            .in1(N__49050),
            .in2(_gnd_net_),
            .in3(N__48960),
            .lcout(\current_shift_inst.PI_CTRL.N_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_24_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_24_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_24_22_2 .LUT_INIT=16'b1111010001010100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_24_22_2  (
            .in0(N__48980),
            .in1(N__49062),
            .in2(N__47762),
            .in3(N__48872),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48723),
            .ce(),
            .sr(N__48241));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_24_23_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_24_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_24_23_0 .LUT_INIT=16'b1111010001010100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_24_23_0  (
            .in0(N__48979),
            .in1(N__49064),
            .in2(N__47704),
            .in3(N__48871),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48714),
            .ce(),
            .sr(N__48246));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_24_23_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_24_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_24_23_1 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_24_23_1  (
            .in0(N__49329),
            .in1(N__49317),
            .in2(N__49288),
            .in3(N__47648),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48714),
            .ce(),
            .sr(N__48246));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_24_23_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_24_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_24_23_2 .LUT_INIT=16'b1111111101010001;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_24_23_2  (
            .in0(N__49316),
            .in1(N__47621),
            .in2(N__49067),
            .in3(N__47604),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48714),
            .ce(),
            .sr(N__48246));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_24_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_24_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_24_23_4 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_24_23_4  (
            .in0(N__49281),
            .in1(N__49361),
            .in2(N__49319),
            .in3(N__49330),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48714),
            .ce(),
            .sr(N__48246));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_24_23_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_24_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_24_23_5 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_24_23_5  (
            .in0(N__49331),
            .in1(N__49318),
            .in2(N__49289),
            .in3(N__49268),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48714),
            .ce(),
            .sr(N__48246));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_24_23_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_24_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_24_23_6 .LUT_INIT=16'b1111010001010100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_24_23_6  (
            .in0(N__48978),
            .in1(N__49063),
            .in2(N__49238),
            .in3(N__48870),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48714),
            .ce(),
            .sr(N__48246));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_24_24_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_24_24_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_24_24_0 .LUT_INIT=16'b1111001000110010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_24_24_0  (
            .in0(N__49054),
            .in1(N__48976),
            .in2(N__49187),
            .in3(N__48867),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48703),
            .ce(),
            .sr(N__48254));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_24_24_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_24_24_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_24_24_2 .LUT_INIT=16'b0101000101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_24_24_2  (
            .in0(N__49145),
            .in1(N__49139),
            .in2(N__49130),
            .in3(N__48869),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48703),
            .ce(),
            .sr(N__48254));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_24_24_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_24_24_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_24_24_6 .LUT_INIT=16'b1111001000110010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_24_24_6  (
            .in0(N__49055),
            .in1(N__48977),
            .in2(N__48908),
            .in3(N__48868),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48703),
            .ce(),
            .sr(N__48254));
endmodule // MAIN
