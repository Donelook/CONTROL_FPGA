-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 18 2025 23:48:52

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    start_stop : in std_logic;
    s2_phy : out std_logic;
    T23 : out std_logic;
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    T45 : out std_logic;
    T12 : out std_logic;
    s4_phy : out std_logic;
    rgb_g : out std_logic;
    T01 : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__50616\ : std_logic;
signal \N__50615\ : std_logic;
signal \N__50614\ : std_logic;
signal \N__50605\ : std_logic;
signal \N__50604\ : std_logic;
signal \N__50603\ : std_logic;
signal \N__50596\ : std_logic;
signal \N__50595\ : std_logic;
signal \N__50594\ : std_logic;
signal \N__50587\ : std_logic;
signal \N__50586\ : std_logic;
signal \N__50585\ : std_logic;
signal \N__50578\ : std_logic;
signal \N__50577\ : std_logic;
signal \N__50576\ : std_logic;
signal \N__50569\ : std_logic;
signal \N__50568\ : std_logic;
signal \N__50567\ : std_logic;
signal \N__50560\ : std_logic;
signal \N__50559\ : std_logic;
signal \N__50558\ : std_logic;
signal \N__50551\ : std_logic;
signal \N__50550\ : std_logic;
signal \N__50549\ : std_logic;
signal \N__50542\ : std_logic;
signal \N__50541\ : std_logic;
signal \N__50540\ : std_logic;
signal \N__50533\ : std_logic;
signal \N__50532\ : std_logic;
signal \N__50531\ : std_logic;
signal \N__50524\ : std_logic;
signal \N__50523\ : std_logic;
signal \N__50522\ : std_logic;
signal \N__50515\ : std_logic;
signal \N__50514\ : std_logic;
signal \N__50513\ : std_logic;
signal \N__50506\ : std_logic;
signal \N__50505\ : std_logic;
signal \N__50504\ : std_logic;
signal \N__50497\ : std_logic;
signal \N__50496\ : std_logic;
signal \N__50495\ : std_logic;
signal \N__50488\ : std_logic;
signal \N__50487\ : std_logic;
signal \N__50486\ : std_logic;
signal \N__50479\ : std_logic;
signal \N__50478\ : std_logic;
signal \N__50477\ : std_logic;
signal \N__50470\ : std_logic;
signal \N__50469\ : std_logic;
signal \N__50468\ : std_logic;
signal \N__50451\ : std_logic;
signal \N__50448\ : std_logic;
signal \N__50447\ : std_logic;
signal \N__50444\ : std_logic;
signal \N__50441\ : std_logic;
signal \N__50436\ : std_logic;
signal \N__50433\ : std_logic;
signal \N__50430\ : std_logic;
signal \N__50427\ : std_logic;
signal \N__50424\ : std_logic;
signal \N__50421\ : std_logic;
signal \N__50420\ : std_logic;
signal \N__50417\ : std_logic;
signal \N__50416\ : std_logic;
signal \N__50413\ : std_logic;
signal \N__50410\ : std_logic;
signal \N__50407\ : std_logic;
signal \N__50400\ : std_logic;
signal \N__50399\ : std_logic;
signal \N__50396\ : std_logic;
signal \N__50395\ : std_logic;
signal \N__50394\ : std_logic;
signal \N__50393\ : std_logic;
signal \N__50392\ : std_logic;
signal \N__50391\ : std_logic;
signal \N__50390\ : std_logic;
signal \N__50387\ : std_logic;
signal \N__50386\ : std_logic;
signal \N__50385\ : std_logic;
signal \N__50384\ : std_logic;
signal \N__50383\ : std_logic;
signal \N__50376\ : std_logic;
signal \N__50371\ : std_logic;
signal \N__50368\ : std_logic;
signal \N__50363\ : std_logic;
signal \N__50360\ : std_logic;
signal \N__50359\ : std_logic;
signal \N__50356\ : std_logic;
signal \N__50353\ : std_logic;
signal \N__50350\ : std_logic;
signal \N__50349\ : std_logic;
signal \N__50348\ : std_logic;
signal \N__50345\ : std_logic;
signal \N__50342\ : std_logic;
signal \N__50337\ : std_logic;
signal \N__50334\ : std_logic;
signal \N__50331\ : std_logic;
signal \N__50326\ : std_logic;
signal \N__50319\ : std_logic;
signal \N__50316\ : std_logic;
signal \N__50309\ : std_logic;
signal \N__50306\ : std_logic;
signal \N__50295\ : std_logic;
signal \N__50292\ : std_logic;
signal \N__50289\ : std_logic;
signal \N__50286\ : std_logic;
signal \N__50285\ : std_logic;
signal \N__50284\ : std_logic;
signal \N__50281\ : std_logic;
signal \N__50280\ : std_logic;
signal \N__50279\ : std_logic;
signal \N__50278\ : std_logic;
signal \N__50277\ : std_logic;
signal \N__50276\ : std_logic;
signal \N__50273\ : std_logic;
signal \N__50270\ : std_logic;
signal \N__50267\ : std_logic;
signal \N__50264\ : std_logic;
signal \N__50263\ : std_logic;
signal \N__50262\ : std_logic;
signal \N__50261\ : std_logic;
signal \N__50260\ : std_logic;
signal \N__50259\ : std_logic;
signal \N__50252\ : std_logic;
signal \N__50251\ : std_logic;
signal \N__50250\ : std_logic;
signal \N__50249\ : std_logic;
signal \N__50248\ : std_logic;
signal \N__50247\ : std_logic;
signal \N__50246\ : std_logic;
signal \N__50245\ : std_logic;
signal \N__50244\ : std_logic;
signal \N__50243\ : std_logic;
signal \N__50242\ : std_logic;
signal \N__50241\ : std_logic;
signal \N__50240\ : std_logic;
signal \N__50239\ : std_logic;
signal \N__50238\ : std_logic;
signal \N__50237\ : std_logic;
signal \N__50234\ : std_logic;
signal \N__50231\ : std_logic;
signal \N__50226\ : std_logic;
signal \N__50223\ : std_logic;
signal \N__50214\ : std_logic;
signal \N__50211\ : std_logic;
signal \N__50208\ : std_logic;
signal \N__50201\ : std_logic;
signal \N__50192\ : std_logic;
signal \N__50183\ : std_logic;
signal \N__50174\ : std_logic;
signal \N__50171\ : std_logic;
signal \N__50170\ : std_logic;
signal \N__50167\ : std_logic;
signal \N__50164\ : std_logic;
signal \N__50163\ : std_logic;
signal \N__50162\ : std_logic;
signal \N__50161\ : std_logic;
signal \N__50160\ : std_logic;
signal \N__50159\ : std_logic;
signal \N__50158\ : std_logic;
signal \N__50157\ : std_logic;
signal \N__50156\ : std_logic;
signal \N__50153\ : std_logic;
signal \N__50150\ : std_logic;
signal \N__50137\ : std_logic;
signal \N__50134\ : std_logic;
signal \N__50131\ : std_logic;
signal \N__50126\ : std_logic;
signal \N__50117\ : std_logic;
signal \N__50108\ : std_logic;
signal \N__50101\ : std_logic;
signal \N__50098\ : std_logic;
signal \N__50087\ : std_logic;
signal \N__50082\ : std_logic;
signal \N__50081\ : std_logic;
signal \N__50078\ : std_logic;
signal \N__50075\ : std_logic;
signal \N__50074\ : std_logic;
signal \N__50071\ : std_logic;
signal \N__50068\ : std_logic;
signal \N__50065\ : std_logic;
signal \N__50058\ : std_logic;
signal \N__50055\ : std_logic;
signal \N__50054\ : std_logic;
signal \N__50051\ : std_logic;
signal \N__50048\ : std_logic;
signal \N__50045\ : std_logic;
signal \N__50042\ : std_logic;
signal \N__50037\ : std_logic;
signal \N__50036\ : std_logic;
signal \N__50033\ : std_logic;
signal \N__50030\ : std_logic;
signal \N__50029\ : std_logic;
signal \N__50026\ : std_logic;
signal \N__50023\ : std_logic;
signal \N__50020\ : std_logic;
signal \N__50013\ : std_logic;
signal \N__50010\ : std_logic;
signal \N__50009\ : std_logic;
signal \N__50008\ : std_logic;
signal \N__50005\ : std_logic;
signal \N__50000\ : std_logic;
signal \N__49997\ : std_logic;
signal \N__49994\ : std_logic;
signal \N__49989\ : std_logic;
signal \N__49988\ : std_logic;
signal \N__49987\ : std_logic;
signal \N__49986\ : std_logic;
signal \N__49985\ : std_logic;
signal \N__49974\ : std_logic;
signal \N__49971\ : std_logic;
signal \N__49968\ : std_logic;
signal \N__49967\ : std_logic;
signal \N__49964\ : std_logic;
signal \N__49963\ : std_logic;
signal \N__49962\ : std_logic;
signal \N__49961\ : std_logic;
signal \N__49958\ : std_logic;
signal \N__49955\ : std_logic;
signal \N__49952\ : std_logic;
signal \N__49951\ : std_logic;
signal \N__49948\ : std_logic;
signal \N__49943\ : std_logic;
signal \N__49940\ : std_logic;
signal \N__49937\ : std_logic;
signal \N__49934\ : std_logic;
signal \N__49931\ : std_logic;
signal \N__49928\ : std_logic;
signal \N__49925\ : std_logic;
signal \N__49922\ : std_logic;
signal \N__49919\ : std_logic;
signal \N__49912\ : std_logic;
signal \N__49905\ : std_logic;
signal \N__49904\ : std_logic;
signal \N__49901\ : std_logic;
signal \N__49900\ : std_logic;
signal \N__49897\ : std_logic;
signal \N__49894\ : std_logic;
signal \N__49893\ : std_logic;
signal \N__49890\ : std_logic;
signal \N__49889\ : std_logic;
signal \N__49888\ : std_logic;
signal \N__49887\ : std_logic;
signal \N__49886\ : std_logic;
signal \N__49883\ : std_logic;
signal \N__49880\ : std_logic;
signal \N__49877\ : std_logic;
signal \N__49876\ : std_logic;
signal \N__49875\ : std_logic;
signal \N__49874\ : std_logic;
signal \N__49871\ : std_logic;
signal \N__49866\ : std_logic;
signal \N__49865\ : std_logic;
signal \N__49864\ : std_logic;
signal \N__49863\ : std_logic;
signal \N__49862\ : std_logic;
signal \N__49861\ : std_logic;
signal \N__49860\ : std_logic;
signal \N__49857\ : std_logic;
signal \N__49854\ : std_logic;
signal \N__49849\ : std_logic;
signal \N__49846\ : std_logic;
signal \N__49845\ : std_logic;
signal \N__49842\ : std_logic;
signal \N__49841\ : std_logic;
signal \N__49840\ : std_logic;
signal \N__49839\ : std_logic;
signal \N__49836\ : std_logic;
signal \N__49833\ : std_logic;
signal \N__49828\ : std_logic;
signal \N__49825\ : std_logic;
signal \N__49822\ : std_logic;
signal \N__49821\ : std_logic;
signal \N__49820\ : std_logic;
signal \N__49819\ : std_logic;
signal \N__49818\ : std_logic;
signal \N__49817\ : std_logic;
signal \N__49816\ : std_logic;
signal \N__49815\ : std_logic;
signal \N__49814\ : std_logic;
signal \N__49813\ : std_logic;
signal \N__49806\ : std_logic;
signal \N__49801\ : std_logic;
signal \N__49798\ : std_logic;
signal \N__49795\ : std_logic;
signal \N__49792\ : std_logic;
signal \N__49783\ : std_logic;
signal \N__49778\ : std_logic;
signal \N__49775\ : std_logic;
signal \N__49772\ : std_logic;
signal \N__49761\ : std_logic;
signal \N__49758\ : std_logic;
signal \N__49755\ : std_logic;
signal \N__49746\ : std_logic;
signal \N__49743\ : std_logic;
signal \N__49716\ : std_logic;
signal \N__49715\ : std_logic;
signal \N__49712\ : std_logic;
signal \N__49711\ : std_logic;
signal \N__49710\ : std_logic;
signal \N__49709\ : std_logic;
signal \N__49706\ : std_logic;
signal \N__49705\ : std_logic;
signal \N__49702\ : std_logic;
signal \N__49701\ : std_logic;
signal \N__49700\ : std_logic;
signal \N__49697\ : std_logic;
signal \N__49696\ : std_logic;
signal \N__49693\ : std_logic;
signal \N__49692\ : std_logic;
signal \N__49691\ : std_logic;
signal \N__49690\ : std_logic;
signal \N__49687\ : std_logic;
signal \N__49686\ : std_logic;
signal \N__49685\ : std_logic;
signal \N__49684\ : std_logic;
signal \N__49683\ : std_logic;
signal \N__49682\ : std_logic;
signal \N__49681\ : std_logic;
signal \N__49680\ : std_logic;
signal \N__49679\ : std_logic;
signal \N__49678\ : std_logic;
signal \N__49675\ : std_logic;
signal \N__49672\ : std_logic;
signal \N__49669\ : std_logic;
signal \N__49666\ : std_logic;
signal \N__49663\ : std_logic;
signal \N__49650\ : std_logic;
signal \N__49645\ : std_logic;
signal \N__49634\ : std_logic;
signal \N__49627\ : std_logic;
signal \N__49608\ : std_logic;
signal \N__49607\ : std_logic;
signal \N__49606\ : std_logic;
signal \N__49603\ : std_logic;
signal \N__49600\ : std_logic;
signal \N__49599\ : std_logic;
signal \N__49598\ : std_logic;
signal \N__49597\ : std_logic;
signal \N__49596\ : std_logic;
signal \N__49589\ : std_logic;
signal \N__49586\ : std_logic;
signal \N__49585\ : std_logic;
signal \N__49584\ : std_logic;
signal \N__49583\ : std_logic;
signal \N__49582\ : std_logic;
signal \N__49581\ : std_logic;
signal \N__49580\ : std_logic;
signal \N__49579\ : std_logic;
signal \N__49578\ : std_logic;
signal \N__49577\ : std_logic;
signal \N__49576\ : std_logic;
signal \N__49575\ : std_logic;
signal \N__49574\ : std_logic;
signal \N__49571\ : std_logic;
signal \N__49568\ : std_logic;
signal \N__49567\ : std_logic;
signal \N__49566\ : std_logic;
signal \N__49565\ : std_logic;
signal \N__49564\ : std_logic;
signal \N__49561\ : std_logic;
signal \N__49558\ : std_logic;
signal \N__49545\ : std_logic;
signal \N__49542\ : std_logic;
signal \N__49539\ : std_logic;
signal \N__49538\ : std_logic;
signal \N__49537\ : std_logic;
signal \N__49534\ : std_logic;
signal \N__49527\ : std_logic;
signal \N__49524\ : std_logic;
signal \N__49517\ : std_logic;
signal \N__49510\ : std_logic;
signal \N__49507\ : std_logic;
signal \N__49502\ : std_logic;
signal \N__49499\ : std_logic;
signal \N__49498\ : std_logic;
signal \N__49491\ : std_logic;
signal \N__49486\ : std_logic;
signal \N__49483\ : std_logic;
signal \N__49480\ : std_logic;
signal \N__49475\ : std_logic;
signal \N__49470\ : std_logic;
signal \N__49469\ : std_logic;
signal \N__49468\ : std_logic;
signal \N__49467\ : std_logic;
signal \N__49466\ : std_logic;
signal \N__49465\ : std_logic;
signal \N__49464\ : std_logic;
signal \N__49461\ : std_logic;
signal \N__49460\ : std_logic;
signal \N__49459\ : std_logic;
signal \N__49458\ : std_logic;
signal \N__49455\ : std_logic;
signal \N__49452\ : std_logic;
signal \N__49451\ : std_logic;
signal \N__49446\ : std_logic;
signal \N__49441\ : std_logic;
signal \N__49432\ : std_logic;
signal \N__49427\ : std_logic;
signal \N__49424\ : std_logic;
signal \N__49421\ : std_logic;
signal \N__49416\ : std_logic;
signal \N__49411\ : std_logic;
signal \N__49408\ : std_logic;
signal \N__49401\ : std_logic;
signal \N__49398\ : std_logic;
signal \N__49383\ : std_logic;
signal \N__49382\ : std_logic;
signal \N__49381\ : std_logic;
signal \N__49378\ : std_logic;
signal \N__49375\ : std_logic;
signal \N__49374\ : std_logic;
signal \N__49373\ : std_logic;
signal \N__49372\ : std_logic;
signal \N__49369\ : std_logic;
signal \N__49368\ : std_logic;
signal \N__49367\ : std_logic;
signal \N__49366\ : std_logic;
signal \N__49365\ : std_logic;
signal \N__49364\ : std_logic;
signal \N__49361\ : std_logic;
signal \N__49358\ : std_logic;
signal \N__49351\ : std_logic;
signal \N__49348\ : std_logic;
signal \N__49343\ : std_logic;
signal \N__49336\ : std_logic;
signal \N__49331\ : std_logic;
signal \N__49326\ : std_logic;
signal \N__49317\ : std_logic;
signal \N__49316\ : std_logic;
signal \N__49315\ : std_logic;
signal \N__49312\ : std_logic;
signal \N__49309\ : std_logic;
signal \N__49306\ : std_logic;
signal \N__49299\ : std_logic;
signal \N__49298\ : std_logic;
signal \N__49295\ : std_logic;
signal \N__49292\ : std_logic;
signal \N__49289\ : std_logic;
signal \N__49284\ : std_logic;
signal \N__49281\ : std_logic;
signal \N__49280\ : std_logic;
signal \N__49277\ : std_logic;
signal \N__49274\ : std_logic;
signal \N__49271\ : std_logic;
signal \N__49266\ : std_logic;
signal \N__49263\ : std_logic;
signal \N__49260\ : std_logic;
signal \N__49257\ : std_logic;
signal \N__49254\ : std_logic;
signal \N__49251\ : std_logic;
signal \N__49250\ : std_logic;
signal \N__49249\ : std_logic;
signal \N__49248\ : std_logic;
signal \N__49247\ : std_logic;
signal \N__49246\ : std_logic;
signal \N__49245\ : std_logic;
signal \N__49244\ : std_logic;
signal \N__49243\ : std_logic;
signal \N__49242\ : std_logic;
signal \N__49241\ : std_logic;
signal \N__49240\ : std_logic;
signal \N__49239\ : std_logic;
signal \N__49238\ : std_logic;
signal \N__49237\ : std_logic;
signal \N__49236\ : std_logic;
signal \N__49235\ : std_logic;
signal \N__49234\ : std_logic;
signal \N__49233\ : std_logic;
signal \N__49232\ : std_logic;
signal \N__49231\ : std_logic;
signal \N__49230\ : std_logic;
signal \N__49229\ : std_logic;
signal \N__49228\ : std_logic;
signal \N__49227\ : std_logic;
signal \N__49226\ : std_logic;
signal \N__49225\ : std_logic;
signal \N__49224\ : std_logic;
signal \N__49223\ : std_logic;
signal \N__49222\ : std_logic;
signal \N__49221\ : std_logic;
signal \N__49220\ : std_logic;
signal \N__49219\ : std_logic;
signal \N__49218\ : std_logic;
signal \N__49217\ : std_logic;
signal \N__49216\ : std_logic;
signal \N__49215\ : std_logic;
signal \N__49214\ : std_logic;
signal \N__49213\ : std_logic;
signal \N__49212\ : std_logic;
signal \N__49211\ : std_logic;
signal \N__49210\ : std_logic;
signal \N__49209\ : std_logic;
signal \N__49208\ : std_logic;
signal \N__49207\ : std_logic;
signal \N__49206\ : std_logic;
signal \N__49205\ : std_logic;
signal \N__49204\ : std_logic;
signal \N__49203\ : std_logic;
signal \N__49202\ : std_logic;
signal \N__49201\ : std_logic;
signal \N__49200\ : std_logic;
signal \N__49199\ : std_logic;
signal \N__49198\ : std_logic;
signal \N__49197\ : std_logic;
signal \N__49196\ : std_logic;
signal \N__49195\ : std_logic;
signal \N__49194\ : std_logic;
signal \N__49193\ : std_logic;
signal \N__49192\ : std_logic;
signal \N__49191\ : std_logic;
signal \N__49190\ : std_logic;
signal \N__49189\ : std_logic;
signal \N__49188\ : std_logic;
signal \N__49187\ : std_logic;
signal \N__49186\ : std_logic;
signal \N__49185\ : std_logic;
signal \N__49184\ : std_logic;
signal \N__49183\ : std_logic;
signal \N__49182\ : std_logic;
signal \N__49181\ : std_logic;
signal \N__49180\ : std_logic;
signal \N__49179\ : std_logic;
signal \N__49178\ : std_logic;
signal \N__49177\ : std_logic;
signal \N__49176\ : std_logic;
signal \N__49175\ : std_logic;
signal \N__49174\ : std_logic;
signal \N__49173\ : std_logic;
signal \N__49172\ : std_logic;
signal \N__49171\ : std_logic;
signal \N__49170\ : std_logic;
signal \N__49169\ : std_logic;
signal \N__49168\ : std_logic;
signal \N__49167\ : std_logic;
signal \N__49166\ : std_logic;
signal \N__49165\ : std_logic;
signal \N__49164\ : std_logic;
signal \N__49163\ : std_logic;
signal \N__49162\ : std_logic;
signal \N__49161\ : std_logic;
signal \N__49160\ : std_logic;
signal \N__49159\ : std_logic;
signal \N__49158\ : std_logic;
signal \N__49157\ : std_logic;
signal \N__49156\ : std_logic;
signal \N__49155\ : std_logic;
signal \N__49154\ : std_logic;
signal \N__49153\ : std_logic;
signal \N__49152\ : std_logic;
signal \N__49151\ : std_logic;
signal \N__49150\ : std_logic;
signal \N__49149\ : std_logic;
signal \N__49148\ : std_logic;
signal \N__49147\ : std_logic;
signal \N__49146\ : std_logic;
signal \N__49145\ : std_logic;
signal \N__49144\ : std_logic;
signal \N__49143\ : std_logic;
signal \N__49142\ : std_logic;
signal \N__49141\ : std_logic;
signal \N__49140\ : std_logic;
signal \N__49139\ : std_logic;
signal \N__49138\ : std_logic;
signal \N__49137\ : std_logic;
signal \N__49136\ : std_logic;
signal \N__49135\ : std_logic;
signal \N__49134\ : std_logic;
signal \N__49133\ : std_logic;
signal \N__49132\ : std_logic;
signal \N__49131\ : std_logic;
signal \N__49130\ : std_logic;
signal \N__49129\ : std_logic;
signal \N__49128\ : std_logic;
signal \N__49127\ : std_logic;
signal \N__49126\ : std_logic;
signal \N__49125\ : std_logic;
signal \N__49124\ : std_logic;
signal \N__49123\ : std_logic;
signal \N__49122\ : std_logic;
signal \N__49121\ : std_logic;
signal \N__49120\ : std_logic;
signal \N__49119\ : std_logic;
signal \N__49118\ : std_logic;
signal \N__49117\ : std_logic;
signal \N__49116\ : std_logic;
signal \N__49115\ : std_logic;
signal \N__49114\ : std_logic;
signal \N__49113\ : std_logic;
signal \N__49112\ : std_logic;
signal \N__49111\ : std_logic;
signal \N__49110\ : std_logic;
signal \N__48825\ : std_logic;
signal \N__48822\ : std_logic;
signal \N__48821\ : std_logic;
signal \N__48820\ : std_logic;
signal \N__48819\ : std_logic;
signal \N__48816\ : std_logic;
signal \N__48815\ : std_logic;
signal \N__48814\ : std_logic;
signal \N__48813\ : std_logic;
signal \N__48812\ : std_logic;
signal \N__48811\ : std_logic;
signal \N__48808\ : std_logic;
signal \N__48807\ : std_logic;
signal \N__48806\ : std_logic;
signal \N__48805\ : std_logic;
signal \N__48804\ : std_logic;
signal \N__48803\ : std_logic;
signal \N__48802\ : std_logic;
signal \N__48801\ : std_logic;
signal \N__48798\ : std_logic;
signal \N__48795\ : std_logic;
signal \N__48792\ : std_logic;
signal \N__48783\ : std_logic;
signal \N__48780\ : std_logic;
signal \N__48777\ : std_logic;
signal \N__48770\ : std_logic;
signal \N__48767\ : std_logic;
signal \N__48764\ : std_logic;
signal \N__48763\ : std_logic;
signal \N__48762\ : std_logic;
signal \N__48761\ : std_logic;
signal \N__48760\ : std_logic;
signal \N__48759\ : std_logic;
signal \N__48758\ : std_logic;
signal \N__48757\ : std_logic;
signal \N__48756\ : std_logic;
signal \N__48755\ : std_logic;
signal \N__48754\ : std_logic;
signal \N__48753\ : std_logic;
signal \N__48752\ : std_logic;
signal \N__48751\ : std_logic;
signal \N__48750\ : std_logic;
signal \N__48749\ : std_logic;
signal \N__48748\ : std_logic;
signal \N__48747\ : std_logic;
signal \N__48746\ : std_logic;
signal \N__48745\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48736\ : std_logic;
signal \N__48733\ : std_logic;
signal \N__48730\ : std_logic;
signal \N__48727\ : std_logic;
signal \N__48722\ : std_logic;
signal \N__48717\ : std_logic;
signal \N__48714\ : std_logic;
signal \N__48705\ : std_logic;
signal \N__48696\ : std_logic;
signal \N__48689\ : std_logic;
signal \N__48680\ : std_logic;
signal \N__48671\ : std_logic;
signal \N__48670\ : std_logic;
signal \N__48669\ : std_logic;
signal \N__48668\ : std_logic;
signal \N__48667\ : std_logic;
signal \N__48666\ : std_logic;
signal \N__48663\ : std_logic;
signal \N__48660\ : std_logic;
signal \N__48655\ : std_logic;
signal \N__48652\ : std_logic;
signal \N__48645\ : std_logic;
signal \N__48638\ : std_logic;
signal \N__48631\ : std_logic;
signal \N__48622\ : std_logic;
signal \N__48619\ : std_logic;
signal \N__48616\ : std_logic;
signal \N__48611\ : std_logic;
signal \N__48602\ : std_logic;
signal \N__48591\ : std_logic;
signal \N__48590\ : std_logic;
signal \N__48589\ : std_logic;
signal \N__48588\ : std_logic;
signal \N__48587\ : std_logic;
signal \N__48586\ : std_logic;
signal \N__48585\ : std_logic;
signal \N__48584\ : std_logic;
signal \N__48583\ : std_logic;
signal \N__48580\ : std_logic;
signal \N__48577\ : std_logic;
signal \N__48574\ : std_logic;
signal \N__48571\ : std_logic;
signal \N__48568\ : std_logic;
signal \N__48565\ : std_logic;
signal \N__48562\ : std_logic;
signal \N__48559\ : std_logic;
signal \N__48556\ : std_logic;
signal \N__48553\ : std_logic;
signal \N__48550\ : std_logic;
signal \N__48547\ : std_logic;
signal \N__48546\ : std_logic;
signal \N__48545\ : std_logic;
signal \N__48544\ : std_logic;
signal \N__48543\ : std_logic;
signal \N__48542\ : std_logic;
signal \N__48541\ : std_logic;
signal \N__48540\ : std_logic;
signal \N__48539\ : std_logic;
signal \N__48538\ : std_logic;
signal \N__48537\ : std_logic;
signal \N__48536\ : std_logic;
signal \N__48535\ : std_logic;
signal \N__48534\ : std_logic;
signal \N__48533\ : std_logic;
signal \N__48532\ : std_logic;
signal \N__48531\ : std_logic;
signal \N__48530\ : std_logic;
signal \N__48529\ : std_logic;
signal \N__48528\ : std_logic;
signal \N__48527\ : std_logic;
signal \N__48526\ : std_logic;
signal \N__48525\ : std_logic;
signal \N__48524\ : std_logic;
signal \N__48523\ : std_logic;
signal \N__48522\ : std_logic;
signal \N__48521\ : std_logic;
signal \N__48520\ : std_logic;
signal \N__48519\ : std_logic;
signal \N__48518\ : std_logic;
signal \N__48517\ : std_logic;
signal \N__48516\ : std_logic;
signal \N__48515\ : std_logic;
signal \N__48514\ : std_logic;
signal \N__48513\ : std_logic;
signal \N__48512\ : std_logic;
signal \N__48511\ : std_logic;
signal \N__48510\ : std_logic;
signal \N__48509\ : std_logic;
signal \N__48508\ : std_logic;
signal \N__48507\ : std_logic;
signal \N__48506\ : std_logic;
signal \N__48505\ : std_logic;
signal \N__48504\ : std_logic;
signal \N__48501\ : std_logic;
signal \N__48500\ : std_logic;
signal \N__48499\ : std_logic;
signal \N__48498\ : std_logic;
signal \N__48497\ : std_logic;
signal \N__48496\ : std_logic;
signal \N__48495\ : std_logic;
signal \N__48494\ : std_logic;
signal \N__48493\ : std_logic;
signal \N__48492\ : std_logic;
signal \N__48489\ : std_logic;
signal \N__48488\ : std_logic;
signal \N__48487\ : std_logic;
signal \N__48486\ : std_logic;
signal \N__48485\ : std_logic;
signal \N__48484\ : std_logic;
signal \N__48483\ : std_logic;
signal \N__48482\ : std_logic;
signal \N__48481\ : std_logic;
signal \N__48480\ : std_logic;
signal \N__48479\ : std_logic;
signal \N__48478\ : std_logic;
signal \N__48477\ : std_logic;
signal \N__48476\ : std_logic;
signal \N__48475\ : std_logic;
signal \N__48474\ : std_logic;
signal \N__48473\ : std_logic;
signal \N__48472\ : std_logic;
signal \N__48471\ : std_logic;
signal \N__48470\ : std_logic;
signal \N__48469\ : std_logic;
signal \N__48468\ : std_logic;
signal \N__48467\ : std_logic;
signal \N__48466\ : std_logic;
signal \N__48465\ : std_logic;
signal \N__48464\ : std_logic;
signal \N__48463\ : std_logic;
signal \N__48462\ : std_logic;
signal \N__48461\ : std_logic;
signal \N__48460\ : std_logic;
signal \N__48459\ : std_logic;
signal \N__48458\ : std_logic;
signal \N__48457\ : std_logic;
signal \N__48456\ : std_logic;
signal \N__48455\ : std_logic;
signal \N__48454\ : std_logic;
signal \N__48453\ : std_logic;
signal \N__48450\ : std_logic;
signal \N__48449\ : std_logic;
signal \N__48448\ : std_logic;
signal \N__48447\ : std_logic;
signal \N__48446\ : std_logic;
signal \N__48445\ : std_logic;
signal \N__48444\ : std_logic;
signal \N__48443\ : std_logic;
signal \N__48442\ : std_logic;
signal \N__48441\ : std_logic;
signal \N__48438\ : std_logic;
signal \N__48437\ : std_logic;
signal \N__48436\ : std_logic;
signal \N__48435\ : std_logic;
signal \N__48434\ : std_logic;
signal \N__48433\ : std_logic;
signal \N__48432\ : std_logic;
signal \N__48431\ : std_logic;
signal \N__48430\ : std_logic;
signal \N__48429\ : std_logic;
signal \N__48428\ : std_logic;
signal \N__48427\ : std_logic;
signal \N__48426\ : std_logic;
signal \N__48423\ : std_logic;
signal \N__48422\ : std_logic;
signal \N__48421\ : std_logic;
signal \N__48420\ : std_logic;
signal \N__48419\ : std_logic;
signal \N__48418\ : std_logic;
signal \N__48417\ : std_logic;
signal \N__48416\ : std_logic;
signal \N__48415\ : std_logic;
signal \N__48414\ : std_logic;
signal \N__48413\ : std_logic;
signal \N__48412\ : std_logic;
signal \N__48409\ : std_logic;
signal \N__48408\ : std_logic;
signal \N__48407\ : std_logic;
signal \N__48406\ : std_logic;
signal \N__48405\ : std_logic;
signal \N__48404\ : std_logic;
signal \N__48403\ : std_logic;
signal \N__48402\ : std_logic;
signal \N__48401\ : std_logic;
signal \N__48400\ : std_logic;
signal \N__48399\ : std_logic;
signal \N__48398\ : std_logic;
signal \N__48397\ : std_logic;
signal \N__48396\ : std_logic;
signal \N__48395\ : std_logic;
signal \N__48394\ : std_logic;
signal \N__48393\ : std_logic;
signal \N__48392\ : std_logic;
signal \N__48391\ : std_logic;
signal \N__48096\ : std_logic;
signal \N__48093\ : std_logic;
signal \N__48090\ : std_logic;
signal \N__48089\ : std_logic;
signal \N__48088\ : std_logic;
signal \N__48087\ : std_logic;
signal \N__48086\ : std_logic;
signal \N__48085\ : std_logic;
signal \N__48084\ : std_logic;
signal \N__48083\ : std_logic;
signal \N__48082\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48080\ : std_logic;
signal \N__48079\ : std_logic;
signal \N__48078\ : std_logic;
signal \N__48077\ : std_logic;
signal \N__48076\ : std_logic;
signal \N__48075\ : std_logic;
signal \N__48074\ : std_logic;
signal \N__48073\ : std_logic;
signal \N__48072\ : std_logic;
signal \N__48071\ : std_logic;
signal \N__48070\ : std_logic;
signal \N__48069\ : std_logic;
signal \N__48068\ : std_logic;
signal \N__48067\ : std_logic;
signal \N__48066\ : std_logic;
signal \N__48065\ : std_logic;
signal \N__48064\ : std_logic;
signal \N__48063\ : std_logic;
signal \N__48062\ : std_logic;
signal \N__48061\ : std_logic;
signal \N__48052\ : std_logic;
signal \N__48043\ : std_logic;
signal \N__48038\ : std_logic;
signal \N__48029\ : std_logic;
signal \N__48020\ : std_logic;
signal \N__48011\ : std_logic;
signal \N__48002\ : std_logic;
signal \N__47993\ : std_logic;
signal \N__47990\ : std_logic;
signal \N__47987\ : std_logic;
signal \N__47974\ : std_logic;
signal \N__47971\ : std_logic;
signal \N__47966\ : std_logic;
signal \N__47961\ : std_logic;
signal \N__47958\ : std_logic;
signal \N__47957\ : std_logic;
signal \N__47954\ : std_logic;
signal \N__47951\ : std_logic;
signal \N__47946\ : std_logic;
signal \N__47945\ : std_logic;
signal \N__47944\ : std_logic;
signal \N__47941\ : std_logic;
signal \N__47938\ : std_logic;
signal \N__47935\ : std_logic;
signal \N__47934\ : std_logic;
signal \N__47929\ : std_logic;
signal \N__47926\ : std_logic;
signal \N__47923\ : std_logic;
signal \N__47920\ : std_logic;
signal \N__47915\ : std_logic;
signal \N__47910\ : std_logic;
signal \N__47907\ : std_logic;
signal \N__47904\ : std_logic;
signal \N__47901\ : std_logic;
signal \N__47898\ : std_logic;
signal \N__47897\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47891\ : std_logic;
signal \N__47886\ : std_logic;
signal \N__47885\ : std_logic;
signal \N__47882\ : std_logic;
signal \N__47881\ : std_logic;
signal \N__47878\ : std_logic;
signal \N__47875\ : std_logic;
signal \N__47872\ : std_logic;
signal \N__47871\ : std_logic;
signal \N__47868\ : std_logic;
signal \N__47863\ : std_logic;
signal \N__47860\ : std_logic;
signal \N__47857\ : std_logic;
signal \N__47854\ : std_logic;
signal \N__47847\ : std_logic;
signal \N__47846\ : std_logic;
signal \N__47843\ : std_logic;
signal \N__47842\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47838\ : std_logic;
signal \N__47835\ : std_logic;
signal \N__47832\ : std_logic;
signal \N__47829\ : std_logic;
signal \N__47828\ : std_logic;
signal \N__47827\ : std_logic;
signal \N__47826\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47822\ : std_logic;
signal \N__47819\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47807\ : std_logic;
signal \N__47804\ : std_logic;
signal \N__47801\ : std_logic;
signal \N__47796\ : std_logic;
signal \N__47787\ : std_logic;
signal \N__47784\ : std_logic;
signal \N__47783\ : std_logic;
signal \N__47782\ : std_logic;
signal \N__47779\ : std_logic;
signal \N__47776\ : std_logic;
signal \N__47773\ : std_logic;
signal \N__47770\ : std_logic;
signal \N__47767\ : std_logic;
signal \N__47766\ : std_logic;
signal \N__47763\ : std_logic;
signal \N__47760\ : std_logic;
signal \N__47757\ : std_logic;
signal \N__47754\ : std_logic;
signal \N__47751\ : std_logic;
signal \N__47742\ : std_logic;
signal \N__47739\ : std_logic;
signal \N__47736\ : std_logic;
signal \N__47735\ : std_logic;
signal \N__47732\ : std_logic;
signal \N__47729\ : std_logic;
signal \N__47728\ : std_logic;
signal \N__47723\ : std_logic;
signal \N__47720\ : std_logic;
signal \N__47715\ : std_logic;
signal \N__47712\ : std_logic;
signal \N__47709\ : std_logic;
signal \N__47706\ : std_logic;
signal \N__47703\ : std_logic;
signal \N__47702\ : std_logic;
signal \N__47701\ : std_logic;
signal \N__47700\ : std_logic;
signal \N__47699\ : std_logic;
signal \N__47698\ : std_logic;
signal \N__47695\ : std_logic;
signal \N__47692\ : std_logic;
signal \N__47691\ : std_logic;
signal \N__47690\ : std_logic;
signal \N__47687\ : std_logic;
signal \N__47684\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47677\ : std_logic;
signal \N__47672\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47668\ : std_logic;
signal \N__47663\ : std_logic;
signal \N__47662\ : std_logic;
signal \N__47659\ : std_logic;
signal \N__47656\ : std_logic;
signal \N__47653\ : std_logic;
signal \N__47650\ : std_logic;
signal \N__47645\ : std_logic;
signal \N__47644\ : std_logic;
signal \N__47641\ : std_logic;
signal \N__47638\ : std_logic;
signal \N__47635\ : std_logic;
signal \N__47634\ : std_logic;
signal \N__47633\ : std_logic;
signal \N__47632\ : std_logic;
signal \N__47631\ : std_logic;
signal \N__47630\ : std_logic;
signal \N__47627\ : std_logic;
signal \N__47626\ : std_logic;
signal \N__47619\ : std_logic;
signal \N__47616\ : std_logic;
signal \N__47615\ : std_logic;
signal \N__47612\ : std_logic;
signal \N__47611\ : std_logic;
signal \N__47610\ : std_logic;
signal \N__47605\ : std_logic;
signal \N__47602\ : std_logic;
signal \N__47597\ : std_logic;
signal \N__47590\ : std_logic;
signal \N__47587\ : std_logic;
signal \N__47584\ : std_logic;
signal \N__47579\ : std_logic;
signal \N__47576\ : std_logic;
signal \N__47569\ : std_logic;
signal \N__47566\ : std_logic;
signal \N__47559\ : std_logic;
signal \N__47544\ : std_logic;
signal \N__47541\ : std_logic;
signal \N__47538\ : std_logic;
signal \N__47537\ : std_logic;
signal \N__47534\ : std_logic;
signal \N__47531\ : std_logic;
signal \N__47528\ : std_logic;
signal \N__47527\ : std_logic;
signal \N__47524\ : std_logic;
signal \N__47521\ : std_logic;
signal \N__47520\ : std_logic;
signal \N__47517\ : std_logic;
signal \N__47512\ : std_logic;
signal \N__47509\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47499\ : std_logic;
signal \N__47496\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47490\ : std_logic;
signal \N__47487\ : std_logic;
signal \N__47484\ : std_logic;
signal \N__47481\ : std_logic;
signal \N__47478\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47476\ : std_logic;
signal \N__47473\ : std_logic;
signal \N__47470\ : std_logic;
signal \N__47467\ : std_logic;
signal \N__47460\ : std_logic;
signal \N__47457\ : std_logic;
signal \N__47454\ : std_logic;
signal \N__47453\ : std_logic;
signal \N__47452\ : std_logic;
signal \N__47449\ : std_logic;
signal \N__47446\ : std_logic;
signal \N__47443\ : std_logic;
signal \N__47436\ : std_logic;
signal \N__47433\ : std_logic;
signal \N__47430\ : std_logic;
signal \N__47429\ : std_logic;
signal \N__47428\ : std_logic;
signal \N__47425\ : std_logic;
signal \N__47422\ : std_logic;
signal \N__47419\ : std_logic;
signal \N__47412\ : std_logic;
signal \N__47409\ : std_logic;
signal \N__47406\ : std_logic;
signal \N__47405\ : std_logic;
signal \N__47404\ : std_logic;
signal \N__47401\ : std_logic;
signal \N__47398\ : std_logic;
signal \N__47395\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47385\ : std_logic;
signal \N__47382\ : std_logic;
signal \N__47381\ : std_logic;
signal \N__47380\ : std_logic;
signal \N__47377\ : std_logic;
signal \N__47374\ : std_logic;
signal \N__47371\ : std_logic;
signal \N__47364\ : std_logic;
signal \N__47361\ : std_logic;
signal \N__47358\ : std_logic;
signal \N__47357\ : std_logic;
signal \N__47356\ : std_logic;
signal \N__47353\ : std_logic;
signal \N__47350\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47340\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47334\ : std_logic;
signal \N__47333\ : std_logic;
signal \N__47332\ : std_logic;
signal \N__47329\ : std_logic;
signal \N__47326\ : std_logic;
signal \N__47323\ : std_logic;
signal \N__47316\ : std_logic;
signal \N__47313\ : std_logic;
signal \N__47312\ : std_logic;
signal \N__47309\ : std_logic;
signal \N__47306\ : std_logic;
signal \N__47301\ : std_logic;
signal \N__47298\ : std_logic;
signal \N__47295\ : std_logic;
signal \N__47294\ : std_logic;
signal \N__47293\ : std_logic;
signal \N__47290\ : std_logic;
signal \N__47287\ : std_logic;
signal \N__47284\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47274\ : std_logic;
signal \N__47271\ : std_logic;
signal \N__47270\ : std_logic;
signal \N__47269\ : std_logic;
signal \N__47266\ : std_logic;
signal \N__47263\ : std_logic;
signal \N__47260\ : std_logic;
signal \N__47253\ : std_logic;
signal \N__47250\ : std_logic;
signal \N__47247\ : std_logic;
signal \N__47246\ : std_logic;
signal \N__47245\ : std_logic;
signal \N__47242\ : std_logic;
signal \N__47239\ : std_logic;
signal \N__47236\ : std_logic;
signal \N__47229\ : std_logic;
signal \N__47226\ : std_logic;
signal \N__47223\ : std_logic;
signal \N__47222\ : std_logic;
signal \N__47221\ : std_logic;
signal \N__47218\ : std_logic;
signal \N__47215\ : std_logic;
signal \N__47212\ : std_logic;
signal \N__47205\ : std_logic;
signal \N__47202\ : std_logic;
signal \N__47199\ : std_logic;
signal \N__47198\ : std_logic;
signal \N__47197\ : std_logic;
signal \N__47194\ : std_logic;
signal \N__47191\ : std_logic;
signal \N__47188\ : std_logic;
signal \N__47181\ : std_logic;
signal \N__47178\ : std_logic;
signal \N__47175\ : std_logic;
signal \N__47174\ : std_logic;
signal \N__47173\ : std_logic;
signal \N__47170\ : std_logic;
signal \N__47167\ : std_logic;
signal \N__47164\ : std_logic;
signal \N__47157\ : std_logic;
signal \N__47154\ : std_logic;
signal \N__47151\ : std_logic;
signal \N__47150\ : std_logic;
signal \N__47149\ : std_logic;
signal \N__47146\ : std_logic;
signal \N__47143\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47133\ : std_logic;
signal \N__47130\ : std_logic;
signal \N__47127\ : std_logic;
signal \N__47126\ : std_logic;
signal \N__47125\ : std_logic;
signal \N__47122\ : std_logic;
signal \N__47119\ : std_logic;
signal \N__47116\ : std_logic;
signal \N__47109\ : std_logic;
signal \N__47106\ : std_logic;
signal \N__47103\ : std_logic;
signal \N__47102\ : std_logic;
signal \N__47101\ : std_logic;
signal \N__47098\ : std_logic;
signal \N__47095\ : std_logic;
signal \N__47092\ : std_logic;
signal \N__47085\ : std_logic;
signal \N__47082\ : std_logic;
signal \N__47079\ : std_logic;
signal \N__47078\ : std_logic;
signal \N__47077\ : std_logic;
signal \N__47074\ : std_logic;
signal \N__47071\ : std_logic;
signal \N__47068\ : std_logic;
signal \N__47061\ : std_logic;
signal \N__47058\ : std_logic;
signal \N__47055\ : std_logic;
signal \N__47054\ : std_logic;
signal \N__47053\ : std_logic;
signal \N__47050\ : std_logic;
signal \N__47047\ : std_logic;
signal \N__47044\ : std_logic;
signal \N__47037\ : std_logic;
signal \N__47034\ : std_logic;
signal \N__47031\ : std_logic;
signal \N__47030\ : std_logic;
signal \N__47029\ : std_logic;
signal \N__47026\ : std_logic;
signal \N__47023\ : std_logic;
signal \N__47020\ : std_logic;
signal \N__47013\ : std_logic;
signal \N__47010\ : std_logic;
signal \N__47007\ : std_logic;
signal \N__47006\ : std_logic;
signal \N__47005\ : std_logic;
signal \N__47002\ : std_logic;
signal \N__46999\ : std_logic;
signal \N__46996\ : std_logic;
signal \N__46989\ : std_logic;
signal \N__46986\ : std_logic;
signal \N__46983\ : std_logic;
signal \N__46982\ : std_logic;
signal \N__46981\ : std_logic;
signal \N__46978\ : std_logic;
signal \N__46975\ : std_logic;
signal \N__46972\ : std_logic;
signal \N__46965\ : std_logic;
signal \N__46962\ : std_logic;
signal \N__46959\ : std_logic;
signal \N__46958\ : std_logic;
signal \N__46957\ : std_logic;
signal \N__46954\ : std_logic;
signal \N__46951\ : std_logic;
signal \N__46948\ : std_logic;
signal \N__46941\ : std_logic;
signal \N__46938\ : std_logic;
signal \N__46935\ : std_logic;
signal \N__46934\ : std_logic;
signal \N__46933\ : std_logic;
signal \N__46930\ : std_logic;
signal \N__46927\ : std_logic;
signal \N__46924\ : std_logic;
signal \N__46917\ : std_logic;
signal \N__46914\ : std_logic;
signal \N__46911\ : std_logic;
signal \N__46910\ : std_logic;
signal \N__46909\ : std_logic;
signal \N__46906\ : std_logic;
signal \N__46903\ : std_logic;
signal \N__46900\ : std_logic;
signal \N__46893\ : std_logic;
signal \N__46890\ : std_logic;
signal \N__46887\ : std_logic;
signal \N__46886\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46882\ : std_logic;
signal \N__46879\ : std_logic;
signal \N__46878\ : std_logic;
signal \N__46875\ : std_logic;
signal \N__46874\ : std_logic;
signal \N__46869\ : std_logic;
signal \N__46868\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46864\ : std_logic;
signal \N__46861\ : std_logic;
signal \N__46860\ : std_logic;
signal \N__46857\ : std_logic;
signal \N__46854\ : std_logic;
signal \N__46851\ : std_logic;
signal \N__46848\ : std_logic;
signal \N__46843\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46827\ : std_logic;
signal \N__46824\ : std_logic;
signal \N__46823\ : std_logic;
signal \N__46822\ : std_logic;
signal \N__46821\ : std_logic;
signal \N__46820\ : std_logic;
signal \N__46819\ : std_logic;
signal \N__46818\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46816\ : std_logic;
signal \N__46815\ : std_logic;
signal \N__46814\ : std_logic;
signal \N__46813\ : std_logic;
signal \N__46812\ : std_logic;
signal \N__46809\ : std_logic;
signal \N__46808\ : std_logic;
signal \N__46807\ : std_logic;
signal \N__46804\ : std_logic;
signal \N__46797\ : std_logic;
signal \N__46794\ : std_logic;
signal \N__46791\ : std_logic;
signal \N__46784\ : std_logic;
signal \N__46779\ : std_logic;
signal \N__46776\ : std_logic;
signal \N__46773\ : std_logic;
signal \N__46772\ : std_logic;
signal \N__46769\ : std_logic;
signal \N__46768\ : std_logic;
signal \N__46767\ : std_logic;
signal \N__46766\ : std_logic;
signal \N__46765\ : std_logic;
signal \N__46764\ : std_logic;
signal \N__46761\ : std_logic;
signal \N__46758\ : std_logic;
signal \N__46753\ : std_logic;
signal \N__46752\ : std_logic;
signal \N__46751\ : std_logic;
signal \N__46750\ : std_logic;
signal \N__46749\ : std_logic;
signal \N__46748\ : std_logic;
signal \N__46745\ : std_logic;
signal \N__46738\ : std_logic;
signal \N__46735\ : std_logic;
signal \N__46728\ : std_logic;
signal \N__46727\ : std_logic;
signal \N__46722\ : std_logic;
signal \N__46715\ : std_logic;
signal \N__46712\ : std_logic;
signal \N__46709\ : std_logic;
signal \N__46698\ : std_logic;
signal \N__46689\ : std_logic;
signal \N__46686\ : std_logic;
signal \N__46671\ : std_logic;
signal \N__46668\ : std_logic;
signal \N__46665\ : std_logic;
signal \N__46662\ : std_logic;
signal \N__46659\ : std_logic;
signal \N__46656\ : std_logic;
signal \N__46653\ : std_logic;
signal \N__46650\ : std_logic;
signal \N__46647\ : std_logic;
signal \N__46644\ : std_logic;
signal \N__46641\ : std_logic;
signal \N__46638\ : std_logic;
signal \N__46635\ : std_logic;
signal \N__46632\ : std_logic;
signal \N__46631\ : std_logic;
signal \N__46630\ : std_logic;
signal \N__46627\ : std_logic;
signal \N__46622\ : std_logic;
signal \N__46617\ : std_logic;
signal \N__46614\ : std_logic;
signal \N__46611\ : std_logic;
signal \N__46608\ : std_logic;
signal \N__46605\ : std_logic;
signal \N__46602\ : std_logic;
signal \N__46599\ : std_logic;
signal \N__46596\ : std_logic;
signal \N__46595\ : std_logic;
signal \N__46594\ : std_logic;
signal \N__46591\ : std_logic;
signal \N__46588\ : std_logic;
signal \N__46585\ : std_logic;
signal \N__46578\ : std_logic;
signal \N__46575\ : std_logic;
signal \N__46572\ : std_logic;
signal \N__46571\ : std_logic;
signal \N__46570\ : std_logic;
signal \N__46567\ : std_logic;
signal \N__46564\ : std_logic;
signal \N__46561\ : std_logic;
signal \N__46554\ : std_logic;
signal \N__46551\ : std_logic;
signal \N__46548\ : std_logic;
signal \N__46547\ : std_logic;
signal \N__46544\ : std_logic;
signal \N__46541\ : std_logic;
signal \N__46538\ : std_logic;
signal \N__46537\ : std_logic;
signal \N__46536\ : std_logic;
signal \N__46533\ : std_logic;
signal \N__46530\ : std_logic;
signal \N__46525\ : std_logic;
signal \N__46518\ : std_logic;
signal \N__46515\ : std_logic;
signal \N__46512\ : std_logic;
signal \N__46509\ : std_logic;
signal \N__46506\ : std_logic;
signal \N__46503\ : std_logic;
signal \N__46500\ : std_logic;
signal \N__46497\ : std_logic;
signal \N__46494\ : std_logic;
signal \N__46491\ : std_logic;
signal \N__46488\ : std_logic;
signal \N__46485\ : std_logic;
signal \N__46484\ : std_logic;
signal \N__46481\ : std_logic;
signal \N__46480\ : std_logic;
signal \N__46477\ : std_logic;
signal \N__46474\ : std_logic;
signal \N__46473\ : std_logic;
signal \N__46472\ : std_logic;
signal \N__46469\ : std_logic;
signal \N__46466\ : std_logic;
signal \N__46463\ : std_logic;
signal \N__46460\ : std_logic;
signal \N__46457\ : std_logic;
signal \N__46446\ : std_logic;
signal \N__46445\ : std_logic;
signal \N__46442\ : std_logic;
signal \N__46437\ : std_logic;
signal \N__46434\ : std_logic;
signal \N__46431\ : std_logic;
signal \N__46428\ : std_logic;
signal \N__46427\ : std_logic;
signal \N__46424\ : std_logic;
signal \N__46423\ : std_logic;
signal \N__46422\ : std_logic;
signal \N__46419\ : std_logic;
signal \N__46416\ : std_logic;
signal \N__46413\ : std_logic;
signal \N__46410\ : std_logic;
signal \N__46401\ : std_logic;
signal \N__46400\ : std_logic;
signal \N__46399\ : std_logic;
signal \N__46396\ : std_logic;
signal \N__46391\ : std_logic;
signal \N__46386\ : std_logic;
signal \N__46383\ : std_logic;
signal \N__46382\ : std_logic;
signal \N__46379\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46373\ : std_logic;
signal \N__46368\ : std_logic;
signal \N__46367\ : std_logic;
signal \N__46366\ : std_logic;
signal \N__46359\ : std_logic;
signal \N__46356\ : std_logic;
signal \N__46353\ : std_logic;
signal \N__46350\ : std_logic;
signal \N__46347\ : std_logic;
signal \N__46346\ : std_logic;
signal \N__46345\ : std_logic;
signal \N__46344\ : std_logic;
signal \N__46341\ : std_logic;
signal \N__46338\ : std_logic;
signal \N__46333\ : std_logic;
signal \N__46326\ : std_logic;
signal \N__46323\ : std_logic;
signal \N__46320\ : std_logic;
signal \N__46317\ : std_logic;
signal \N__46314\ : std_logic;
signal \N__46311\ : std_logic;
signal \N__46310\ : std_logic;
signal \N__46307\ : std_logic;
signal \N__46304\ : std_logic;
signal \N__46299\ : std_logic;
signal \N__46298\ : std_logic;
signal \N__46295\ : std_logic;
signal \N__46294\ : std_logic;
signal \N__46291\ : std_logic;
signal \N__46284\ : std_logic;
signal \N__46281\ : std_logic;
signal \N__46278\ : std_logic;
signal \N__46277\ : std_logic;
signal \N__46274\ : std_logic;
signal \N__46273\ : std_logic;
signal \N__46270\ : std_logic;
signal \N__46269\ : std_logic;
signal \N__46266\ : std_logic;
signal \N__46263\ : std_logic;
signal \N__46258\ : std_logic;
signal \N__46255\ : std_logic;
signal \N__46252\ : std_logic;
signal \N__46249\ : std_logic;
signal \N__46246\ : std_logic;
signal \N__46241\ : std_logic;
signal \N__46236\ : std_logic;
signal \N__46233\ : std_logic;
signal \N__46232\ : std_logic;
signal \N__46231\ : std_logic;
signal \N__46228\ : std_logic;
signal \N__46225\ : std_logic;
signal \N__46222\ : std_logic;
signal \N__46215\ : std_logic;
signal \N__46212\ : std_logic;
signal \N__46209\ : std_logic;
signal \N__46206\ : std_logic;
signal \N__46203\ : std_logic;
signal \N__46200\ : std_logic;
signal \N__46197\ : std_logic;
signal \N__46194\ : std_logic;
signal \N__46193\ : std_logic;
signal \N__46190\ : std_logic;
signal \N__46189\ : std_logic;
signal \N__46186\ : std_logic;
signal \N__46183\ : std_logic;
signal \N__46180\ : std_logic;
signal \N__46177\ : std_logic;
signal \N__46174\ : std_logic;
signal \N__46171\ : std_logic;
signal \N__46166\ : std_logic;
signal \N__46163\ : std_logic;
signal \N__46162\ : std_logic;
signal \N__46159\ : std_logic;
signal \N__46156\ : std_logic;
signal \N__46153\ : std_logic;
signal \N__46146\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46140\ : std_logic;
signal \N__46139\ : std_logic;
signal \N__46138\ : std_logic;
signal \N__46135\ : std_logic;
signal \N__46132\ : std_logic;
signal \N__46129\ : std_logic;
signal \N__46122\ : std_logic;
signal \N__46119\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46112\ : std_logic;
signal \N__46109\ : std_logic;
signal \N__46106\ : std_logic;
signal \N__46105\ : std_logic;
signal \N__46102\ : std_logic;
signal \N__46099\ : std_logic;
signal \N__46096\ : std_logic;
signal \N__46095\ : std_logic;
signal \N__46092\ : std_logic;
signal \N__46089\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46083\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46077\ : std_logic;
signal \N__46074\ : std_logic;
signal \N__46071\ : std_logic;
signal \N__46068\ : std_logic;
signal \N__46063\ : std_logic;
signal \N__46056\ : std_logic;
signal \N__46053\ : std_logic;
signal \N__46052\ : std_logic;
signal \N__46049\ : std_logic;
signal \N__46046\ : std_logic;
signal \N__46045\ : std_logic;
signal \N__46042\ : std_logic;
signal \N__46039\ : std_logic;
signal \N__46036\ : std_logic;
signal \N__46029\ : std_logic;
signal \N__46026\ : std_logic;
signal \N__46023\ : std_logic;
signal \N__46020\ : std_logic;
signal \N__46017\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46013\ : std_logic;
signal \N__46012\ : std_logic;
signal \N__46011\ : std_logic;
signal \N__46010\ : std_logic;
signal \N__46009\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46007\ : std_logic;
signal \N__46006\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46004\ : std_logic;
signal \N__46003\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__46001\ : std_logic;
signal \N__46000\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45998\ : std_logic;
signal \N__45997\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45995\ : std_logic;
signal \N__45994\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45992\ : std_logic;
signal \N__45989\ : std_logic;
signal \N__45988\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45986\ : std_logic;
signal \N__45983\ : std_logic;
signal \N__45982\ : std_logic;
signal \N__45981\ : std_logic;
signal \N__45980\ : std_logic;
signal \N__45977\ : std_logic;
signal \N__45976\ : std_logic;
signal \N__45975\ : std_logic;
signal \N__45974\ : std_logic;
signal \N__45965\ : std_logic;
signal \N__45956\ : std_logic;
signal \N__45955\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45953\ : std_logic;
signal \N__45952\ : std_logic;
signal \N__45949\ : std_logic;
signal \N__45948\ : std_logic;
signal \N__45947\ : std_logic;
signal \N__45946\ : std_logic;
signal \N__45945\ : std_logic;
signal \N__45944\ : std_logic;
signal \N__45943\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45941\ : std_logic;
signal \N__45940\ : std_logic;
signal \N__45939\ : std_logic;
signal \N__45936\ : std_logic;
signal \N__45935\ : std_logic;
signal \N__45932\ : std_logic;
signal \N__45931\ : std_logic;
signal \N__45928\ : std_logic;
signal \N__45927\ : std_logic;
signal \N__45924\ : std_logic;
signal \N__45923\ : std_logic;
signal \N__45920\ : std_logic;
signal \N__45919\ : std_logic;
signal \N__45916\ : std_logic;
signal \N__45915\ : std_logic;
signal \N__45912\ : std_logic;
signal \N__45911\ : std_logic;
signal \N__45910\ : std_logic;
signal \N__45909\ : std_logic;
signal \N__45908\ : std_logic;
signal \N__45907\ : std_logic;
signal \N__45906\ : std_logic;
signal \N__45905\ : std_logic;
signal \N__45904\ : std_logic;
signal \N__45903\ : std_logic;
signal \N__45902\ : std_logic;
signal \N__45901\ : std_logic;
signal \N__45900\ : std_logic;
signal \N__45897\ : std_logic;
signal \N__45896\ : std_logic;
signal \N__45893\ : std_logic;
signal \N__45892\ : std_logic;
signal \N__45889\ : std_logic;
signal \N__45888\ : std_logic;
signal \N__45887\ : std_logic;
signal \N__45886\ : std_logic;
signal \N__45885\ : std_logic;
signal \N__45884\ : std_logic;
signal \N__45883\ : std_logic;
signal \N__45882\ : std_logic;
signal \N__45877\ : std_logic;
signal \N__45876\ : std_logic;
signal \N__45875\ : std_logic;
signal \N__45874\ : std_logic;
signal \N__45871\ : std_logic;
signal \N__45864\ : std_logic;
signal \N__45853\ : std_logic;
signal \N__45852\ : std_logic;
signal \N__45849\ : std_logic;
signal \N__45848\ : std_logic;
signal \N__45845\ : std_logic;
signal \N__45844\ : std_logic;
signal \N__45843\ : std_logic;
signal \N__45842\ : std_logic;
signal \N__45841\ : std_logic;
signal \N__45840\ : std_logic;
signal \N__45835\ : std_logic;
signal \N__45822\ : std_logic;
signal \N__45811\ : std_logic;
signal \N__45806\ : std_logic;
signal \N__45805\ : std_logic;
signal \N__45804\ : std_logic;
signal \N__45803\ : std_logic;
signal \N__45802\ : std_logic;
signal \N__45801\ : std_logic;
signal \N__45784\ : std_logic;
signal \N__45767\ : std_logic;
signal \N__45764\ : std_logic;
signal \N__45763\ : std_logic;
signal \N__45760\ : std_logic;
signal \N__45759\ : std_logic;
signal \N__45756\ : std_logic;
signal \N__45755\ : std_logic;
signal \N__45752\ : std_logic;
signal \N__45751\ : std_logic;
signal \N__45750\ : std_logic;
signal \N__45749\ : std_logic;
signal \N__45748\ : std_logic;
signal \N__45747\ : std_logic;
signal \N__45744\ : std_logic;
signal \N__45743\ : std_logic;
signal \N__45740\ : std_logic;
signal \N__45739\ : std_logic;
signal \N__45736\ : std_logic;
signal \N__45735\ : std_logic;
signal \N__45732\ : std_logic;
signal \N__45731\ : std_logic;
signal \N__45728\ : std_logic;
signal \N__45727\ : std_logic;
signal \N__45724\ : std_logic;
signal \N__45723\ : std_logic;
signal \N__45720\ : std_logic;
signal \N__45719\ : std_logic;
signal \N__45706\ : std_logic;
signal \N__45697\ : std_logic;
signal \N__45692\ : std_logic;
signal \N__45689\ : std_logic;
signal \N__45686\ : std_logic;
signal \N__45685\ : std_logic;
signal \N__45682\ : std_logic;
signal \N__45681\ : std_logic;
signal \N__45680\ : std_logic;
signal \N__45679\ : std_logic;
signal \N__45676\ : std_logic;
signal \N__45675\ : std_logic;
signal \N__45674\ : std_logic;
signal \N__45673\ : std_logic;
signal \N__45672\ : std_logic;
signal \N__45667\ : std_logic;
signal \N__45664\ : std_logic;
signal \N__45653\ : std_logic;
signal \N__45650\ : std_logic;
signal \N__45649\ : std_logic;
signal \N__45646\ : std_logic;
signal \N__45645\ : std_logic;
signal \N__45642\ : std_logic;
signal \N__45641\ : std_logic;
signal \N__45638\ : std_logic;
signal \N__45637\ : std_logic;
signal \N__45628\ : std_logic;
signal \N__45617\ : std_logic;
signal \N__45612\ : std_logic;
signal \N__45595\ : std_logic;
signal \N__45592\ : std_logic;
signal \N__45591\ : std_logic;
signal \N__45588\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45584\ : std_logic;
signal \N__45583\ : std_logic;
signal \N__45568\ : std_logic;
signal \N__45551\ : std_logic;
signal \N__45548\ : std_logic;
signal \N__45543\ : std_logic;
signal \N__45538\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45516\ : std_logic;
signal \N__45509\ : std_logic;
signal \N__45492\ : std_logic;
signal \N__45483\ : std_logic;
signal \N__45470\ : std_logic;
signal \N__45463\ : std_logic;
signal \N__45444\ : std_logic;
signal \N__45443\ : std_logic;
signal \N__45442\ : std_logic;
signal \N__45441\ : std_logic;
signal \N__45440\ : std_logic;
signal \N__45439\ : std_logic;
signal \N__45438\ : std_logic;
signal \N__45437\ : std_logic;
signal \N__45436\ : std_logic;
signal \N__45435\ : std_logic;
signal \N__45434\ : std_logic;
signal \N__45433\ : std_logic;
signal \N__45432\ : std_logic;
signal \N__45431\ : std_logic;
signal \N__45430\ : std_logic;
signal \N__45429\ : std_logic;
signal \N__45428\ : std_logic;
signal \N__45427\ : std_logic;
signal \N__45426\ : std_logic;
signal \N__45425\ : std_logic;
signal \N__45424\ : std_logic;
signal \N__45423\ : std_logic;
signal \N__45422\ : std_logic;
signal \N__45421\ : std_logic;
signal \N__45420\ : std_logic;
signal \N__45419\ : std_logic;
signal \N__45418\ : std_logic;
signal \N__45417\ : std_logic;
signal \N__45416\ : std_logic;
signal \N__45415\ : std_logic;
signal \N__45414\ : std_logic;
signal \N__45413\ : std_logic;
signal \N__45412\ : std_logic;
signal \N__45411\ : std_logic;
signal \N__45410\ : std_logic;
signal \N__45409\ : std_logic;
signal \N__45408\ : std_logic;
signal \N__45407\ : std_logic;
signal \N__45406\ : std_logic;
signal \N__45405\ : std_logic;
signal \N__45404\ : std_logic;
signal \N__45403\ : std_logic;
signal \N__45400\ : std_logic;
signal \N__45399\ : std_logic;
signal \N__45398\ : std_logic;
signal \N__45397\ : std_logic;
signal \N__45396\ : std_logic;
signal \N__45395\ : std_logic;
signal \N__45394\ : std_logic;
signal \N__45393\ : std_logic;
signal \N__45392\ : std_logic;
signal \N__45389\ : std_logic;
signal \N__45378\ : std_logic;
signal \N__45365\ : std_logic;
signal \N__45364\ : std_logic;
signal \N__45355\ : std_logic;
signal \N__45346\ : std_logic;
signal \N__45345\ : std_logic;
signal \N__45344\ : std_logic;
signal \N__45343\ : std_logic;
signal \N__45342\ : std_logic;
signal \N__45341\ : std_logic;
signal \N__45340\ : std_logic;
signal \N__45339\ : std_logic;
signal \N__45338\ : std_logic;
signal \N__45333\ : std_logic;
signal \N__45324\ : std_logic;
signal \N__45313\ : std_logic;
signal \N__45306\ : std_logic;
signal \N__45303\ : std_logic;
signal \N__45302\ : std_logic;
signal \N__45301\ : std_logic;
signal \N__45300\ : std_logic;
signal \N__45299\ : std_logic;
signal \N__45298\ : std_logic;
signal \N__45297\ : std_logic;
signal \N__45286\ : std_logic;
signal \N__45283\ : std_logic;
signal \N__45268\ : std_logic;
signal \N__45267\ : std_logic;
signal \N__45266\ : std_logic;
signal \N__45263\ : std_logic;
signal \N__45260\ : std_logic;
signal \N__45257\ : std_logic;
signal \N__45252\ : std_logic;
signal \N__45251\ : std_logic;
signal \N__45250\ : std_logic;
signal \N__45249\ : std_logic;
signal \N__45246\ : std_logic;
signal \N__45245\ : std_logic;
signal \N__45242\ : std_logic;
signal \N__45239\ : std_logic;
signal \N__45236\ : std_logic;
signal \N__45221\ : std_logic;
signal \N__45216\ : std_logic;
signal \N__45213\ : std_logic;
signal \N__45208\ : std_logic;
signal \N__45195\ : std_logic;
signal \N__45192\ : std_logic;
signal \N__45187\ : std_logic;
signal \N__45182\ : std_logic;
signal \N__45173\ : std_logic;
signal \N__45162\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45156\ : std_logic;
signal \N__45145\ : std_logic;
signal \N__45126\ : std_logic;
signal \N__45123\ : std_logic;
signal \N__45122\ : std_logic;
signal \N__45119\ : std_logic;
signal \N__45116\ : std_logic;
signal \N__45115\ : std_logic;
signal \N__45112\ : std_logic;
signal \N__45107\ : std_logic;
signal \N__45102\ : std_logic;
signal \N__45101\ : std_logic;
signal \N__45096\ : std_logic;
signal \N__45095\ : std_logic;
signal \N__45094\ : std_logic;
signal \N__45091\ : std_logic;
signal \N__45086\ : std_logic;
signal \N__45083\ : std_logic;
signal \N__45080\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45072\ : std_logic;
signal \N__45069\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45063\ : std_logic;
signal \N__45060\ : std_logic;
signal \N__45057\ : std_logic;
signal \N__45054\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45048\ : std_logic;
signal \N__45045\ : std_logic;
signal \N__45042\ : std_logic;
signal \N__45039\ : std_logic;
signal \N__45036\ : std_logic;
signal \N__45033\ : std_logic;
signal \N__45032\ : std_logic;
signal \N__45029\ : std_logic;
signal \N__45026\ : std_logic;
signal \N__45021\ : std_logic;
signal \N__45018\ : std_logic;
signal \N__45015\ : std_logic;
signal \N__45012\ : std_logic;
signal \N__45009\ : std_logic;
signal \N__45006\ : std_logic;
signal \N__45003\ : std_logic;
signal \N__45002\ : std_logic;
signal \N__44999\ : std_logic;
signal \N__44998\ : std_logic;
signal \N__44995\ : std_logic;
signal \N__44994\ : std_logic;
signal \N__44991\ : std_logic;
signal \N__44988\ : std_logic;
signal \N__44985\ : std_logic;
signal \N__44982\ : std_logic;
signal \N__44977\ : std_logic;
signal \N__44974\ : std_logic;
signal \N__44969\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44961\ : std_logic;
signal \N__44958\ : std_logic;
signal \N__44957\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44950\ : std_logic;
signal \N__44947\ : std_logic;
signal \N__44940\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44928\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44924\ : std_logic;
signal \N__44921\ : std_logic;
signal \N__44918\ : std_logic;
signal \N__44917\ : std_logic;
signal \N__44912\ : std_logic;
signal \N__44909\ : std_logic;
signal \N__44906\ : std_logic;
signal \N__44901\ : std_logic;
signal \N__44900\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44890\ : std_logic;
signal \N__44887\ : std_logic;
signal \N__44884\ : std_logic;
signal \N__44881\ : std_logic;
signal \N__44878\ : std_logic;
signal \N__44875\ : std_logic;
signal \N__44872\ : std_logic;
signal \N__44869\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44859\ : std_logic;
signal \N__44858\ : std_logic;
signal \N__44857\ : std_logic;
signal \N__44852\ : std_logic;
signal \N__44849\ : std_logic;
signal \N__44846\ : std_logic;
signal \N__44841\ : std_logic;
signal \N__44838\ : std_logic;
signal \N__44835\ : std_logic;
signal \N__44832\ : std_logic;
signal \N__44829\ : std_logic;
signal \N__44826\ : std_logic;
signal \N__44825\ : std_logic;
signal \N__44822\ : std_logic;
signal \N__44819\ : std_logic;
signal \N__44816\ : std_logic;
signal \N__44813\ : std_logic;
signal \N__44812\ : std_logic;
signal \N__44809\ : std_logic;
signal \N__44806\ : std_logic;
signal \N__44803\ : std_logic;
signal \N__44802\ : std_logic;
signal \N__44797\ : std_logic;
signal \N__44792\ : std_logic;
signal \N__44789\ : std_logic;
signal \N__44786\ : std_logic;
signal \N__44781\ : std_logic;
signal \N__44778\ : std_logic;
signal \N__44775\ : std_logic;
signal \N__44774\ : std_logic;
signal \N__44773\ : std_logic;
signal \N__44770\ : std_logic;
signal \N__44767\ : std_logic;
signal \N__44764\ : std_logic;
signal \N__44757\ : std_logic;
signal \N__44754\ : std_logic;
signal \N__44751\ : std_logic;
signal \N__44748\ : std_logic;
signal \N__44745\ : std_logic;
signal \N__44742\ : std_logic;
signal \N__44741\ : std_logic;
signal \N__44740\ : std_logic;
signal \N__44737\ : std_logic;
signal \N__44734\ : std_logic;
signal \N__44733\ : std_logic;
signal \N__44732\ : std_logic;
signal \N__44729\ : std_logic;
signal \N__44726\ : std_logic;
signal \N__44723\ : std_logic;
signal \N__44718\ : std_logic;
signal \N__44715\ : std_logic;
signal \N__44712\ : std_logic;
signal \N__44709\ : std_logic;
signal \N__44706\ : std_logic;
signal \N__44701\ : std_logic;
signal \N__44694\ : std_logic;
signal \N__44691\ : std_logic;
signal \N__44688\ : std_logic;
signal \N__44685\ : std_logic;
signal \N__44682\ : std_logic;
signal \N__44679\ : std_logic;
signal \N__44676\ : std_logic;
signal \N__44675\ : std_logic;
signal \N__44672\ : std_logic;
signal \N__44671\ : std_logic;
signal \N__44668\ : std_logic;
signal \N__44665\ : std_logic;
signal \N__44662\ : std_logic;
signal \N__44659\ : std_logic;
signal \N__44656\ : std_logic;
signal \N__44653\ : std_logic;
signal \N__44652\ : std_logic;
signal \N__44649\ : std_logic;
signal \N__44644\ : std_logic;
signal \N__44641\ : std_logic;
signal \N__44634\ : std_logic;
signal \N__44631\ : std_logic;
signal \N__44628\ : std_logic;
signal \N__44627\ : std_logic;
signal \N__44626\ : std_logic;
signal \N__44623\ : std_logic;
signal \N__44620\ : std_logic;
signal \N__44617\ : std_logic;
signal \N__44610\ : std_logic;
signal \N__44607\ : std_logic;
signal \N__44604\ : std_logic;
signal \N__44601\ : std_logic;
signal \N__44598\ : std_logic;
signal \N__44597\ : std_logic;
signal \N__44596\ : std_logic;
signal \N__44595\ : std_logic;
signal \N__44594\ : std_logic;
signal \N__44593\ : std_logic;
signal \N__44592\ : std_logic;
signal \N__44591\ : std_logic;
signal \N__44590\ : std_logic;
signal \N__44589\ : std_logic;
signal \N__44588\ : std_logic;
signal \N__44587\ : std_logic;
signal \N__44586\ : std_logic;
signal \N__44585\ : std_logic;
signal \N__44584\ : std_logic;
signal \N__44583\ : std_logic;
signal \N__44582\ : std_logic;
signal \N__44581\ : std_logic;
signal \N__44580\ : std_logic;
signal \N__44577\ : std_logic;
signal \N__44576\ : std_logic;
signal \N__44575\ : std_logic;
signal \N__44574\ : std_logic;
signal \N__44571\ : std_logic;
signal \N__44570\ : std_logic;
signal \N__44569\ : std_logic;
signal \N__44566\ : std_logic;
signal \N__44565\ : std_logic;
signal \N__44560\ : std_logic;
signal \N__44559\ : std_logic;
signal \N__44556\ : std_logic;
signal \N__44555\ : std_logic;
signal \N__44554\ : std_logic;
signal \N__44551\ : std_logic;
signal \N__44548\ : std_logic;
signal \N__44545\ : std_logic;
signal \N__44542\ : std_logic;
signal \N__44539\ : std_logic;
signal \N__44536\ : std_logic;
signal \N__44535\ : std_logic;
signal \N__44532\ : std_logic;
signal \N__44531\ : std_logic;
signal \N__44528\ : std_logic;
signal \N__44525\ : std_logic;
signal \N__44524\ : std_logic;
signal \N__44523\ : std_logic;
signal \N__44522\ : std_logic;
signal \N__44519\ : std_logic;
signal \N__44518\ : std_logic;
signal \N__44517\ : std_logic;
signal \N__44516\ : std_logic;
signal \N__44515\ : std_logic;
signal \N__44514\ : std_logic;
signal \N__44513\ : std_logic;
signal \N__44512\ : std_logic;
signal \N__44511\ : std_logic;
signal \N__44510\ : std_logic;
signal \N__44505\ : std_logic;
signal \N__44502\ : std_logic;
signal \N__44499\ : std_logic;
signal \N__44496\ : std_logic;
signal \N__44495\ : std_logic;
signal \N__44492\ : std_logic;
signal \N__44481\ : std_logic;
signal \N__44478\ : std_logic;
signal \N__44475\ : std_logic;
signal \N__44474\ : std_logic;
signal \N__44461\ : std_logic;
signal \N__44458\ : std_logic;
signal \N__44453\ : std_logic;
signal \N__44450\ : std_logic;
signal \N__44447\ : std_logic;
signal \N__44444\ : std_logic;
signal \N__44427\ : std_logic;
signal \N__44420\ : std_logic;
signal \N__44417\ : std_logic;
signal \N__44414\ : std_logic;
signal \N__44407\ : std_logic;
signal \N__44404\ : std_logic;
signal \N__44401\ : std_logic;
signal \N__44400\ : std_logic;
signal \N__44397\ : std_logic;
signal \N__44394\ : std_logic;
signal \N__44391\ : std_logic;
signal \N__44386\ : std_logic;
signal \N__44381\ : std_logic;
signal \N__44380\ : std_logic;
signal \N__44377\ : std_logic;
signal \N__44376\ : std_logic;
signal \N__44375\ : std_logic;
signal \N__44374\ : std_logic;
signal \N__44371\ : std_logic;
signal \N__44368\ : std_logic;
signal \N__44365\ : std_logic;
signal \N__44358\ : std_logic;
signal \N__44353\ : std_logic;
signal \N__44342\ : std_logic;
signal \N__44339\ : std_logic;
signal \N__44336\ : std_logic;
signal \N__44333\ : std_logic;
signal \N__44330\ : std_logic;
signal \N__44325\ : std_logic;
signal \N__44314\ : std_logic;
signal \N__44305\ : std_logic;
signal \N__44300\ : std_logic;
signal \N__44283\ : std_logic;
signal \N__44282\ : std_logic;
signal \N__44279\ : std_logic;
signal \N__44276\ : std_logic;
signal \N__44273\ : std_logic;
signal \N__44270\ : std_logic;
signal \N__44269\ : std_logic;
signal \N__44266\ : std_logic;
signal \N__44263\ : std_logic;
signal \N__44260\ : std_logic;
signal \N__44257\ : std_logic;
signal \N__44254\ : std_logic;
signal \N__44247\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44243\ : std_logic;
signal \N__44240\ : std_logic;
signal \N__44237\ : std_logic;
signal \N__44236\ : std_logic;
signal \N__44233\ : std_logic;
signal \N__44230\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44220\ : std_logic;
signal \N__44217\ : std_logic;
signal \N__44216\ : std_logic;
signal \N__44213\ : std_logic;
signal \N__44212\ : std_logic;
signal \N__44209\ : std_logic;
signal \N__44206\ : std_logic;
signal \N__44203\ : std_logic;
signal \N__44200\ : std_logic;
signal \N__44199\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44191\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44181\ : std_logic;
signal \N__44178\ : std_logic;
signal \N__44175\ : std_logic;
signal \N__44172\ : std_logic;
signal \N__44169\ : std_logic;
signal \N__44166\ : std_logic;
signal \N__44163\ : std_logic;
signal \N__44160\ : std_logic;
signal \N__44159\ : std_logic;
signal \N__44156\ : std_logic;
signal \N__44155\ : std_logic;
signal \N__44152\ : std_logic;
signal \N__44149\ : std_logic;
signal \N__44146\ : std_logic;
signal \N__44143\ : std_logic;
signal \N__44136\ : std_logic;
signal \N__44135\ : std_logic;
signal \N__44134\ : std_logic;
signal \N__44133\ : std_logic;
signal \N__44132\ : std_logic;
signal \N__44131\ : std_logic;
signal \N__44130\ : std_logic;
signal \N__44129\ : std_logic;
signal \N__44128\ : std_logic;
signal \N__44109\ : std_logic;
signal \N__44106\ : std_logic;
signal \N__44103\ : std_logic;
signal \N__44102\ : std_logic;
signal \N__44099\ : std_logic;
signal \N__44094\ : std_logic;
signal \N__44093\ : std_logic;
signal \N__44090\ : std_logic;
signal \N__44087\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44081\ : std_logic;
signal \N__44078\ : std_logic;
signal \N__44075\ : std_logic;
signal \N__44070\ : std_logic;
signal \N__44067\ : std_logic;
signal \N__44064\ : std_logic;
signal \N__44061\ : std_logic;
signal \N__44058\ : std_logic;
signal \N__44055\ : std_logic;
signal \N__44054\ : std_logic;
signal \N__44053\ : std_logic;
signal \N__44052\ : std_logic;
signal \N__44051\ : std_logic;
signal \N__44050\ : std_logic;
signal \N__44049\ : std_logic;
signal \N__44048\ : std_logic;
signal \N__44047\ : std_logic;
signal \N__44046\ : std_logic;
signal \N__44045\ : std_logic;
signal \N__44042\ : std_logic;
signal \N__44041\ : std_logic;
signal \N__44040\ : std_logic;
signal \N__44039\ : std_logic;
signal \N__44038\ : std_logic;
signal \N__44037\ : std_logic;
signal \N__44036\ : std_logic;
signal \N__44033\ : std_logic;
signal \N__44028\ : std_logic;
signal \N__44025\ : std_logic;
signal \N__44024\ : std_logic;
signal \N__44023\ : std_logic;
signal \N__44022\ : std_logic;
signal \N__44021\ : std_logic;
signal \N__44020\ : std_logic;
signal \N__44019\ : std_logic;
signal \N__44018\ : std_logic;
signal \N__44017\ : std_logic;
signal \N__44004\ : std_logic;
signal \N__44001\ : std_logic;
signal \N__43992\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43984\ : std_logic;
signal \N__43981\ : std_logic;
signal \N__43978\ : std_logic;
signal \N__43975\ : std_logic;
signal \N__43960\ : std_logic;
signal \N__43955\ : std_logic;
signal \N__43952\ : std_logic;
signal \N__43945\ : std_logic;
signal \N__43932\ : std_logic;
signal \N__43931\ : std_logic;
signal \N__43928\ : std_logic;
signal \N__43927\ : std_logic;
signal \N__43920\ : std_logic;
signal \N__43917\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43915\ : std_logic;
signal \N__43914\ : std_logic;
signal \N__43907\ : std_logic;
signal \N__43904\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43896\ : std_logic;
signal \N__43893\ : std_logic;
signal \N__43890\ : std_logic;
signal \N__43887\ : std_logic;
signal \N__43884\ : std_logic;
signal \N__43881\ : std_logic;
signal \N__43878\ : std_logic;
signal \N__43875\ : std_logic;
signal \N__43872\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43863\ : std_logic;
signal \N__43860\ : std_logic;
signal \N__43857\ : std_logic;
signal \N__43854\ : std_logic;
signal \N__43851\ : std_logic;
signal \N__43850\ : std_logic;
signal \N__43847\ : std_logic;
signal \N__43844\ : std_logic;
signal \N__43843\ : std_logic;
signal \N__43842\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43836\ : std_logic;
signal \N__43831\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43823\ : std_logic;
signal \N__43818\ : std_logic;
signal \N__43817\ : std_logic;
signal \N__43816\ : std_logic;
signal \N__43813\ : std_logic;
signal \N__43808\ : std_logic;
signal \N__43803\ : std_logic;
signal \N__43800\ : std_logic;
signal \N__43797\ : std_logic;
signal \N__43794\ : std_logic;
signal \N__43791\ : std_logic;
signal \N__43788\ : std_logic;
signal \N__43785\ : std_logic;
signal \N__43782\ : std_logic;
signal \N__43779\ : std_logic;
signal \N__43776\ : std_logic;
signal \N__43775\ : std_logic;
signal \N__43774\ : std_logic;
signal \N__43773\ : std_logic;
signal \N__43770\ : std_logic;
signal \N__43765\ : std_logic;
signal \N__43762\ : std_logic;
signal \N__43759\ : std_logic;
signal \N__43756\ : std_logic;
signal \N__43753\ : std_logic;
signal \N__43750\ : std_logic;
signal \N__43747\ : std_logic;
signal \N__43740\ : std_logic;
signal \N__43737\ : std_logic;
signal \N__43736\ : std_logic;
signal \N__43733\ : std_logic;
signal \N__43732\ : std_logic;
signal \N__43729\ : std_logic;
signal \N__43726\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43718\ : std_logic;
signal \N__43713\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43707\ : std_logic;
signal \N__43704\ : std_logic;
signal \N__43701\ : std_logic;
signal \N__43700\ : std_logic;
signal \N__43697\ : std_logic;
signal \N__43694\ : std_logic;
signal \N__43693\ : std_logic;
signal \N__43690\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43684\ : std_logic;
signal \N__43683\ : std_logic;
signal \N__43680\ : std_logic;
signal \N__43677\ : std_logic;
signal \N__43674\ : std_logic;
signal \N__43671\ : std_logic;
signal \N__43668\ : std_logic;
signal \N__43663\ : std_logic;
signal \N__43660\ : std_logic;
signal \N__43657\ : std_logic;
signal \N__43654\ : std_logic;
signal \N__43647\ : std_logic;
signal \N__43646\ : std_logic;
signal \N__43643\ : std_logic;
signal \N__43642\ : std_logic;
signal \N__43639\ : std_logic;
signal \N__43636\ : std_logic;
signal \N__43633\ : std_logic;
signal \N__43626\ : std_logic;
signal \N__43623\ : std_logic;
signal \N__43620\ : std_logic;
signal \N__43617\ : std_logic;
signal \N__43614\ : std_logic;
signal \N__43611\ : std_logic;
signal \N__43608\ : std_logic;
signal \N__43607\ : std_logic;
signal \N__43604\ : std_logic;
signal \N__43603\ : std_logic;
signal \N__43600\ : std_logic;
signal \N__43597\ : std_logic;
signal \N__43594\ : std_logic;
signal \N__43591\ : std_logic;
signal \N__43588\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43580\ : std_logic;
signal \N__43579\ : std_logic;
signal \N__43576\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43570\ : std_logic;
signal \N__43563\ : std_logic;
signal \N__43560\ : std_logic;
signal \N__43557\ : std_logic;
signal \N__43554\ : std_logic;
signal \N__43553\ : std_logic;
signal \N__43552\ : std_logic;
signal \N__43549\ : std_logic;
signal \N__43546\ : std_logic;
signal \N__43543\ : std_logic;
signal \N__43536\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43530\ : std_logic;
signal \N__43527\ : std_logic;
signal \N__43524\ : std_logic;
signal \N__43521\ : std_logic;
signal \N__43518\ : std_logic;
signal \N__43515\ : std_logic;
signal \N__43512\ : std_logic;
signal \N__43509\ : std_logic;
signal \N__43506\ : std_logic;
signal \N__43503\ : std_logic;
signal \N__43502\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43496\ : std_logic;
signal \N__43493\ : std_logic;
signal \N__43490\ : std_logic;
signal \N__43489\ : std_logic;
signal \N__43488\ : std_logic;
signal \N__43485\ : std_logic;
signal \N__43482\ : std_logic;
signal \N__43477\ : std_logic;
signal \N__43474\ : std_logic;
signal \N__43469\ : std_logic;
signal \N__43464\ : std_logic;
signal \N__43461\ : std_logic;
signal \N__43458\ : std_logic;
signal \N__43457\ : std_logic;
signal \N__43456\ : std_logic;
signal \N__43453\ : std_logic;
signal \N__43450\ : std_logic;
signal \N__43447\ : std_logic;
signal \N__43440\ : std_logic;
signal \N__43437\ : std_logic;
signal \N__43434\ : std_logic;
signal \N__43431\ : std_logic;
signal \N__43428\ : std_logic;
signal \N__43425\ : std_logic;
signal \N__43422\ : std_logic;
signal \N__43421\ : std_logic;
signal \N__43418\ : std_logic;
signal \N__43415\ : std_logic;
signal \N__43414\ : std_logic;
signal \N__43413\ : std_logic;
signal \N__43410\ : std_logic;
signal \N__43407\ : std_logic;
signal \N__43402\ : std_logic;
signal \N__43399\ : std_logic;
signal \N__43396\ : std_logic;
signal \N__43393\ : std_logic;
signal \N__43386\ : std_logic;
signal \N__43385\ : std_logic;
signal \N__43382\ : std_logic;
signal \N__43379\ : std_logic;
signal \N__43378\ : std_logic;
signal \N__43375\ : std_logic;
signal \N__43372\ : std_logic;
signal \N__43369\ : std_logic;
signal \N__43364\ : std_logic;
signal \N__43359\ : std_logic;
signal \N__43356\ : std_logic;
signal \N__43353\ : std_logic;
signal \N__43350\ : std_logic;
signal \N__43347\ : std_logic;
signal \N__43344\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43338\ : std_logic;
signal \N__43335\ : std_logic;
signal \N__43334\ : std_logic;
signal \N__43331\ : std_logic;
signal \N__43328\ : std_logic;
signal \N__43327\ : std_logic;
signal \N__43322\ : std_logic;
signal \N__43319\ : std_logic;
signal \N__43314\ : std_logic;
signal \N__43313\ : std_logic;
signal \N__43312\ : std_logic;
signal \N__43309\ : std_logic;
signal \N__43306\ : std_logic;
signal \N__43303\ : std_logic;
signal \N__43302\ : std_logic;
signal \N__43299\ : std_logic;
signal \N__43296\ : std_logic;
signal \N__43291\ : std_logic;
signal \N__43284\ : std_logic;
signal \N__43281\ : std_logic;
signal \N__43278\ : std_logic;
signal \N__43275\ : std_logic;
signal \N__43272\ : std_logic;
signal \N__43269\ : std_logic;
signal \N__43266\ : std_logic;
signal \N__43263\ : std_logic;
signal \N__43260\ : std_logic;
signal \N__43257\ : std_logic;
signal \N__43254\ : std_logic;
signal \N__43251\ : std_logic;
signal \N__43248\ : std_logic;
signal \N__43245\ : std_logic;
signal \N__43242\ : std_logic;
signal \N__43241\ : std_logic;
signal \N__43238\ : std_logic;
signal \N__43235\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43227\ : std_logic;
signal \N__43224\ : std_logic;
signal \N__43221\ : std_logic;
signal \N__43220\ : std_logic;
signal \N__43217\ : std_logic;
signal \N__43214\ : std_logic;
signal \N__43209\ : std_logic;
signal \N__43206\ : std_logic;
signal \N__43203\ : std_logic;
signal \N__43200\ : std_logic;
signal \N__43199\ : std_logic;
signal \N__43196\ : std_logic;
signal \N__43193\ : std_logic;
signal \N__43190\ : std_logic;
signal \N__43187\ : std_logic;
signal \N__43182\ : std_logic;
signal \N__43179\ : std_logic;
signal \N__43176\ : std_logic;
signal \N__43173\ : std_logic;
signal \N__43170\ : std_logic;
signal \N__43169\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43163\ : std_logic;
signal \N__43158\ : std_logic;
signal \N__43155\ : std_logic;
signal \N__43152\ : std_logic;
signal \N__43151\ : std_logic;
signal \N__43148\ : std_logic;
signal \N__43145\ : std_logic;
signal \N__43142\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43134\ : std_logic;
signal \N__43131\ : std_logic;
signal \N__43128\ : std_logic;
signal \N__43125\ : std_logic;
signal \N__43124\ : std_logic;
signal \N__43121\ : std_logic;
signal \N__43118\ : std_logic;
signal \N__43113\ : std_logic;
signal \N__43110\ : std_logic;
signal \N__43109\ : std_logic;
signal \N__43106\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43100\ : std_logic;
signal \N__43097\ : std_logic;
signal \N__43092\ : std_logic;
signal \N__43089\ : std_logic;
signal \N__43088\ : std_logic;
signal \N__43085\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43076\ : std_logic;
signal \N__43071\ : std_logic;
signal \N__43068\ : std_logic;
signal \N__43067\ : std_logic;
signal \N__43066\ : std_logic;
signal \N__43063\ : std_logic;
signal \N__43062\ : std_logic;
signal \N__43057\ : std_logic;
signal \N__43054\ : std_logic;
signal \N__43051\ : std_logic;
signal \N__43048\ : std_logic;
signal \N__43041\ : std_logic;
signal \N__43038\ : std_logic;
signal \N__43037\ : std_logic;
signal \N__43034\ : std_logic;
signal \N__43031\ : std_logic;
signal \N__43028\ : std_logic;
signal \N__43025\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43019\ : std_logic;
signal \N__43016\ : std_logic;
signal \N__43011\ : std_logic;
signal \N__43008\ : std_logic;
signal \N__43007\ : std_logic;
signal \N__43006\ : std_logic;
signal \N__43003\ : std_logic;
signal \N__43000\ : std_logic;
signal \N__42997\ : std_logic;
signal \N__42994\ : std_logic;
signal \N__42991\ : std_logic;
signal \N__42988\ : std_logic;
signal \N__42981\ : std_logic;
signal \N__42978\ : std_logic;
signal \N__42975\ : std_logic;
signal \N__42974\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42967\ : std_logic;
signal \N__42964\ : std_logic;
signal \N__42961\ : std_logic;
signal \N__42958\ : std_logic;
signal \N__42951\ : std_logic;
signal \N__42948\ : std_logic;
signal \N__42945\ : std_logic;
signal \N__42942\ : std_logic;
signal \N__42941\ : std_logic;
signal \N__42940\ : std_logic;
signal \N__42937\ : std_logic;
signal \N__42934\ : std_logic;
signal \N__42931\ : std_logic;
signal \N__42924\ : std_logic;
signal \N__42921\ : std_logic;
signal \N__42918\ : std_logic;
signal \N__42915\ : std_logic;
signal \N__42912\ : std_logic;
signal \N__42909\ : std_logic;
signal \N__42908\ : std_logic;
signal \N__42905\ : std_logic;
signal \N__42902\ : std_logic;
signal \N__42897\ : std_logic;
signal \N__42894\ : std_logic;
signal \N__42891\ : std_logic;
signal \N__42890\ : std_logic;
signal \N__42889\ : std_logic;
signal \N__42886\ : std_logic;
signal \N__42881\ : std_logic;
signal \N__42876\ : std_logic;
signal \N__42873\ : std_logic;
signal \N__42870\ : std_logic;
signal \N__42869\ : std_logic;
signal \N__42868\ : std_logic;
signal \N__42865\ : std_logic;
signal \N__42860\ : std_logic;
signal \N__42857\ : std_logic;
signal \N__42854\ : std_logic;
signal \N__42849\ : std_logic;
signal \N__42846\ : std_logic;
signal \N__42843\ : std_logic;
signal \N__42840\ : std_logic;
signal \N__42837\ : std_logic;
signal \N__42834\ : std_logic;
signal \N__42831\ : std_logic;
signal \N__42830\ : std_logic;
signal \N__42829\ : std_logic;
signal \N__42826\ : std_logic;
signal \N__42825\ : std_logic;
signal \N__42822\ : std_logic;
signal \N__42819\ : std_logic;
signal \N__42816\ : std_logic;
signal \N__42813\ : std_logic;
signal \N__42810\ : std_logic;
signal \N__42807\ : std_logic;
signal \N__42798\ : std_logic;
signal \N__42795\ : std_logic;
signal \N__42792\ : std_logic;
signal \N__42791\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42785\ : std_logic;
signal \N__42780\ : std_logic;
signal \N__42777\ : std_logic;
signal \N__42774\ : std_logic;
signal \N__42773\ : std_logic;
signal \N__42770\ : std_logic;
signal \N__42767\ : std_logic;
signal \N__42762\ : std_logic;
signal \N__42759\ : std_logic;
signal \N__42756\ : std_logic;
signal \N__42755\ : std_logic;
signal \N__42752\ : std_logic;
signal \N__42749\ : std_logic;
signal \N__42746\ : std_logic;
signal \N__42743\ : std_logic;
signal \N__42738\ : std_logic;
signal \N__42735\ : std_logic;
signal \N__42732\ : std_logic;
signal \N__42729\ : std_logic;
signal \N__42728\ : std_logic;
signal \N__42725\ : std_logic;
signal \N__42722\ : std_logic;
signal \N__42717\ : std_logic;
signal \N__42714\ : std_logic;
signal \N__42711\ : std_logic;
signal \N__42708\ : std_logic;
signal \N__42705\ : std_logic;
signal \N__42702\ : std_logic;
signal \N__42699\ : std_logic;
signal \N__42696\ : std_logic;
signal \N__42693\ : std_logic;
signal \N__42690\ : std_logic;
signal \N__42687\ : std_logic;
signal \N__42684\ : std_logic;
signal \N__42681\ : std_logic;
signal \N__42678\ : std_logic;
signal \N__42675\ : std_logic;
signal \N__42672\ : std_logic;
signal \N__42671\ : std_logic;
signal \N__42668\ : std_logic;
signal \N__42665\ : std_logic;
signal \N__42660\ : std_logic;
signal \N__42657\ : std_logic;
signal \N__42654\ : std_logic;
signal \N__42653\ : std_logic;
signal \N__42652\ : std_logic;
signal \N__42649\ : std_logic;
signal \N__42644\ : std_logic;
signal \N__42639\ : std_logic;
signal \N__42636\ : std_logic;
signal \N__42635\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42629\ : std_logic;
signal \N__42624\ : std_logic;
signal \N__42621\ : std_logic;
signal \N__42618\ : std_logic;
signal \N__42617\ : std_logic;
signal \N__42614\ : std_logic;
signal \N__42611\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42603\ : std_logic;
signal \N__42600\ : std_logic;
signal \N__42599\ : std_logic;
signal \N__42596\ : std_logic;
signal \N__42593\ : std_logic;
signal \N__42588\ : std_logic;
signal \N__42585\ : std_logic;
signal \N__42582\ : std_logic;
signal \N__42579\ : std_logic;
signal \N__42578\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42572\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42564\ : std_logic;
signal \N__42561\ : std_logic;
signal \N__42560\ : std_logic;
signal \N__42557\ : std_logic;
signal \N__42556\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42554\ : std_logic;
signal \N__42551\ : std_logic;
signal \N__42548\ : std_logic;
signal \N__42545\ : std_logic;
signal \N__42542\ : std_logic;
signal \N__42539\ : std_logic;
signal \N__42528\ : std_logic;
signal \N__42525\ : std_logic;
signal \N__42522\ : std_logic;
signal \N__42521\ : std_logic;
signal \N__42518\ : std_logic;
signal \N__42517\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42515\ : std_logic;
signal \N__42512\ : std_logic;
signal \N__42509\ : std_logic;
signal \N__42506\ : std_logic;
signal \N__42503\ : std_logic;
signal \N__42500\ : std_logic;
signal \N__42489\ : std_logic;
signal \N__42486\ : std_logic;
signal \N__42485\ : std_logic;
signal \N__42482\ : std_logic;
signal \N__42479\ : std_logic;
signal \N__42474\ : std_logic;
signal \N__42471\ : std_logic;
signal \N__42468\ : std_logic;
signal \N__42467\ : std_logic;
signal \N__42464\ : std_logic;
signal \N__42461\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42450\ : std_logic;
signal \N__42449\ : std_logic;
signal \N__42446\ : std_logic;
signal \N__42443\ : std_logic;
signal \N__42442\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42436\ : std_logic;
signal \N__42433\ : std_logic;
signal \N__42430\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42417\ : std_logic;
signal \N__42414\ : std_logic;
signal \N__42411\ : std_logic;
signal \N__42408\ : std_logic;
signal \N__42405\ : std_logic;
signal \N__42404\ : std_logic;
signal \N__42401\ : std_logic;
signal \N__42398\ : std_logic;
signal \N__42397\ : std_logic;
signal \N__42392\ : std_logic;
signal \N__42389\ : std_logic;
signal \N__42388\ : std_logic;
signal \N__42385\ : std_logic;
signal \N__42382\ : std_logic;
signal \N__42379\ : std_logic;
signal \N__42372\ : std_logic;
signal \N__42369\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42360\ : std_logic;
signal \N__42357\ : std_logic;
signal \N__42356\ : std_logic;
signal \N__42353\ : std_logic;
signal \N__42350\ : std_logic;
signal \N__42345\ : std_logic;
signal \N__42342\ : std_logic;
signal \N__42339\ : std_logic;
signal \N__42336\ : std_logic;
signal \N__42335\ : std_logic;
signal \N__42334\ : std_logic;
signal \N__42331\ : std_logic;
signal \N__42328\ : std_logic;
signal \N__42325\ : std_logic;
signal \N__42322\ : std_logic;
signal \N__42321\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42315\ : std_logic;
signal \N__42312\ : std_logic;
signal \N__42309\ : std_logic;
signal \N__42300\ : std_logic;
signal \N__42297\ : std_logic;
signal \N__42294\ : std_logic;
signal \N__42291\ : std_logic;
signal \N__42288\ : std_logic;
signal \N__42285\ : std_logic;
signal \N__42282\ : std_logic;
signal \N__42279\ : std_logic;
signal \N__42276\ : std_logic;
signal \N__42273\ : std_logic;
signal \N__42270\ : std_logic;
signal \N__42267\ : std_logic;
signal \N__42266\ : std_logic;
signal \N__42263\ : std_logic;
signal \N__42260\ : std_logic;
signal \N__42257\ : std_logic;
signal \N__42254\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42248\ : std_logic;
signal \N__42245\ : std_logic;
signal \N__42242\ : std_logic;
signal \N__42239\ : std_logic;
signal \N__42234\ : std_logic;
signal \N__42231\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42229\ : std_logic;
signal \N__42226\ : std_logic;
signal \N__42225\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42216\ : std_logic;
signal \N__42213\ : std_logic;
signal \N__42204\ : std_logic;
signal \N__42203\ : std_logic;
signal \N__42200\ : std_logic;
signal \N__42199\ : std_logic;
signal \N__42196\ : std_logic;
signal \N__42193\ : std_logic;
signal \N__42190\ : std_logic;
signal \N__42183\ : std_logic;
signal \N__42180\ : std_logic;
signal \N__42177\ : std_logic;
signal \N__42174\ : std_logic;
signal \N__42171\ : std_logic;
signal \N__42170\ : std_logic;
signal \N__42169\ : std_logic;
signal \N__42168\ : std_logic;
signal \N__42165\ : std_logic;
signal \N__42162\ : std_logic;
signal \N__42159\ : std_logic;
signal \N__42158\ : std_logic;
signal \N__42155\ : std_logic;
signal \N__42152\ : std_logic;
signal \N__42149\ : std_logic;
signal \N__42146\ : std_logic;
signal \N__42143\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42129\ : std_logic;
signal \N__42128\ : std_logic;
signal \N__42127\ : std_logic;
signal \N__42124\ : std_logic;
signal \N__42123\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42117\ : std_logic;
signal \N__42114\ : std_logic;
signal \N__42111\ : std_logic;
signal \N__42106\ : std_logic;
signal \N__42105\ : std_logic;
signal \N__42102\ : std_logic;
signal \N__42097\ : std_logic;
signal \N__42094\ : std_logic;
signal \N__42087\ : std_logic;
signal \N__42084\ : std_logic;
signal \N__42081\ : std_logic;
signal \N__42078\ : std_logic;
signal \N__42075\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42069\ : std_logic;
signal \N__42066\ : std_logic;
signal \N__42063\ : std_logic;
signal \N__42060\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42051\ : std_logic;
signal \N__42048\ : std_logic;
signal \N__42045\ : std_logic;
signal \N__42042\ : std_logic;
signal \N__42039\ : std_logic;
signal \N__42036\ : std_logic;
signal \N__42033\ : std_logic;
signal \N__42030\ : std_logic;
signal \N__42027\ : std_logic;
signal \N__42024\ : std_logic;
signal \N__42021\ : std_logic;
signal \N__42018\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42009\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__42000\ : std_logic;
signal \N__41997\ : std_logic;
signal \N__41994\ : std_logic;
signal \N__41991\ : std_logic;
signal \N__41988\ : std_logic;
signal \N__41985\ : std_logic;
signal \N__41982\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41976\ : std_logic;
signal \N__41973\ : std_logic;
signal \N__41970\ : std_logic;
signal \N__41967\ : std_logic;
signal \N__41964\ : std_logic;
signal \N__41961\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41955\ : std_logic;
signal \N__41952\ : std_logic;
signal \N__41949\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41940\ : std_logic;
signal \N__41937\ : std_logic;
signal \N__41934\ : std_logic;
signal \N__41931\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41925\ : std_logic;
signal \N__41922\ : std_logic;
signal \N__41919\ : std_logic;
signal \N__41916\ : std_logic;
signal \N__41913\ : std_logic;
signal \N__41910\ : std_logic;
signal \N__41907\ : std_logic;
signal \N__41904\ : std_logic;
signal \N__41901\ : std_logic;
signal \N__41898\ : std_logic;
signal \N__41895\ : std_logic;
signal \N__41892\ : std_logic;
signal \N__41889\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41877\ : std_logic;
signal \N__41874\ : std_logic;
signal \N__41871\ : std_logic;
signal \N__41868\ : std_logic;
signal \N__41865\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41859\ : std_logic;
signal \N__41856\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41850\ : std_logic;
signal \N__41847\ : std_logic;
signal \N__41844\ : std_logic;
signal \N__41841\ : std_logic;
signal \N__41838\ : std_logic;
signal \N__41835\ : std_logic;
signal \N__41832\ : std_logic;
signal \N__41829\ : std_logic;
signal \N__41826\ : std_logic;
signal \N__41823\ : std_logic;
signal \N__41820\ : std_logic;
signal \N__41817\ : std_logic;
signal \N__41814\ : std_logic;
signal \N__41811\ : std_logic;
signal \N__41808\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41802\ : std_logic;
signal \N__41799\ : std_logic;
signal \N__41796\ : std_logic;
signal \N__41793\ : std_logic;
signal \N__41790\ : std_logic;
signal \N__41787\ : std_logic;
signal \N__41784\ : std_logic;
signal \N__41781\ : std_logic;
signal \N__41780\ : std_logic;
signal \N__41777\ : std_logic;
signal \N__41774\ : std_logic;
signal \N__41771\ : std_logic;
signal \N__41768\ : std_logic;
signal \N__41765\ : std_logic;
signal \N__41762\ : std_logic;
signal \N__41761\ : std_logic;
signal \N__41756\ : std_logic;
signal \N__41753\ : std_logic;
signal \N__41752\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41744\ : std_logic;
signal \N__41739\ : std_logic;
signal \N__41736\ : std_logic;
signal \N__41735\ : std_logic;
signal \N__41734\ : std_logic;
signal \N__41731\ : std_logic;
signal \N__41728\ : std_logic;
signal \N__41725\ : std_logic;
signal \N__41720\ : std_logic;
signal \N__41717\ : std_logic;
signal \N__41714\ : std_logic;
signal \N__41709\ : std_logic;
signal \N__41708\ : std_logic;
signal \N__41705\ : std_logic;
signal \N__41702\ : std_logic;
signal \N__41701\ : std_logic;
signal \N__41698\ : std_logic;
signal \N__41697\ : std_logic;
signal \N__41694\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41680\ : std_logic;
signal \N__41677\ : std_logic;
signal \N__41674\ : std_logic;
signal \N__41671\ : std_logic;
signal \N__41666\ : std_logic;
signal \N__41661\ : std_logic;
signal \N__41658\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41656\ : std_logic;
signal \N__41653\ : std_logic;
signal \N__41650\ : std_logic;
signal \N__41647\ : std_logic;
signal \N__41642\ : std_logic;
signal \N__41637\ : std_logic;
signal \N__41634\ : std_logic;
signal \N__41633\ : std_logic;
signal \N__41630\ : std_logic;
signal \N__41627\ : std_logic;
signal \N__41624\ : std_logic;
signal \N__41621\ : std_logic;
signal \N__41616\ : std_logic;
signal \N__41613\ : std_logic;
signal \N__41612\ : std_logic;
signal \N__41609\ : std_logic;
signal \N__41606\ : std_logic;
signal \N__41603\ : std_logic;
signal \N__41600\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41592\ : std_logic;
signal \N__41589\ : std_logic;
signal \N__41586\ : std_logic;
signal \N__41583\ : std_logic;
signal \N__41580\ : std_logic;
signal \N__41577\ : std_logic;
signal \N__41574\ : std_logic;
signal \N__41571\ : std_logic;
signal \N__41568\ : std_logic;
signal \N__41565\ : std_logic;
signal \N__41562\ : std_logic;
signal \N__41559\ : std_logic;
signal \N__41556\ : std_logic;
signal \N__41553\ : std_logic;
signal \N__41550\ : std_logic;
signal \N__41549\ : std_logic;
signal \N__41548\ : std_logic;
signal \N__41541\ : std_logic;
signal \N__41538\ : std_logic;
signal \N__41535\ : std_logic;
signal \N__41532\ : std_logic;
signal \N__41529\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41520\ : std_logic;
signal \N__41517\ : std_logic;
signal \N__41514\ : std_logic;
signal \N__41511\ : std_logic;
signal \N__41508\ : std_logic;
signal \N__41505\ : std_logic;
signal \N__41502\ : std_logic;
signal \N__41499\ : std_logic;
signal \N__41496\ : std_logic;
signal \N__41493\ : std_logic;
signal \N__41490\ : std_logic;
signal \N__41487\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41481\ : std_logic;
signal \N__41480\ : std_logic;
signal \N__41477\ : std_logic;
signal \N__41474\ : std_logic;
signal \N__41473\ : std_logic;
signal \N__41468\ : std_logic;
signal \N__41465\ : std_logic;
signal \N__41462\ : std_logic;
signal \N__41459\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41451\ : std_logic;
signal \N__41448\ : std_logic;
signal \N__41445\ : std_logic;
signal \N__41442\ : std_logic;
signal \N__41439\ : std_logic;
signal \N__41438\ : std_logic;
signal \N__41435\ : std_logic;
signal \N__41432\ : std_logic;
signal \N__41431\ : std_logic;
signal \N__41428\ : std_logic;
signal \N__41425\ : std_logic;
signal \N__41422\ : std_logic;
signal \N__41419\ : std_logic;
signal \N__41414\ : std_logic;
signal \N__41409\ : std_logic;
signal \N__41406\ : std_logic;
signal \N__41403\ : std_logic;
signal \N__41400\ : std_logic;
signal \N__41397\ : std_logic;
signal \N__41394\ : std_logic;
signal \N__41391\ : std_logic;
signal \N__41390\ : std_logic;
signal \N__41387\ : std_logic;
signal \N__41384\ : std_logic;
signal \N__41383\ : std_logic;
signal \N__41380\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41367\ : std_logic;
signal \N__41364\ : std_logic;
signal \N__41361\ : std_logic;
signal \N__41358\ : std_logic;
signal \N__41357\ : std_logic;
signal \N__41356\ : std_logic;
signal \N__41349\ : std_logic;
signal \N__41346\ : std_logic;
signal \N__41343\ : std_logic;
signal \N__41340\ : std_logic;
signal \N__41337\ : std_logic;
signal \N__41334\ : std_logic;
signal \N__41331\ : std_logic;
signal \N__41328\ : std_logic;
signal \N__41325\ : std_logic;
signal \N__41322\ : std_logic;
signal \N__41319\ : std_logic;
signal \N__41316\ : std_logic;
signal \N__41313\ : std_logic;
signal \N__41310\ : std_logic;
signal \N__41307\ : std_logic;
signal \N__41304\ : std_logic;
signal \N__41301\ : std_logic;
signal \N__41298\ : std_logic;
signal \N__41295\ : std_logic;
signal \N__41292\ : std_logic;
signal \N__41289\ : std_logic;
signal \N__41286\ : std_logic;
signal \N__41283\ : std_logic;
signal \N__41280\ : std_logic;
signal \N__41277\ : std_logic;
signal \N__41274\ : std_logic;
signal \N__41271\ : std_logic;
signal \N__41268\ : std_logic;
signal \N__41265\ : std_logic;
signal \N__41262\ : std_logic;
signal \N__41259\ : std_logic;
signal \N__41256\ : std_logic;
signal \N__41253\ : std_logic;
signal \N__41252\ : std_logic;
signal \N__41251\ : std_logic;
signal \N__41248\ : std_logic;
signal \N__41245\ : std_logic;
signal \N__41242\ : std_logic;
signal \N__41235\ : std_logic;
signal \N__41232\ : std_logic;
signal \N__41229\ : std_logic;
signal \N__41226\ : std_logic;
signal \N__41223\ : std_logic;
signal \N__41220\ : std_logic;
signal \N__41217\ : std_logic;
signal \N__41214\ : std_logic;
signal \N__41211\ : std_logic;
signal \N__41208\ : std_logic;
signal \N__41205\ : std_logic;
signal \N__41204\ : std_logic;
signal \N__41203\ : std_logic;
signal \N__41200\ : std_logic;
signal \N__41197\ : std_logic;
signal \N__41194\ : std_logic;
signal \N__41189\ : std_logic;
signal \N__41184\ : std_logic;
signal \N__41181\ : std_logic;
signal \N__41178\ : std_logic;
signal \N__41175\ : std_logic;
signal \N__41172\ : std_logic;
signal \N__41169\ : std_logic;
signal \N__41166\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41160\ : std_logic;
signal \N__41157\ : std_logic;
signal \N__41156\ : std_logic;
signal \N__41153\ : std_logic;
signal \N__41150\ : std_logic;
signal \N__41149\ : std_logic;
signal \N__41146\ : std_logic;
signal \N__41141\ : std_logic;
signal \N__41138\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41130\ : std_logic;
signal \N__41127\ : std_logic;
signal \N__41124\ : std_logic;
signal \N__41121\ : std_logic;
signal \N__41118\ : std_logic;
signal \N__41115\ : std_logic;
signal \N__41112\ : std_logic;
signal \N__41109\ : std_logic;
signal \N__41106\ : std_logic;
signal \N__41103\ : std_logic;
signal \N__41102\ : std_logic;
signal \N__41099\ : std_logic;
signal \N__41096\ : std_logic;
signal \N__41093\ : std_logic;
signal \N__41090\ : std_logic;
signal \N__41089\ : std_logic;
signal \N__41088\ : std_logic;
signal \N__41085\ : std_logic;
signal \N__41082\ : std_logic;
signal \N__41077\ : std_logic;
signal \N__41074\ : std_logic;
signal \N__41069\ : std_logic;
signal \N__41064\ : std_logic;
signal \N__41063\ : std_logic;
signal \N__41060\ : std_logic;
signal \N__41057\ : std_logic;
signal \N__41056\ : std_logic;
signal \N__41053\ : std_logic;
signal \N__41050\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41041\ : std_logic;
signal \N__41038\ : std_logic;
signal \N__41035\ : std_logic;
signal \N__41028\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41019\ : std_logic;
signal \N__41018\ : std_logic;
signal \N__41013\ : std_logic;
signal \N__41010\ : std_logic;
signal \N__41009\ : std_logic;
signal \N__41006\ : std_logic;
signal \N__41003\ : std_logic;
signal \N__40998\ : std_logic;
signal \N__40995\ : std_logic;
signal \N__40992\ : std_logic;
signal \N__40989\ : std_logic;
signal \N__40986\ : std_logic;
signal \N__40983\ : std_logic;
signal \N__40980\ : std_logic;
signal \N__40979\ : std_logic;
signal \N__40978\ : std_logic;
signal \N__40975\ : std_logic;
signal \N__40972\ : std_logic;
signal \N__40969\ : std_logic;
signal \N__40962\ : std_logic;
signal \N__40959\ : std_logic;
signal \N__40956\ : std_logic;
signal \N__40953\ : std_logic;
signal \N__40950\ : std_logic;
signal \N__40947\ : std_logic;
signal \N__40944\ : std_logic;
signal \N__40943\ : std_logic;
signal \N__40942\ : std_logic;
signal \N__40939\ : std_logic;
signal \N__40934\ : std_logic;
signal \N__40931\ : std_logic;
signal \N__40926\ : std_logic;
signal \N__40923\ : std_logic;
signal \N__40922\ : std_logic;
signal \N__40921\ : std_logic;
signal \N__40918\ : std_logic;
signal \N__40915\ : std_logic;
signal \N__40914\ : std_logic;
signal \N__40911\ : std_logic;
signal \N__40908\ : std_logic;
signal \N__40905\ : std_logic;
signal \N__40902\ : std_logic;
signal \N__40899\ : std_logic;
signal \N__40896\ : std_logic;
signal \N__40893\ : std_logic;
signal \N__40884\ : std_logic;
signal \N__40881\ : std_logic;
signal \N__40878\ : std_logic;
signal \N__40875\ : std_logic;
signal \N__40872\ : std_logic;
signal \N__40869\ : std_logic;
signal \N__40868\ : std_logic;
signal \N__40867\ : std_logic;
signal \N__40866\ : std_logic;
signal \N__40865\ : std_logic;
signal \N__40864\ : std_logic;
signal \N__40861\ : std_logic;
signal \N__40860\ : std_logic;
signal \N__40859\ : std_logic;
signal \N__40858\ : std_logic;
signal \N__40855\ : std_logic;
signal \N__40850\ : std_logic;
signal \N__40845\ : std_logic;
signal \N__40842\ : std_logic;
signal \N__40839\ : std_logic;
signal \N__40838\ : std_logic;
signal \N__40835\ : std_logic;
signal \N__40832\ : std_logic;
signal \N__40831\ : std_logic;
signal \N__40828\ : std_logic;
signal \N__40825\ : std_logic;
signal \N__40820\ : std_logic;
signal \N__40815\ : std_logic;
signal \N__40812\ : std_logic;
signal \N__40807\ : std_logic;
signal \N__40804\ : std_logic;
signal \N__40801\ : std_logic;
signal \N__40798\ : std_logic;
signal \N__40785\ : std_logic;
signal \N__40782\ : std_logic;
signal \N__40779\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40775\ : std_logic;
signal \N__40770\ : std_logic;
signal \N__40767\ : std_logic;
signal \N__40766\ : std_logic;
signal \N__40763\ : std_logic;
signal \N__40760\ : std_logic;
signal \N__40757\ : std_logic;
signal \N__40754\ : std_logic;
signal \N__40751\ : std_logic;
signal \N__40746\ : std_logic;
signal \N__40745\ : std_logic;
signal \N__40742\ : std_logic;
signal \N__40739\ : std_logic;
signal \N__40734\ : std_logic;
signal \N__40733\ : std_logic;
signal \N__40730\ : std_logic;
signal \N__40727\ : std_logic;
signal \N__40726\ : std_logic;
signal \N__40723\ : std_logic;
signal \N__40720\ : std_logic;
signal \N__40717\ : std_logic;
signal \N__40714\ : std_logic;
signal \N__40707\ : std_logic;
signal \N__40704\ : std_logic;
signal \N__40703\ : std_logic;
signal \N__40702\ : std_logic;
signal \N__40699\ : std_logic;
signal \N__40696\ : std_logic;
signal \N__40693\ : std_logic;
signal \N__40692\ : std_logic;
signal \N__40689\ : std_logic;
signal \N__40686\ : std_logic;
signal \N__40681\ : std_logic;
signal \N__40678\ : std_logic;
signal \N__40673\ : std_logic;
signal \N__40668\ : std_logic;
signal \N__40667\ : std_logic;
signal \N__40666\ : std_logic;
signal \N__40661\ : std_logic;
signal \N__40658\ : std_logic;
signal \N__40655\ : std_logic;
signal \N__40652\ : std_logic;
signal \N__40651\ : std_logic;
signal \N__40648\ : std_logic;
signal \N__40645\ : std_logic;
signal \N__40642\ : std_logic;
signal \N__40635\ : std_logic;
signal \N__40632\ : std_logic;
signal \N__40631\ : std_logic;
signal \N__40628\ : std_logic;
signal \N__40625\ : std_logic;
signal \N__40620\ : std_logic;
signal \N__40617\ : std_logic;
signal \N__40616\ : std_logic;
signal \N__40613\ : std_logic;
signal \N__40610\ : std_logic;
signal \N__40605\ : std_logic;
signal \N__40604\ : std_logic;
signal \N__40599\ : std_logic;
signal \N__40596\ : std_logic;
signal \N__40593\ : std_logic;
signal \N__40590\ : std_logic;
signal \N__40587\ : std_logic;
signal \N__40586\ : std_logic;
signal \N__40583\ : std_logic;
signal \N__40580\ : std_logic;
signal \N__40577\ : std_logic;
signal \N__40574\ : std_logic;
signal \N__40569\ : std_logic;
signal \N__40566\ : std_logic;
signal \N__40563\ : std_logic;
signal \N__40560\ : std_logic;
signal \N__40559\ : std_logic;
signal \N__40556\ : std_logic;
signal \N__40553\ : std_logic;
signal \N__40548\ : std_logic;
signal \N__40545\ : std_logic;
signal \N__40542\ : std_logic;
signal \N__40539\ : std_logic;
signal \N__40538\ : std_logic;
signal \N__40533\ : std_logic;
signal \N__40530\ : std_logic;
signal \N__40527\ : std_logic;
signal \N__40524\ : std_logic;
signal \N__40521\ : std_logic;
signal \N__40518\ : std_logic;
signal \N__40515\ : std_logic;
signal \N__40512\ : std_logic;
signal \N__40509\ : std_logic;
signal \N__40506\ : std_logic;
signal \N__40505\ : std_logic;
signal \N__40500\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40494\ : std_logic;
signal \N__40493\ : std_logic;
signal \N__40488\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40481\ : std_logic;
signal \N__40476\ : std_logic;
signal \N__40473\ : std_logic;
signal \N__40470\ : std_logic;
signal \N__40469\ : std_logic;
signal \N__40466\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40458\ : std_logic;
signal \N__40455\ : std_logic;
signal \N__40452\ : std_logic;
signal \N__40449\ : std_logic;
signal \N__40446\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40442\ : std_logic;
signal \N__40439\ : std_logic;
signal \N__40434\ : std_logic;
signal \N__40433\ : std_logic;
signal \N__40430\ : std_logic;
signal \N__40427\ : std_logic;
signal \N__40424\ : std_logic;
signal \N__40419\ : std_logic;
signal \N__40416\ : std_logic;
signal \N__40415\ : std_logic;
signal \N__40414\ : std_logic;
signal \N__40411\ : std_logic;
signal \N__40408\ : std_logic;
signal \N__40405\ : std_logic;
signal \N__40398\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40394\ : std_logic;
signal \N__40391\ : std_logic;
signal \N__40386\ : std_logic;
signal \N__40383\ : std_logic;
signal \N__40380\ : std_logic;
signal \N__40377\ : std_logic;
signal \N__40374\ : std_logic;
signal \N__40371\ : std_logic;
signal \N__40368\ : std_logic;
signal \N__40365\ : std_logic;
signal \N__40362\ : std_logic;
signal \N__40359\ : std_logic;
signal \N__40356\ : std_logic;
signal \N__40353\ : std_logic;
signal \N__40350\ : std_logic;
signal \N__40347\ : std_logic;
signal \N__40344\ : std_logic;
signal \N__40341\ : std_logic;
signal \N__40338\ : std_logic;
signal \N__40335\ : std_logic;
signal \N__40332\ : std_logic;
signal \N__40329\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40320\ : std_logic;
signal \N__40319\ : std_logic;
signal \N__40318\ : std_logic;
signal \N__40315\ : std_logic;
signal \N__40314\ : std_logic;
signal \N__40311\ : std_logic;
signal \N__40308\ : std_logic;
signal \N__40305\ : std_logic;
signal \N__40302\ : std_logic;
signal \N__40297\ : std_logic;
signal \N__40294\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40288\ : std_logic;
signal \N__40285\ : std_logic;
signal \N__40278\ : std_logic;
signal \N__40275\ : std_logic;
signal \N__40272\ : std_logic;
signal \N__40269\ : std_logic;
signal \N__40266\ : std_logic;
signal \N__40263\ : std_logic;
signal \N__40260\ : std_logic;
signal \N__40257\ : std_logic;
signal \N__40256\ : std_logic;
signal \N__40253\ : std_logic;
signal \N__40250\ : std_logic;
signal \N__40245\ : std_logic;
signal \N__40244\ : std_logic;
signal \N__40243\ : std_logic;
signal \N__40240\ : std_logic;
signal \N__40235\ : std_logic;
signal \N__40230\ : std_logic;
signal \N__40227\ : std_logic;
signal \N__40224\ : std_logic;
signal \N__40223\ : std_logic;
signal \N__40222\ : std_logic;
signal \N__40219\ : std_logic;
signal \N__40216\ : std_logic;
signal \N__40213\ : std_logic;
signal \N__40208\ : std_logic;
signal \N__40205\ : std_logic;
signal \N__40204\ : std_logic;
signal \N__40201\ : std_logic;
signal \N__40198\ : std_logic;
signal \N__40195\ : std_logic;
signal \N__40188\ : std_logic;
signal \N__40185\ : std_logic;
signal \N__40182\ : std_logic;
signal \N__40179\ : std_logic;
signal \N__40176\ : std_logic;
signal \N__40173\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40167\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40161\ : std_logic;
signal \N__40158\ : std_logic;
signal \N__40155\ : std_logic;
signal \N__40152\ : std_logic;
signal \N__40149\ : std_logic;
signal \N__40146\ : std_logic;
signal \N__40143\ : std_logic;
signal \N__40140\ : std_logic;
signal \N__40137\ : std_logic;
signal \N__40134\ : std_logic;
signal \N__40131\ : std_logic;
signal \N__40130\ : std_logic;
signal \N__40127\ : std_logic;
signal \N__40124\ : std_logic;
signal \N__40123\ : std_logic;
signal \N__40120\ : std_logic;
signal \N__40117\ : std_logic;
signal \N__40114\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40110\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40104\ : std_logic;
signal \N__40101\ : std_logic;
signal \N__40092\ : std_logic;
signal \N__40089\ : std_logic;
signal \N__40086\ : std_logic;
signal \N__40083\ : std_logic;
signal \N__40080\ : std_logic;
signal \N__40077\ : std_logic;
signal \N__40074\ : std_logic;
signal \N__40073\ : std_logic;
signal \N__40072\ : std_logic;
signal \N__40069\ : std_logic;
signal \N__40066\ : std_logic;
signal \N__40063\ : std_logic;
signal \N__40062\ : std_logic;
signal \N__40059\ : std_logic;
signal \N__40056\ : std_logic;
signal \N__40053\ : std_logic;
signal \N__40050\ : std_logic;
signal \N__40049\ : std_logic;
signal \N__40046\ : std_logic;
signal \N__40043\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40035\ : std_logic;
signal \N__40030\ : std_logic;
signal \N__40027\ : std_logic;
signal \N__40024\ : std_logic;
signal \N__40017\ : std_logic;
signal \N__40014\ : std_logic;
signal \N__40011\ : std_logic;
signal \N__40008\ : std_logic;
signal \N__40005\ : std_logic;
signal \N__40002\ : std_logic;
signal \N__39999\ : std_logic;
signal \N__39996\ : std_logic;
signal \N__39993\ : std_logic;
signal \N__39990\ : std_logic;
signal \N__39987\ : std_logic;
signal \N__39984\ : std_logic;
signal \N__39981\ : std_logic;
signal \N__39980\ : std_logic;
signal \N__39977\ : std_logic;
signal \N__39974\ : std_logic;
signal \N__39973\ : std_logic;
signal \N__39968\ : std_logic;
signal \N__39965\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39954\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39948\ : std_logic;
signal \N__39947\ : std_logic;
signal \N__39942\ : std_logic;
signal \N__39941\ : std_logic;
signal \N__39940\ : std_logic;
signal \N__39937\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39927\ : std_logic;
signal \N__39924\ : std_logic;
signal \N__39921\ : std_logic;
signal \N__39918\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39912\ : std_logic;
signal \N__39909\ : std_logic;
signal \N__39906\ : std_logic;
signal \N__39903\ : std_logic;
signal \N__39900\ : std_logic;
signal \N__39897\ : std_logic;
signal \N__39894\ : std_logic;
signal \N__39891\ : std_logic;
signal \N__39888\ : std_logic;
signal \N__39885\ : std_logic;
signal \N__39882\ : std_logic;
signal \N__39879\ : std_logic;
signal \N__39876\ : std_logic;
signal \N__39873\ : std_logic;
signal \N__39870\ : std_logic;
signal \N__39867\ : std_logic;
signal \N__39864\ : std_logic;
signal \N__39863\ : std_logic;
signal \N__39860\ : std_logic;
signal \N__39859\ : std_logic;
signal \N__39852\ : std_logic;
signal \N__39851\ : std_logic;
signal \N__39848\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39840\ : std_logic;
signal \N__39837\ : std_logic;
signal \N__39834\ : std_logic;
signal \N__39831\ : std_logic;
signal \N__39828\ : std_logic;
signal \N__39825\ : std_logic;
signal \N__39822\ : std_logic;
signal \N__39819\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39813\ : std_logic;
signal \N__39810\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39806\ : std_logic;
signal \N__39803\ : std_logic;
signal \N__39802\ : std_logic;
signal \N__39795\ : std_logic;
signal \N__39792\ : std_logic;
signal \N__39791\ : std_logic;
signal \N__39788\ : std_logic;
signal \N__39785\ : std_logic;
signal \N__39780\ : std_logic;
signal \N__39777\ : std_logic;
signal \N__39774\ : std_logic;
signal \N__39771\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39762\ : std_logic;
signal \N__39759\ : std_logic;
signal \N__39756\ : std_logic;
signal \N__39753\ : std_logic;
signal \N__39750\ : std_logic;
signal \N__39747\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39741\ : std_logic;
signal \N__39738\ : std_logic;
signal \N__39735\ : std_logic;
signal \N__39732\ : std_logic;
signal \N__39729\ : std_logic;
signal \N__39726\ : std_logic;
signal \N__39723\ : std_logic;
signal \N__39720\ : std_logic;
signal \N__39717\ : std_logic;
signal \N__39714\ : std_logic;
signal \N__39711\ : std_logic;
signal \N__39708\ : std_logic;
signal \N__39705\ : std_logic;
signal \N__39702\ : std_logic;
signal \N__39699\ : std_logic;
signal \N__39696\ : std_logic;
signal \N__39693\ : std_logic;
signal \N__39690\ : std_logic;
signal \N__39687\ : std_logic;
signal \N__39684\ : std_logic;
signal \N__39683\ : std_logic;
signal \N__39682\ : std_logic;
signal \N__39681\ : std_logic;
signal \N__39678\ : std_logic;
signal \N__39673\ : std_logic;
signal \N__39668\ : std_logic;
signal \N__39665\ : std_logic;
signal \N__39662\ : std_logic;
signal \N__39659\ : std_logic;
signal \N__39654\ : std_logic;
signal \N__39651\ : std_logic;
signal \N__39648\ : std_logic;
signal \N__39645\ : std_logic;
signal \N__39642\ : std_logic;
signal \N__39639\ : std_logic;
signal \N__39636\ : std_logic;
signal \N__39633\ : std_logic;
signal \N__39630\ : std_logic;
signal \N__39627\ : std_logic;
signal \N__39624\ : std_logic;
signal \N__39621\ : std_logic;
signal \N__39618\ : std_logic;
signal \N__39615\ : std_logic;
signal \N__39612\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39608\ : std_logic;
signal \N__39605\ : std_logic;
signal \N__39600\ : std_logic;
signal \N__39599\ : std_logic;
signal \N__39596\ : std_logic;
signal \N__39593\ : std_logic;
signal \N__39588\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39582\ : std_logic;
signal \N__39579\ : std_logic;
signal \N__39578\ : std_logic;
signal \N__39577\ : std_logic;
signal \N__39574\ : std_logic;
signal \N__39571\ : std_logic;
signal \N__39568\ : std_logic;
signal \N__39561\ : std_logic;
signal \N__39560\ : std_logic;
signal \N__39559\ : std_logic;
signal \N__39556\ : std_logic;
signal \N__39553\ : std_logic;
signal \N__39550\ : std_logic;
signal \N__39543\ : std_logic;
signal \N__39540\ : std_logic;
signal \N__39537\ : std_logic;
signal \N__39534\ : std_logic;
signal \N__39531\ : std_logic;
signal \N__39528\ : std_logic;
signal \N__39525\ : std_logic;
signal \N__39524\ : std_logic;
signal \N__39523\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39515\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39511\ : std_logic;
signal \N__39508\ : std_logic;
signal \N__39505\ : std_logic;
signal \N__39498\ : std_logic;
signal \N__39495\ : std_logic;
signal \N__39492\ : std_logic;
signal \N__39489\ : std_logic;
signal \N__39486\ : std_logic;
signal \N__39483\ : std_logic;
signal \N__39480\ : std_logic;
signal \N__39477\ : std_logic;
signal \N__39474\ : std_logic;
signal \N__39471\ : std_logic;
signal \N__39468\ : std_logic;
signal \N__39465\ : std_logic;
signal \N__39462\ : std_logic;
signal \N__39459\ : std_logic;
signal \N__39456\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39446\ : std_logic;
signal \N__39443\ : std_logic;
signal \N__39440\ : std_logic;
signal \N__39435\ : std_logic;
signal \N__39432\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39425\ : std_logic;
signal \N__39424\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39416\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39408\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39406\ : std_logic;
signal \N__39403\ : std_logic;
signal \N__39398\ : std_logic;
signal \N__39393\ : std_logic;
signal \N__39390\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39384\ : std_logic;
signal \N__39381\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39375\ : std_logic;
signal \N__39374\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39366\ : std_logic;
signal \N__39363\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39359\ : std_logic;
signal \N__39358\ : std_logic;
signal \N__39355\ : std_logic;
signal \N__39354\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39348\ : std_logic;
signal \N__39345\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39339\ : std_logic;
signal \N__39330\ : std_logic;
signal \N__39327\ : std_logic;
signal \N__39324\ : std_logic;
signal \N__39323\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39319\ : std_logic;
signal \N__39316\ : std_logic;
signal \N__39313\ : std_logic;
signal \N__39310\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39300\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39294\ : std_logic;
signal \N__39291\ : std_logic;
signal \N__39290\ : std_logic;
signal \N__39287\ : std_logic;
signal \N__39284\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39278\ : std_logic;
signal \N__39275\ : std_logic;
signal \N__39272\ : std_logic;
signal \N__39267\ : std_logic;
signal \N__39264\ : std_logic;
signal \N__39261\ : std_logic;
signal \N__39258\ : std_logic;
signal \N__39255\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39249\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39245\ : std_logic;
signal \N__39242\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39234\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39222\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39215\ : std_logic;
signal \N__39212\ : std_logic;
signal \N__39209\ : std_logic;
signal \N__39204\ : std_logic;
signal \N__39201\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39186\ : std_logic;
signal \N__39183\ : std_logic;
signal \N__39180\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39171\ : std_logic;
signal \N__39168\ : std_logic;
signal \N__39167\ : std_logic;
signal \N__39164\ : std_logic;
signal \N__39161\ : std_logic;
signal \N__39158\ : std_logic;
signal \N__39153\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39141\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39131\ : std_logic;
signal \N__39128\ : std_logic;
signal \N__39123\ : std_logic;
signal \N__39120\ : std_logic;
signal \N__39117\ : std_logic;
signal \N__39116\ : std_logic;
signal \N__39113\ : std_logic;
signal \N__39110\ : std_logic;
signal \N__39105\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39099\ : std_logic;
signal \N__39096\ : std_logic;
signal \N__39093\ : std_logic;
signal \N__39090\ : std_logic;
signal \N__39089\ : std_logic;
signal \N__39086\ : std_logic;
signal \N__39083\ : std_logic;
signal \N__39078\ : std_logic;
signal \N__39075\ : std_logic;
signal \N__39072\ : std_logic;
signal \N__39069\ : std_logic;
signal \N__39068\ : std_logic;
signal \N__39065\ : std_logic;
signal \N__39062\ : std_logic;
signal \N__39057\ : std_logic;
signal \N__39054\ : std_logic;
signal \N__39051\ : std_logic;
signal \N__39048\ : std_logic;
signal \N__39045\ : std_logic;
signal \N__39042\ : std_logic;
signal \N__39039\ : std_logic;
signal \N__39036\ : std_logic;
signal \N__39033\ : std_logic;
signal \N__39030\ : std_logic;
signal \N__39027\ : std_logic;
signal \N__39024\ : std_logic;
signal \N__39021\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39014\ : std_logic;
signal \N__39009\ : std_logic;
signal \N__39006\ : std_logic;
signal \N__39003\ : std_logic;
signal \N__39000\ : std_logic;
signal \N__38999\ : std_logic;
signal \N__38996\ : std_logic;
signal \N__38993\ : std_logic;
signal \N__38988\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38982\ : std_logic;
signal \N__38979\ : std_logic;
signal \N__38978\ : std_logic;
signal \N__38975\ : std_logic;
signal \N__38972\ : std_logic;
signal \N__38967\ : std_logic;
signal \N__38964\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38958\ : std_logic;
signal \N__38957\ : std_logic;
signal \N__38954\ : std_logic;
signal \N__38951\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38947\ : std_logic;
signal \N__38944\ : std_logic;
signal \N__38941\ : std_logic;
signal \N__38938\ : std_logic;
signal \N__38931\ : std_logic;
signal \N__38928\ : std_logic;
signal \N__38925\ : std_logic;
signal \N__38922\ : std_logic;
signal \N__38921\ : std_logic;
signal \N__38918\ : std_logic;
signal \N__38915\ : std_logic;
signal \N__38910\ : std_logic;
signal \N__38907\ : std_logic;
signal \N__38904\ : std_logic;
signal \N__38901\ : std_logic;
signal \N__38900\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38894\ : std_logic;
signal \N__38889\ : std_logic;
signal \N__38886\ : std_logic;
signal \N__38883\ : std_logic;
signal \N__38880\ : std_logic;
signal \N__38879\ : std_logic;
signal \N__38876\ : std_logic;
signal \N__38873\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38865\ : std_logic;
signal \N__38862\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38858\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38852\ : std_logic;
signal \N__38847\ : std_logic;
signal \N__38844\ : std_logic;
signal \N__38841\ : std_logic;
signal \N__38838\ : std_logic;
signal \N__38835\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38823\ : std_logic;
signal \N__38820\ : std_logic;
signal \N__38817\ : std_logic;
signal \N__38814\ : std_logic;
signal \N__38813\ : std_logic;
signal \N__38812\ : std_logic;
signal \N__38807\ : std_logic;
signal \N__38804\ : std_logic;
signal \N__38801\ : std_logic;
signal \N__38796\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38792\ : std_logic;
signal \N__38787\ : std_logic;
signal \N__38784\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38782\ : std_logic;
signal \N__38779\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38769\ : std_logic;
signal \N__38766\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38757\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38739\ : std_logic;
signal \N__38736\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38727\ : std_logic;
signal \N__38724\ : std_logic;
signal \N__38721\ : std_logic;
signal \N__38718\ : std_logic;
signal \N__38715\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38709\ : std_logic;
signal \N__38706\ : std_logic;
signal \N__38703\ : std_logic;
signal \N__38700\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38691\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38672\ : std_logic;
signal \N__38669\ : std_logic;
signal \N__38666\ : std_logic;
signal \N__38661\ : std_logic;
signal \N__38660\ : std_logic;
signal \N__38659\ : std_logic;
signal \N__38656\ : std_logic;
signal \N__38653\ : std_logic;
signal \N__38648\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38642\ : std_logic;
signal \N__38641\ : std_logic;
signal \N__38638\ : std_logic;
signal \N__38635\ : std_logic;
signal \N__38632\ : std_logic;
signal \N__38625\ : std_logic;
signal \N__38622\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38610\ : std_logic;
signal \N__38609\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38601\ : std_logic;
signal \N__38598\ : std_logic;
signal \N__38595\ : std_logic;
signal \N__38592\ : std_logic;
signal \N__38589\ : std_logic;
signal \N__38586\ : std_logic;
signal \N__38583\ : std_logic;
signal \N__38580\ : std_logic;
signal \N__38577\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38562\ : std_logic;
signal \N__38559\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38547\ : std_logic;
signal \N__38544\ : std_logic;
signal \N__38541\ : std_logic;
signal \N__38538\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38529\ : std_logic;
signal \N__38528\ : std_logic;
signal \N__38525\ : std_logic;
signal \N__38522\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38520\ : std_logic;
signal \N__38519\ : std_logic;
signal \N__38518\ : std_logic;
signal \N__38515\ : std_logic;
signal \N__38514\ : std_logic;
signal \N__38513\ : std_logic;
signal \N__38512\ : std_logic;
signal \N__38509\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38499\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38496\ : std_logic;
signal \N__38495\ : std_logic;
signal \N__38494\ : std_logic;
signal \N__38491\ : std_logic;
signal \N__38484\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38468\ : std_logic;
signal \N__38465\ : std_logic;
signal \N__38454\ : std_logic;
signal \N__38451\ : std_logic;
signal \N__38448\ : std_logic;
signal \N__38445\ : std_logic;
signal \N__38442\ : std_logic;
signal \N__38439\ : std_logic;
signal \N__38436\ : std_logic;
signal \N__38433\ : std_logic;
signal \N__38430\ : std_logic;
signal \N__38427\ : std_logic;
signal \N__38424\ : std_logic;
signal \N__38421\ : std_logic;
signal \N__38418\ : std_logic;
signal \N__38415\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38409\ : std_logic;
signal \N__38406\ : std_logic;
signal \N__38403\ : std_logic;
signal \N__38400\ : std_logic;
signal \N__38397\ : std_logic;
signal \N__38394\ : std_logic;
signal \N__38391\ : std_logic;
signal \N__38388\ : std_logic;
signal \N__38385\ : std_logic;
signal \N__38382\ : std_logic;
signal \N__38379\ : std_logic;
signal \N__38376\ : std_logic;
signal \N__38373\ : std_logic;
signal \N__38370\ : std_logic;
signal \N__38367\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38361\ : std_logic;
signal \N__38358\ : std_logic;
signal \N__38355\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38349\ : std_logic;
signal \N__38346\ : std_logic;
signal \N__38343\ : std_logic;
signal \N__38340\ : std_logic;
signal \N__38337\ : std_logic;
signal \N__38334\ : std_logic;
signal \N__38331\ : std_logic;
signal \N__38328\ : std_logic;
signal \N__38325\ : std_logic;
signal \N__38322\ : std_logic;
signal \N__38319\ : std_logic;
signal \N__38316\ : std_logic;
signal \N__38313\ : std_logic;
signal \N__38310\ : std_logic;
signal \N__38307\ : std_logic;
signal \N__38304\ : std_logic;
signal \N__38301\ : std_logic;
signal \N__38298\ : std_logic;
signal \N__38295\ : std_logic;
signal \N__38292\ : std_logic;
signal \N__38289\ : std_logic;
signal \N__38286\ : std_logic;
signal \N__38283\ : std_logic;
signal \N__38282\ : std_logic;
signal \N__38281\ : std_logic;
signal \N__38280\ : std_logic;
signal \N__38279\ : std_logic;
signal \N__38278\ : std_logic;
signal \N__38277\ : std_logic;
signal \N__38276\ : std_logic;
signal \N__38275\ : std_logic;
signal \N__38274\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38270\ : std_logic;
signal \N__38267\ : std_logic;
signal \N__38260\ : std_logic;
signal \N__38251\ : std_logic;
signal \N__38250\ : std_logic;
signal \N__38249\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38247\ : std_logic;
signal \N__38246\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38244\ : std_logic;
signal \N__38243\ : std_logic;
signal \N__38240\ : std_logic;
signal \N__38237\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38226\ : std_logic;
signal \N__38223\ : std_logic;
signal \N__38216\ : std_logic;
signal \N__38207\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38200\ : std_logic;
signal \N__38199\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38194\ : std_logic;
signal \N__38193\ : std_logic;
signal \N__38192\ : std_logic;
signal \N__38189\ : std_logic;
signal \N__38180\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38172\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38162\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38158\ : std_logic;
signal \N__38157\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38153\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38149\ : std_logic;
signal \N__38148\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38146\ : std_logic;
signal \N__38145\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38143\ : std_logic;
signal \N__38142\ : std_logic;
signal \N__38141\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38139\ : std_logic;
signal \N__38138\ : std_logic;
signal \N__38135\ : std_logic;
signal \N__38132\ : std_logic;
signal \N__38125\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38117\ : std_logic;
signal \N__38102\ : std_logic;
signal \N__38099\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38094\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38090\ : std_logic;
signal \N__38087\ : std_logic;
signal \N__38086\ : std_logic;
signal \N__38083\ : std_logic;
signal \N__38082\ : std_logic;
signal \N__38079\ : std_logic;
signal \N__38078\ : std_logic;
signal \N__38075\ : std_logic;
signal \N__38074\ : std_logic;
signal \N__38071\ : std_logic;
signal \N__38070\ : std_logic;
signal \N__38069\ : std_logic;
signal \N__38066\ : std_logic;
signal \N__38065\ : std_logic;
signal \N__38062\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38058\ : std_logic;
signal \N__38057\ : std_logic;
signal \N__38054\ : std_logic;
signal \N__38051\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38043\ : std_logic;
signal \N__38040\ : std_logic;
signal \N__38023\ : std_logic;
signal \N__38006\ : std_logic;
signal \N__37991\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37981\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37965\ : std_logic;
signal \N__37962\ : std_logic;
signal \N__37959\ : std_logic;
signal \N__37956\ : std_logic;
signal \N__37953\ : std_logic;
signal \N__37950\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37944\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37926\ : std_logic;
signal \N__37923\ : std_logic;
signal \N__37922\ : std_logic;
signal \N__37919\ : std_logic;
signal \N__37916\ : std_logic;
signal \N__37915\ : std_logic;
signal \N__37910\ : std_logic;
signal \N__37907\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37896\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37892\ : std_logic;
signal \N__37891\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37882\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37877\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37869\ : std_logic;
signal \N__37866\ : std_logic;
signal \N__37863\ : std_logic;
signal \N__37860\ : std_logic;
signal \N__37855\ : std_logic;
signal \N__37848\ : std_logic;
signal \N__37845\ : std_logic;
signal \N__37842\ : std_logic;
signal \N__37839\ : std_logic;
signal \N__37836\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37829\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37821\ : std_logic;
signal \N__37818\ : std_logic;
signal \N__37817\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37811\ : std_logic;
signal \N__37808\ : std_logic;
signal \N__37803\ : std_logic;
signal \N__37800\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37788\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37782\ : std_logic;
signal \N__37779\ : std_logic;
signal \N__37776\ : std_logic;
signal \N__37773\ : std_logic;
signal \N__37770\ : std_logic;
signal \N__37767\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37755\ : std_logic;
signal \N__37752\ : std_logic;
signal \N__37751\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37745\ : std_logic;
signal \N__37740\ : std_logic;
signal \N__37737\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37733\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37727\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37719\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37712\ : std_logic;
signal \N__37709\ : std_logic;
signal \N__37706\ : std_logic;
signal \N__37701\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37695\ : std_logic;
signal \N__37692\ : std_logic;
signal \N__37689\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37680\ : std_logic;
signal \N__37677\ : std_logic;
signal \N__37674\ : std_logic;
signal \N__37671\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37662\ : std_logic;
signal \N__37659\ : std_logic;
signal \N__37656\ : std_logic;
signal \N__37655\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37652\ : std_logic;
signal \N__37649\ : std_logic;
signal \N__37644\ : std_logic;
signal \N__37639\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37631\ : std_logic;
signal \N__37630\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37625\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37608\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37587\ : std_logic;
signal \N__37584\ : std_logic;
signal \N__37581\ : std_logic;
signal \N__37578\ : std_logic;
signal \N__37575\ : std_logic;
signal \N__37572\ : std_logic;
signal \N__37569\ : std_logic;
signal \N__37566\ : std_logic;
signal \N__37563\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37553\ : std_logic;
signal \N__37550\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37546\ : std_logic;
signal \N__37545\ : std_logic;
signal \N__37540\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37532\ : std_logic;
signal \N__37527\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37507\ : std_logic;
signal \N__37504\ : std_logic;
signal \N__37501\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37491\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37485\ : std_logic;
signal \N__37484\ : std_logic;
signal \N__37483\ : std_logic;
signal \N__37482\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37473\ : std_logic;
signal \N__37470\ : std_logic;
signal \N__37467\ : std_logic;
signal \N__37458\ : std_logic;
signal \N__37457\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37453\ : std_logic;
signal \N__37450\ : std_logic;
signal \N__37447\ : std_logic;
signal \N__37444\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37421\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37401\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37392\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37386\ : std_logic;
signal \N__37383\ : std_logic;
signal \N__37380\ : std_logic;
signal \N__37377\ : std_logic;
signal \N__37374\ : std_logic;
signal \N__37371\ : std_logic;
signal \N__37368\ : std_logic;
signal \N__37365\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37359\ : std_logic;
signal \N__37356\ : std_logic;
signal \N__37355\ : std_logic;
signal \N__37352\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37338\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37320\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37314\ : std_logic;
signal \N__37311\ : std_logic;
signal \N__37308\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37263\ : std_logic;
signal \N__37260\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37253\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37245\ : std_logic;
signal \N__37242\ : std_logic;
signal \N__37239\ : std_logic;
signal \N__37236\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37229\ : std_logic;
signal \N__37226\ : std_logic;
signal \N__37221\ : std_logic;
signal \N__37218\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37208\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37199\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37185\ : std_logic;
signal \N__37182\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37175\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37167\ : std_logic;
signal \N__37164\ : std_logic;
signal \N__37161\ : std_logic;
signal \N__37158\ : std_logic;
signal \N__37155\ : std_logic;
signal \N__37152\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37137\ : std_logic;
signal \N__37134\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37104\ : std_logic;
signal \N__37101\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37094\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37086\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37073\ : std_logic;
signal \N__37068\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37058\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37050\ : std_logic;
signal \N__37047\ : std_logic;
signal \N__37046\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37032\ : std_logic;
signal \N__37029\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37025\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37014\ : std_logic;
signal \N__37011\ : std_logic;
signal \N__37008\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36975\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36962\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36933\ : std_logic;
signal \N__36930\ : std_logic;
signal \N__36927\ : std_logic;
signal \N__36924\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36915\ : std_logic;
signal \N__36914\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36907\ : std_logic;
signal \N__36904\ : std_logic;
signal \N__36897\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36891\ : std_logic;
signal \N__36888\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36870\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36860\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36851\ : std_logic;
signal \N__36846\ : std_logic;
signal \N__36843\ : std_logic;
signal \N__36840\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36836\ : std_logic;
signal \N__36833\ : std_logic;
signal \N__36830\ : std_logic;
signal \N__36827\ : std_logic;
signal \N__36824\ : std_logic;
signal \N__36821\ : std_logic;
signal \N__36818\ : std_logic;
signal \N__36813\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36798\ : std_logic;
signal \N__36795\ : std_logic;
signal \N__36792\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36787\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36778\ : std_logic;
signal \N__36775\ : std_logic;
signal \N__36768\ : std_logic;
signal \N__36765\ : std_logic;
signal \N__36762\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36756\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36747\ : std_logic;
signal \N__36744\ : std_logic;
signal \N__36741\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36730\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36714\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36709\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36683\ : std_logic;
signal \N__36680\ : std_logic;
signal \N__36675\ : std_logic;
signal \N__36672\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36669\ : std_logic;
signal \N__36668\ : std_logic;
signal \N__36667\ : std_logic;
signal \N__36666\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36658\ : std_logic;
signal \N__36657\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36654\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36652\ : std_logic;
signal \N__36651\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36648\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36637\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36634\ : std_logic;
signal \N__36633\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36631\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36578\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36539\ : std_logic;
signal \N__36536\ : std_logic;
signal \N__36533\ : std_logic;
signal \N__36528\ : std_logic;
signal \N__36525\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36523\ : std_logic;
signal \N__36520\ : std_logic;
signal \N__36517\ : std_logic;
signal \N__36516\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36508\ : std_logic;
signal \N__36505\ : std_logic;
signal \N__36502\ : std_logic;
signal \N__36497\ : std_logic;
signal \N__36494\ : std_logic;
signal \N__36489\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36480\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36474\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36466\ : std_logic;
signal \N__36463\ : std_logic;
signal \N__36460\ : std_logic;
signal \N__36453\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36449\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36443\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36425\ : std_logic;
signal \N__36424\ : std_logic;
signal \N__36419\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36408\ : std_logic;
signal \N__36405\ : std_logic;
signal \N__36404\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36398\ : std_logic;
signal \N__36393\ : std_logic;
signal \N__36392\ : std_logic;
signal \N__36389\ : std_logic;
signal \N__36386\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36378\ : std_logic;
signal \N__36375\ : std_logic;
signal \N__36374\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36351\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36347\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36330\ : std_logic;
signal \N__36327\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36323\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36313\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36305\ : std_logic;
signal \N__36300\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36292\ : std_logic;
signal \N__36289\ : std_logic;
signal \N__36286\ : std_logic;
signal \N__36283\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36267\ : std_logic;
signal \N__36264\ : std_logic;
signal \N__36261\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36240\ : std_logic;
signal \N__36237\ : std_logic;
signal \N__36234\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36226\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36220\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36210\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36186\ : std_logic;
signal \N__36183\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36176\ : std_logic;
signal \N__36173\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36162\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36150\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36135\ : std_logic;
signal \N__36132\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36128\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36119\ : std_logic;
signal \N__36116\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36105\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36103\ : std_logic;
signal \N__36098\ : std_logic;
signal \N__36095\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36087\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36051\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36043\ : std_logic;
signal \N__36040\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36017\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36008\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__35997\ : std_logic;
signal \N__35994\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35987\ : std_logic;
signal \N__35986\ : std_logic;
signal \N__35983\ : std_logic;
signal \N__35980\ : std_logic;
signal \N__35977\ : std_logic;
signal \N__35974\ : std_logic;
signal \N__35971\ : std_logic;
signal \N__35964\ : std_logic;
signal \N__35961\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35959\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35948\ : std_logic;
signal \N__35943\ : std_logic;
signal \N__35940\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35932\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35921\ : std_logic;
signal \N__35916\ : std_logic;
signal \N__35913\ : std_logic;
signal \N__35912\ : std_logic;
signal \N__35909\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35901\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35879\ : std_logic;
signal \N__35876\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35866\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35856\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35850\ : std_logic;
signal \N__35849\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35845\ : std_logic;
signal \N__35842\ : std_logic;
signal \N__35839\ : std_logic;
signal \N__35836\ : std_logic;
signal \N__35829\ : std_logic;
signal \N__35826\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35807\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35801\ : std_logic;
signal \N__35800\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35794\ : std_logic;
signal \N__35791\ : std_logic;
signal \N__35784\ : std_logic;
signal \N__35781\ : std_logic;
signal \N__35780\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35770\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35764\ : std_logic;
signal \N__35757\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35751\ : std_logic;
signal \N__35750\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35740\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35727\ : std_logic;
signal \N__35724\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35700\ : std_logic;
signal \N__35697\ : std_logic;
signal \N__35694\ : std_logic;
signal \N__35691\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35687\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35679\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35673\ : std_logic;
signal \N__35670\ : std_logic;
signal \N__35669\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35665\ : std_logic;
signal \N__35662\ : std_logic;
signal \N__35659\ : std_logic;
signal \N__35652\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35650\ : std_logic;
signal \N__35649\ : std_logic;
signal \N__35646\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35639\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35625\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35592\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35557\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35505\ : std_logic;
signal \N__35502\ : std_logic;
signal \N__35499\ : std_logic;
signal \N__35496\ : std_logic;
signal \N__35493\ : std_logic;
signal \N__35490\ : std_logic;
signal \N__35487\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35475\ : std_logic;
signal \N__35474\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35463\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35457\ : std_logic;
signal \N__35454\ : std_logic;
signal \N__35451\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35412\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35397\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35355\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35352\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35331\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35313\ : std_logic;
signal \N__35310\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35286\ : std_logic;
signal \N__35283\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35253\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35247\ : std_logic;
signal \N__35244\ : std_logic;
signal \N__35241\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35229\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35217\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35205\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35193\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35172\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35163\ : std_logic;
signal \N__35158\ : std_logic;
signal \N__35155\ : std_logic;
signal \N__35152\ : std_logic;
signal \N__35149\ : std_logic;
signal \N__35142\ : std_logic;
signal \N__35139\ : std_logic;
signal \N__35138\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35118\ : std_logic;
signal \N__35115\ : std_logic;
signal \N__35112\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35106\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35067\ : std_logic;
signal \N__35064\ : std_logic;
signal \N__35061\ : std_logic;
signal \N__35058\ : std_logic;
signal \N__35055\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35049\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35043\ : std_logic;
signal \N__35040\ : std_logic;
signal \N__35037\ : std_logic;
signal \N__35034\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35028\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35022\ : std_logic;
signal \N__35019\ : std_logic;
signal \N__35016\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35010\ : std_logic;
signal \N__35007\ : std_logic;
signal \N__35004\ : std_logic;
signal \N__35001\ : std_logic;
signal \N__34998\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34992\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34985\ : std_logic;
signal \N__34984\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34970\ : std_logic;
signal \N__34965\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34954\ : std_logic;
signal \N__34951\ : std_logic;
signal \N__34948\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34918\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34904\ : std_logic;
signal \N__34899\ : std_logic;
signal \N__34898\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34890\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34876\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34824\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34818\ : std_logic;
signal \N__34815\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34791\ : std_logic;
signal \N__34790\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34779\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34770\ : std_logic;
signal \N__34767\ : std_logic;
signal \N__34764\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34749\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34713\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34689\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34671\ : std_logic;
signal \N__34668\ : std_logic;
signal \N__34665\ : std_logic;
signal \N__34662\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34656\ : std_logic;
signal \N__34653\ : std_logic;
signal \N__34650\ : std_logic;
signal \N__34647\ : std_logic;
signal \N__34644\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34629\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34623\ : std_logic;
signal \N__34620\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34599\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34559\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34554\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34531\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34510\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34507\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34492\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34477\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34465\ : std_logic;
signal \N__34460\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34438\ : std_logic;
signal \N__34435\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34407\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34391\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34378\ : std_logic;
signal \N__34375\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34365\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34361\ : std_logic;
signal \N__34358\ : std_logic;
signal \N__34357\ : std_logic;
signal \N__34354\ : std_logic;
signal \N__34351\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34341\ : std_logic;
signal \N__34338\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34316\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34310\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34299\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34287\ : std_logic;
signal \N__34278\ : std_logic;
signal \N__34275\ : std_logic;
signal \N__34272\ : std_logic;
signal \N__34269\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34254\ : std_logic;
signal \N__34253\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34240\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34232\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34218\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34213\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34204\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34185\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34179\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34172\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34151\ : std_logic;
signal \N__34148\ : std_logic;
signal \N__34145\ : std_logic;
signal \N__34140\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34118\ : std_logic;
signal \N__34115\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34100\ : std_logic;
signal \N__34097\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34068\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34022\ : std_logic;
signal \N__34019\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33995\ : std_logic;
signal \N__33992\ : std_logic;
signal \N__33989\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33978\ : std_logic;
signal \N__33975\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33957\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33900\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33890\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33879\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33843\ : std_logic;
signal \N__33840\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33834\ : std_logic;
signal \N__33831\ : std_logic;
signal \N__33828\ : std_logic;
signal \N__33825\ : std_logic;
signal \N__33822\ : std_logic;
signal \N__33819\ : std_logic;
signal \N__33816\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33810\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33801\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33795\ : std_logic;
signal \N__33792\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33756\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33729\ : std_logic;
signal \N__33726\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33720\ : std_logic;
signal \N__33717\ : std_logic;
signal \N__33714\ : std_logic;
signal \N__33711\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33705\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33690\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33684\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33672\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33660\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33654\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33624\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33618\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33591\ : std_logic;
signal \N__33588\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33579\ : std_logic;
signal \N__33576\ : std_logic;
signal \N__33573\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33567\ : std_logic;
signal \N__33564\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33552\ : std_logic;
signal \N__33549\ : std_logic;
signal \N__33546\ : std_logic;
signal \N__33543\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33528\ : std_logic;
signal \N__33525\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33498\ : std_logic;
signal \N__33495\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33486\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33480\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33462\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33431\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33425\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33399\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33351\ : std_logic;
signal \N__33348\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33327\ : std_logic;
signal \N__33324\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33309\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33306\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33283\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33239\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33230\ : std_logic;
signal \N__33229\ : std_logic;
signal \N__33228\ : std_logic;
signal \N__33227\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33216\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33190\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33119\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33107\ : std_logic;
signal \N__33104\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33036\ : std_logic;
signal \N__33035\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33026\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__33003\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32998\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32968\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32930\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32913\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32907\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32890\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32845\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32841\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32803\ : std_logic;
signal \N__32794\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32766\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32758\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32743\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32685\ : std_logic;
signal \N__32682\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32654\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32574\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32557\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32544\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32540\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32536\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32520\ : std_logic;
signal \N__32517\ : std_logic;
signal \N__32514\ : std_logic;
signal \N__32511\ : std_logic;
signal \N__32508\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32487\ : std_logic;
signal \N__32486\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32480\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32388\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32344\ : std_logic;
signal \N__32341\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32326\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32295\ : std_logic;
signal \N__32292\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32271\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32233\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32144\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32124\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32118\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32061\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32028\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31962\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31930\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31899\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31893\ : std_logic;
signal \N__31890\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31875\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31860\ : std_logic;
signal \N__31857\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31844\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31821\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31813\ : std_logic;
signal \N__31810\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31742\ : std_logic;
signal \N__31739\ : std_logic;
signal \N__31736\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31717\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31708\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31676\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31650\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31644\ : std_logic;
signal \N__31641\ : std_logic;
signal \N__31638\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31620\ : std_logic;
signal \N__31617\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31613\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31567\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31558\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31531\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31504\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31495\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31490\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31467\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31438\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31399\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31396\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31382\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31371\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31318\ : std_logic;
signal \N__31305\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31292\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31247\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31235\ : std_logic;
signal \N__31232\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31213\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31184\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31172\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31099\ : std_logic;
signal \N__31094\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31081\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31063\ : std_logic;
signal \N__31058\ : std_logic;
signal \N__31057\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31055\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31036\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31019\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30977\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30949\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30906\ : std_logic;
signal \N__30903\ : std_logic;
signal \N__30900\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30866\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30831\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30822\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30803\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30678\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30674\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30672\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30667\ : std_logic;
signal \N__30666\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30663\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30641\ : std_logic;
signal \N__30634\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30604\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30566\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30545\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30539\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30513\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30483\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30464\ : std_logic;
signal \N__30461\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30408\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30363\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30351\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30333\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30253\ : std_logic;
signal \N__30252\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30242\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30216\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30183\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30155\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30087\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30079\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30063\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30009\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29950\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29925\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29904\ : std_logic;
signal \N__29901\ : std_logic;
signal \N__29898\ : std_logic;
signal \N__29895\ : std_logic;
signal \N__29892\ : std_logic;
signal \N__29889\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29854\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29798\ : std_logic;
signal \N__29795\ : std_logic;
signal \N__29792\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29776\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29751\ : std_logic;
signal \N__29748\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29697\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29687\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29670\ : std_logic;
signal \N__29667\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29429\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29373\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29343\ : std_logic;
signal \N__29340\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29184\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29169\ : std_logic;
signal \N__29166\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29157\ : std_logic;
signal \N__29154\ : std_logic;
signal \N__29151\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29145\ : std_logic;
signal \N__29142\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29094\ : std_logic;
signal \N__29091\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29064\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29058\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29024\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29013\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28883\ : std_logic;
signal \N__28880\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28869\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28860\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28793\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28710\ : std_logic;
signal \N__28709\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28688\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28671\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28644\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28634\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28620\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28565\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28538\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28526\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28496\ : std_logic;
signal \N__28491\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28460\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28448\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28424\ : std_logic;
signal \N__28421\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28400\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28380\ : std_logic;
signal \N__28377\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28370\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28239\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28232\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28124\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28101\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28022\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27986\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27900\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27722\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27705\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27638\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27581\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27547\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27515\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27512\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27499\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27478\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27475\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27437\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27420\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27369\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27355\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27274\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27244\ : std_logic;
signal \N__27241\ : std_logic;
signal \N__27238\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27198\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27191\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27178\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27167\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27164\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27040\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26994\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26973\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26949\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26930\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26897\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26872\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26687\ : std_logic;
signal \N__26684\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26640\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26547\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26481\ : std_logic;
signal \N__26478\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26430\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26424\ : std_logic;
signal \N__26421\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26301\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26238\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26217\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26109\ : std_logic;
signal \N__26106\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26094\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26037\ : std_logic;
signal \N__26034\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26014\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25908\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25710\ : std_logic;
signal \N__25707\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25491\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25481\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25448\ : std_logic;
signal \N__25445\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25323\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25203\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25122\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24990\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24978\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24897\ : std_logic;
signal \N__24894\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24735\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24576\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24522\ : std_logic;
signal \N__24519\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24504\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24444\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24396\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24253\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23970\ : std_logic;
signal \N__23967\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23943\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23895\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23760\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23559\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23451\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23442\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23280\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23115\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22749\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21534\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21000\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20919\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20715\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20613\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20556\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20538\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20529\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20460\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20010\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19647\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19515\ : std_logic;
signal delay_tr_input_ibuf_gb_io_gb_input : std_logic;
signal delay_hc_input_ibuf_gb_io_gb_input : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_149\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_15\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_20\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_21\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_22\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_23\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_24\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_25\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\ : std_logic;
signal \bfn_1_16_0_\ : std_logic;
signal un7_start_stop_0_a2 : std_logic;
signal \N_38_i_i\ : std_logic;
signal pwm_duty_input_0 : std_logic;
signal pwm_duty_input_1 : std_logic;
signal pwm_duty_input_2 : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_3\ : std_logic;
signal pwm_duty_input_7 : std_logic;
signal pwm_duty_input_8 : std_logic;
signal pwm_duty_input_9 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\ : std_logic;
signal pwm_duty_input_6 : std_logic;
signal \current_shift_inst.PI_CTRL.N_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_153\ : std_logic;
signal pwm_duty_input_5 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\ : std_logic;
signal pwm_duty_input_4 : std_logic;
signal pwm_duty_input_3 : std_logic;
signal \pwm_generator_inst.un1_duty_inputlt3\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_154\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_155\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_7\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_6\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_4\ : std_logic;
signal \bfn_2_14_0_\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_0\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_1\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_2\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\ : std_logic;
signal \bfn_2_15_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\ : std_logic;
signal \bfn_2_16_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_19\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_0\ : std_logic;
signal \bfn_2_18_0_\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_2\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_4\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_6\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_7\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_7\ : std_logic;
signal \bfn_2_19_0_\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_118\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_1\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_3_11_0_\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_3_12_0_\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\ : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_0\ : std_logic;
signal \bfn_3_15_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_8\ : std_logic;
signal \bfn_3_16_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\ : std_logic;
signal \bfn_3_17_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_5\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_0\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_0\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_5\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_9\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_9\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_8\ : std_logic;
signal \pwm_generator_inst.N_16\ : std_logic;
signal \N_19_1\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\ : std_logic;
signal \pwm_generator_inst.N_17\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_53\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \bfn_4_12_0_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \bfn_4_13_0_\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_10\ : std_logic;
signal il_max_comp2_c : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal \bfn_5_9_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal \bfn_5_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \bfn_5_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \bfn_5_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \il_max_comp2_D1\ : std_logic;
signal il_min_comp2_c : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\ : std_logic;
signal \il_min_comp2_D1\ : std_logic;
signal \phase_controller_inst2.start_timer_tr_0_sqmuxa\ : std_logic;
signal \il_max_comp2_D2\ : std_logic;
signal \il_min_comp2_D2\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_393_i\ : std_logic;
signal \phase_controller_inst2.start_timer_hc_RNO_0_0\ : std_logic;
signal \phase_controller_inst2.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_inst2.start_timer_hcZ0\ : std_logic;
signal start_stop_c : std_logic;
signal \phase_controller_inst2.stateZ0Z_1\ : std_logic;
signal s4_phy_c : std_logic;
signal il_max_comp1_c : std_logic;
signal \il_max_comp1_D1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_13_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_72\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst2.state_RNI9M3OZ0Z_0\ : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \bfn_8_16_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \bfn_8_17_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \bfn_8_18_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_394_i\ : std_logic;
signal \phase_controller_inst1.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\ : std_logic;
signal \bfn_8_23_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIM9HS1Z0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \bfn_8_24_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_8_25_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\ : std_logic;
signal \bfn_8_26_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_3\ : std_logic;
signal s3_phy_c : std_logic;
signal il_min_comp1_c : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal delay_hc_input_c_g : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNID56UZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNILF8UZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIISQ01Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \bfn_9_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_30\ : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIUE3CP1_0_6_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIFFC6P1_0_16_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \elapsed_time_ns_1_RNILGKEE1_0_4_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_342_i_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIHHC6P1_0_18_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17\ : std_logic;
signal \elapsed_time_ns_1_RNIFFC6P1_0_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_267_iZ0Z_1_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_267_iZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_9_22_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_9_23_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_16\ : std_logic;
signal \bfn_9_24_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_df24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_df20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_df22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_df26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_df28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_71\ : std_logic;
signal \pll_inst.red_c_i\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI1M2UZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_enablelt3_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVHZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIM1S01Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIHA7UZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI905UZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIQ6T01Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_i_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI7T941Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_75\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_74\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIJEKEE1_0_2_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_284\ : std_logic;
signal \elapsed_time_ns_1_RNIJEKEE1_0_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\ : std_logic;
signal \elapsed_time_ns_1_RNI1I3CP1_0_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_326_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_308\ : std_logic;
signal \elapsed_time_ns_1_RNILGKEE1_0_4\ : std_logic;
signal \elapsed_time_ns_1_RNIAMU8E1_0_27\ : std_logic;
signal \elapsed_time_ns_1_RNIAMU8E1_0_27_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI6IU8E1_0_23\ : std_logic;
signal \elapsed_time_ns_1_RNI6IU8E1_0_23_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_1\ : std_logic;
signal \elapsed_time_ns_1_RNI9LU8E1_0_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlt31_0_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI5HU8E1_0_22\ : std_logic;
signal \elapsed_time_ns_1_RNI7JU8E1_0_24\ : std_logic;
signal \elapsed_time_ns_1_RNIBNU8E1_0_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_365_clk_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_367\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIDDC6P1_0_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14\ : std_logic;
signal \elapsed_time_ns_1_RNIMHKEE1_0_5\ : std_logic;
signal \elapsed_time_ns_1_RNI5IV8E1_0_31_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\ : std_logic;
signal \bfn_10_19_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \bfn_10_20_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_10_21_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \bfn_10_22_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_393_i_g\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \elapsed_time_ns_1_RNIGGC6P1_0_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_8\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74KZ0\ : std_logic;
signal \il_min_comp1_D1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_i_0_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7JZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3\ : std_logic;
signal \elapsed_time_ns_1_RNIRB3CP1_0_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIOJKEE1_0_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2\ : std_logic;
signal \elapsed_time_ns_1_RNI7IT8E1_0_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIUE3CP1_0_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_328_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst2.hc_time_passed\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \elapsed_time_ns_1_RNICOU8E1_0_29\ : std_logic;
signal \elapsed_time_ns_1_RNI4GU8E1_0_21\ : std_logic;
signal \elapsed_time_ns_1_RNICOU8E1_0_29_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un2_start_0\ : std_logic;
signal \elapsed_time_ns_1_RNI8KU8E1_0_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\ : std_logic;
signal \elapsed_time_ns_1_RNI2DT8E1_0_10_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\ : std_logic;
signal \elapsed_time_ns_1_RNI4HV8E1_0_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_342_i\ : std_logic;
signal \elapsed_time_ns_1_RNIP93CP1_0_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_16_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31\ : std_logic;
signal \elapsed_time_ns_1_RNI3FU8E1_0_20\ : std_logic;
signal \elapsed_time_ns_1_RNI2DT8E1_0_10\ : std_logic;
signal \elapsed_time_ns_1_RNI3ET8E1_0_11\ : std_logic;
signal \elapsed_time_ns_1_RNI4FT8E1_0_12\ : std_logic;
signal \elapsed_time_ns_1_RNI5GT8E1_0_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_316\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\ : std_logic;
signal \elapsed_time_ns_1_RNIHHC6P1_0_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \elapsed_time_ns_1_RNIPKKEE1_0_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_365_clk\ : std_logic;
signal \elapsed_time_ns_1_RNIIIC6P1_0_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latchedZ0\ : std_logic;
signal state_ns_i_a2_1 : std_logic;
signal \phase_controller_inst1.start_timer_hc_RNOZ0Z_0\ : std_logic;
signal \phase_controller_inst1.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \il_max_comp1_D2\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_395_i\ : std_logic;
signal delay_tr_input_c_g : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI5R3UZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axb_0\ : std_logic;
signal \bfn_12_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_7\ : std_logic;
signal \bfn_12_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_328\ : std_logic;
signal \elapsed_time_ns_1_RNI5IV8E1_0_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_326\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_12_14_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_12_15_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\ : std_logic;
signal \bfn_12_16_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\ : std_logic;
signal \bfn_12_17_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNITOIN1Z0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_12_18_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \bfn_12_19_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\ : std_logic;
signal \bfn_12_20_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\ : std_logic;
signal \il_min_comp1_D2\ : std_logic;
signal \T12_c\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \T01_c\ : std_logic;
signal \bfn_13_7_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \bfn_13_8_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \bfn_13_9_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.control_input_18\ : std_logic;
signal \bfn_13_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\ : std_logic;
signal \current_shift_inst.control_input_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\ : std_logic;
signal \current_shift_inst.control_input_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\ : std_logic;
signal \current_shift_inst.control_input_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\ : std_logic;
signal \current_shift_inst.control_input_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\ : std_logic;
signal \current_shift_inst.control_input_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\ : std_logic;
signal \current_shift_inst.control_input_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\ : std_logic;
signal \current_shift_inst.control_input_cry_6\ : std_logic;
signal \current_shift_inst.control_input_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\ : std_logic;
signal \bfn_13_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\ : std_logic;
signal \current_shift_inst.control_input_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\ : std_logic;
signal \current_shift_inst.control_input_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\ : std_logic;
signal \current_shift_inst.control_input_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\ : std_logic;
signal \current_shift_inst.control_input_cry_11\ : std_logic;
signal \current_shift_inst.control_input_cry_12\ : std_logic;
signal \current_shift_inst.control_input_31\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst2.tr_time_passed\ : std_logic;
signal \phase_controller_inst2.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_13_16_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_13_17_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_16\ : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_df26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_df28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_df22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_df24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_df26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_df28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_df20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_df22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_df20\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \phase_controller_inst1.start_timer_tr_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.time_passed_RNI7NN7\ : std_logic;
signal phase_controller_inst1_state_4 : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \current_shift_inst.timer_s1.N_166_i\ : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal s1_phy_c : std_logic;
signal \T23_c\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal state_3 : std_logic;
signal \T45_c\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal s2_phy_c : std_logic;
signal \bfn_14_5_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \bfn_14_6_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \bfn_14_7_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \bfn_14_8_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.timer_s1.N_167_i\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINRRH_1_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\ : std_logic;
signal \current_shift_inst.control_input_axb_0\ : std_logic;
signal \current_shift_inst.control_input_axb_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_fast_31\ : std_logic;
signal \current_shift_inst.control_input_axb_1\ : std_logic;
signal \current_shift_inst.control_input_axb_12\ : std_logic;
signal \current_shift_inst.N_1460_i\ : std_logic;
signal \current_shift_inst.control_input_axb_2\ : std_logic;
signal \current_shift_inst.control_input_axb_3\ : std_logic;
signal \current_shift_inst.control_input_axb_4\ : std_logic;
signal \current_shift_inst.control_input_axb_5\ : std_logic;
signal \current_shift_inst.control_input_axb_6\ : std_logic;
signal \current_shift_inst.control_input_axb_7\ : std_logic;
signal \current_shift_inst.control_input_axb_8\ : std_logic;
signal \current_shift_inst.control_input_axb_9\ : std_logic;
signal \current_shift_inst.control_input_axb_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIQU8A2Z0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_df24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\ : std_logic;
signal \bfn_14_21_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIJF7V2Z0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \bfn_14_22_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_14_23_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\ : std_logic;
signal \bfn_14_24_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\ : std_logic;
signal \bfn_15_8_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7\ : std_logic;
signal \bfn_15_9_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15\ : std_logic;
signal \bfn_15_10_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23\ : std_logic;
signal \bfn_15_11_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30\ : std_logic;
signal \bfn_15_12_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\ : std_logic;
signal \bfn_15_13_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0\ : std_logic;
signal \bfn_15_14_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_24\ : std_logic;
signal \bfn_15_15_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s0\ : std_logic;
signal \current_shift_inst.control_input_axb_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_242_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt16\ : std_logic;
signal \elapsed_time_ns_1_RNIQENQL1_0_9_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_15_20_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_15_21_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_16\ : std_logic;
signal \bfn_15_22_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_df20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_df22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_df24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_df28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_df26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_axb_31_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0_sf\ : std_logic;
signal \current_shift_inst.un4_control_input1_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_1_cascade_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\ : std_logic;
signal \elapsed_time_ns_1_RNISAHF91_0_13_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \elapsed_time_ns_1_RNIVEIF91_0_25\ : std_logic;
signal \elapsed_time_ns_1_RNI1HIF91_0_27\ : std_logic;
signal \elapsed_time_ns_1_RNIVEIF91_0_25_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNISBIF91_0_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI2IIF91_0_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI0GIF91_0_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17\ : std_logic;
signal \delay_measurement_inst.delay_tr9_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_390\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_390_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_391_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI6565M1_0_14_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_382\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_382_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_371\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_356\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_351_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_378\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_360\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_242\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1\ : std_logic;
signal \bfn_17_7_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.un4_control_input1_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.un4_control_input1_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un4_control_input1_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input1_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un4_control_input1_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_9\ : std_logic;
signal \current_shift_inst.un4_control_input1_10\ : std_logic;
signal \bfn_17_8_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_17\ : std_logic;
signal \bfn_17_9_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.un4_control_input1_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_25\ : std_logic;
signal \current_shift_inst.un4_control_input1_26\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_26\ : std_logic;
signal \current_shift_inst.un4_control_input1_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_27\ : std_logic;
signal \current_shift_inst.un4_control_input1_28\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_29\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_29\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.un4_control_input1_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.un4_control_input1_25\ : std_logic;
signal \current_shift_inst.un38_control_input_5_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\ : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1\ : std_logic;
signal \bfn_17_12_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1\ : std_logic;
signal \bfn_17_13_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_24\ : std_logic;
signal \bfn_17_14_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_26\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_28\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_31\ : std_logic;
signal \elapsed_time_ns_1_RNIP7HF91_0_10\ : std_logic;
signal \elapsed_time_ns_1_RNIR9HF91_0_12\ : std_logic;
signal \elapsed_time_ns_1_RNISAHF91_0_13\ : std_logic;
signal \elapsed_time_ns_1_RNIP7HF91_0_10_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI6565M1_0_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIQENQL1_0_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_0_6_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIK8NQL1_0_3_cascade_\ : std_logic;
signal \delay_measurement_inst.N_363\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIBA65M1_0_19_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_9\ : std_logic;
signal \elapsed_time_ns_1_RNIQ9IF91_0_20\ : std_logic;
signal \elapsed_time_ns_1_RNIQ9IF91_0_20_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIRAIF91_0_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15\ : std_logic;
signal \elapsed_time_ns_1_RNIQ8HF91_0_11\ : std_logic;
signal \elapsed_time_ns_1_RNI3JIF91_0_29\ : std_logic;
signal \elapsed_time_ns_1_RNITCIF91_0_23\ : std_logic;
signal \elapsed_time_ns_1_RNITCIF91_0_23_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIUDIF91_0_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15\ : std_logic;
signal \elapsed_time_ns_1_RNIA965M1_0_18\ : std_logic;
signal \elapsed_time_ns_1_RNICG2591_0_4_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI9865M1_0_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIRBJF91_0_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_344\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_344_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_347\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_347_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_373_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_351\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_353\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_348\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\ : std_logic;
signal \bfn_17_19_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\ : std_logic;
signal \bfn_17_20_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \bfn_17_21_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \bfn_17_22_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.un4_control_input1_17\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.un4_control_input1_14\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.un4_control_input1_7\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.un4_control_input1_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.timer_s1.N_166_i_g\ : std_logic;
signal \current_shift_inst.un38_control_input_5_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31_rep1\ : std_logic;
signal \current_shift_inst.un4_control_input1_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.un4_control_input1_16\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.un4_control_input1_13\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.un4_control_input1_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.un4_control_input1_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_11\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.un4_control_input1_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\ : std_logic;
signal \current_shift_inst.un4_control_input1_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_19\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.un4_control_input1_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.un4_control_input1_18\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.un4_control_input1_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_5_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \elapsed_time_ns_1_RNIDH2591_0_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \elapsed_time_ns_1_RNI8765M1_0_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \elapsed_time_ns_1_RNIK8NQL1_0_3\ : std_logic;
signal \elapsed_time_ns_1_RNIAE2591_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2Z0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNINBNQL1_0_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2\ : std_logic;
signal \elapsed_time_ns_1_RNIUCHF91_0_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \elapsed_time_ns_1_RNINBNQL1_0_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \bfn_18_18_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \bfn_18_19_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \bfn_18_20_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \bfn_18_21_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_396_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\ : std_logic;
signal \elapsed_time_ns_1_RNIGK2591_0_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\ : std_logic;
signal \elapsed_time_ns_1_RNII6NQL1_0_1_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIBA65M1_0_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19\ : std_logic;
signal \delay_measurement_inst.delay_tr9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1\ : std_logic;
signal \elapsed_time_ns_1_RNIFJ2591_0_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \elapsed_time_ns_1_RNICG2591_0_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_395_i_g\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\ : std_logic;
signal \elapsed_time_ns_1_RNISCJF91_0_31\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\ : std_logic;
signal \elapsed_time_ns_1_RNII6NQL1_0_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5Z0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_100mhz_0 : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\ : std_logic;
signal red_c_g : std_logic;

signal reset_wire : std_logic;
signal \T01_wire\ : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal \T23_wire\ : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal \T12_wire\ : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal \T45_wire\ : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal rgb_r_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    T01 <= \T01_wire\;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    T23 <= \T23_wire\;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    s2_phy <= s2_phy_wire;
    T12 <= \T12_wire\;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    T45 <= \T45_wire\;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    rgb_r <= rgb_r_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\ <= '0'&\N__21925\&\N__21918\&\N__21923\&\N__21917\&\N__21924\&\N__21916\&\N__21926\&\N__21913\&\N__21919\&\N__21912\&\N__21920\&\N__21914\&\N__21921\&\N__21915\&\N__21922\;
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__38281\&\N__38278\&'0'&'0'&'0'&\N__38276\&\N__38280\&\N__38277\&\N__38279\;
    \pwm_generator_inst.un2_threshold_acc_2_1_16\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_acc_2_1_15\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.un2_threshold_acc_2_14\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.un2_threshold_acc_2_13\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.un2_threshold_acc_2_12\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_acc_2_11\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_acc_2_10\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_acc_2_9\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_acc_2_8\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_acc_2_7\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_acc_2_6\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_acc_2_5\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_acc_2_4\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_acc_2_3\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_acc_2_2\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_acc_2_1\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_acc_2_0\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\ <= '0'&\N__21853\&\N__21891\&\N__21854\&\N__21892\&\N__21855\&\N__20353\&\N__20368\&\N__20079\&\N__20337\&\N__20261\&\N__20218\&\N__20204\&\N__20105\&\N__20121\&\N__20136\;
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__38249\&\N__38246\&'0'&'0'&'0'&\N__38244\&\N__38248\&\N__38245\&\N__38247\;
    \pwm_generator_inst.un2_threshold_acc_1_25\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(25);
    \pwm_generator_inst.un2_threshold_acc_1_24\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(24);
    \pwm_generator_inst.un2_threshold_acc_1_23\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(23);
    \pwm_generator_inst.un2_threshold_acc_1_22\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(22);
    \pwm_generator_inst.un2_threshold_acc_1_21\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(21);
    \pwm_generator_inst.un2_threshold_acc_1_20\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(20);
    \pwm_generator_inst.un2_threshold_acc_1_19\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_acc_1_18\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_acc_1_17\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_acc_1_16\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_acc_1_15\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un3_threshold_acc\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__32022\,
            RESETB => \N__25983\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clk_100mhz_0
        );

    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__38282\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__38275\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__38250\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__38243\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__50614\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50616\,
            DIN => \N__50615\,
            DOUT => \N__50614\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50616\,
            PADOUT => \N__50615\,
            PADIN => \N__50614\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T01_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50605\,
            DIN => \N__50604\,
            DOUT => \N__50603\,
            PACKAGEPIN => \T01_wire\
        );

    \T01_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50605\,
            PADOUT => \N__50604\,
            PADIN => \N__50603\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__34278\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50596\,
            DIN => \N__50595\,
            DOUT => \N__50594\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50596\,
            PADOUT => \N__50595\,
            PADIN => \N__50594\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50587\,
            DIN => \N__50586\,
            DOUT => \N__50585\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50587\,
            PADOUT => \N__50586\,
            PADIN => \N__50585\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T23_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50578\,
            DIN => \N__50577\,
            DOUT => \N__50576\,
            PACKAGEPIN => \T23_wire\
        );

    \T23_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50578\,
            PADOUT => \N__50577\,
            PADIN => \N__50576\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35700\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50569\,
            DIN => \N__50568\,
            DOUT => \N__50567\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50569\,
            PADOUT => \N__50568\,
            PADIN => \N__50567\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21009\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50560\,
            DIN => \N__50559\,
            DOUT => \N__50558\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50560\,
            PADOUT => \N__50559\,
            PADIN => \N__50558\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50551\,
            DIN => \N__50550\,
            DOUT => \N__50549\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50551\,
            PADOUT => \N__50550\,
            PADIN => \N__50549\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35508\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T12_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50542\,
            DIN => \N__50541\,
            DOUT => \N__50540\,
            PACKAGEPIN => \T12_wire\
        );

    \T12_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50542\,
            PADOUT => \N__50541\,
            PADIN => \N__50540\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__34335\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50533\,
            DIN => \N__50532\,
            DOUT => \N__50531\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50533\,
            PADOUT => \N__50532\,
            PADIN => \N__50531\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50524\,
            DIN => \N__50523\,
            DOUT => \N__50522\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50524\,
            PADOUT => \N__50523\,
            PADIN => \N__50522\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35727\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50515\,
            DIN => \N__50514\,
            DOUT => \N__50513\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50515\,
            PADOUT => \N__50514\,
            PADIN => \N__50513\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23532\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50506\,
            DIN => \N__50505\,
            DOUT => \N__50504\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50506\,
            PADOUT => \N__50505\,
            PADIN => \N__50504\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50497\,
            DIN => \N__50496\,
            DOUT => \N__50495\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50497\,
            PADOUT => \N__50496\,
            PADIN => \N__50495\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24522\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T45_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50488\,
            DIN => \N__50487\,
            DOUT => \N__50486\,
            PACKAGEPIN => \T45_wire\
        );

    \T45_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50488\,
            PADOUT => \N__50487\,
            PADIN => \N__50486\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35592\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50479\,
            DIN => \N__50478\,
            DOUT => \N__50477\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50479\,
            PADOUT => \N__50478\,
            PADIN => \N__50477\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50470\,
            DIN => \N__50469\,
            DOUT => \N__50468\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50470\,
            PADOUT => \N__50469\,
            PADIN => \N__50468\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__11944\ : InMux
    port map (
            O => \N__50451\,
            I => \N__50448\
        );

    \I__11943\ : LocalMux
    port map (
            O => \N__50448\,
            I => \N__50444\
        );

    \I__11942\ : InMux
    port map (
            O => \N__50447\,
            I => \N__50441\
        );

    \I__11941\ : Odrv4
    port map (
            O => \N__50444\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2\
        );

    \I__11940\ : LocalMux
    port map (
            O => \N__50441\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2\
        );

    \I__11939\ : InMux
    port map (
            O => \N__50436\,
            I => \N__50433\
        );

    \I__11938\ : LocalMux
    port map (
            O => \N__50433\,
            I => \N__50430\
        );

    \I__11937\ : Odrv12
    port map (
            O => \N__50430\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\
        );

    \I__11936\ : CascadeMux
    port map (
            O => \N__50427\,
            I => \N__50424\
        );

    \I__11935\ : InMux
    port map (
            O => \N__50424\,
            I => \N__50421\
        );

    \I__11934\ : LocalMux
    port map (
            O => \N__50421\,
            I => \N__50417\
        );

    \I__11933\ : InMux
    port map (
            O => \N__50420\,
            I => \N__50413\
        );

    \I__11932\ : Span4Mux_h
    port map (
            O => \N__50417\,
            I => \N__50410\
        );

    \I__11931\ : InMux
    port map (
            O => \N__50416\,
            I => \N__50407\
        );

    \I__11930\ : LocalMux
    port map (
            O => \N__50413\,
            I => \elapsed_time_ns_1_RNICG2591_0_4\
        );

    \I__11929\ : Odrv4
    port map (
            O => \N__50410\,
            I => \elapsed_time_ns_1_RNICG2591_0_4\
        );

    \I__11928\ : LocalMux
    port map (
            O => \N__50407\,
            I => \elapsed_time_ns_1_RNICG2591_0_4\
        );

    \I__11927\ : CascadeMux
    port map (
            O => \N__50400\,
            I => \N__50396\
        );

    \I__11926\ : CascadeMux
    port map (
            O => \N__50399\,
            I => \N__50387\
        );

    \I__11925\ : InMux
    port map (
            O => \N__50396\,
            I => \N__50376\
        );

    \I__11924\ : InMux
    port map (
            O => \N__50395\,
            I => \N__50376\
        );

    \I__11923\ : InMux
    port map (
            O => \N__50394\,
            I => \N__50376\
        );

    \I__11922\ : InMux
    port map (
            O => \N__50393\,
            I => \N__50371\
        );

    \I__11921\ : InMux
    port map (
            O => \N__50392\,
            I => \N__50371\
        );

    \I__11920\ : InMux
    port map (
            O => \N__50391\,
            I => \N__50368\
        );

    \I__11919\ : InMux
    port map (
            O => \N__50390\,
            I => \N__50363\
        );

    \I__11918\ : InMux
    port map (
            O => \N__50387\,
            I => \N__50363\
        );

    \I__11917\ : InMux
    port map (
            O => \N__50386\,
            I => \N__50360\
        );

    \I__11916\ : InMux
    port map (
            O => \N__50385\,
            I => \N__50356\
        );

    \I__11915\ : InMux
    port map (
            O => \N__50384\,
            I => \N__50353\
        );

    \I__11914\ : CascadeMux
    port map (
            O => \N__50383\,
            I => \N__50350\
        );

    \I__11913\ : LocalMux
    port map (
            O => \N__50376\,
            I => \N__50345\
        );

    \I__11912\ : LocalMux
    port map (
            O => \N__50371\,
            I => \N__50342\
        );

    \I__11911\ : LocalMux
    port map (
            O => \N__50368\,
            I => \N__50337\
        );

    \I__11910\ : LocalMux
    port map (
            O => \N__50363\,
            I => \N__50337\
        );

    \I__11909\ : LocalMux
    port map (
            O => \N__50360\,
            I => \N__50334\
        );

    \I__11908\ : InMux
    port map (
            O => \N__50359\,
            I => \N__50331\
        );

    \I__11907\ : LocalMux
    port map (
            O => \N__50356\,
            I => \N__50326\
        );

    \I__11906\ : LocalMux
    port map (
            O => \N__50353\,
            I => \N__50326\
        );

    \I__11905\ : InMux
    port map (
            O => \N__50350\,
            I => \N__50319\
        );

    \I__11904\ : InMux
    port map (
            O => \N__50349\,
            I => \N__50319\
        );

    \I__11903\ : InMux
    port map (
            O => \N__50348\,
            I => \N__50319\
        );

    \I__11902\ : Span4Mux_v
    port map (
            O => \N__50345\,
            I => \N__50316\
        );

    \I__11901\ : Span4Mux_v
    port map (
            O => \N__50342\,
            I => \N__50309\
        );

    \I__11900\ : Span4Mux_v
    port map (
            O => \N__50337\,
            I => \N__50309\
        );

    \I__11899\ : Span4Mux_v
    port map (
            O => \N__50334\,
            I => \N__50309\
        );

    \I__11898\ : LocalMux
    port map (
            O => \N__50331\,
            I => \N__50306\
        );

    \I__11897\ : Odrv4
    port map (
            O => \N__50326\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6\
        );

    \I__11896\ : LocalMux
    port map (
            O => \N__50319\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6\
        );

    \I__11895\ : Odrv4
    port map (
            O => \N__50316\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6\
        );

    \I__11894\ : Odrv4
    port map (
            O => \N__50309\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6\
        );

    \I__11893\ : Odrv4
    port map (
            O => \N__50306\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6\
        );

    \I__11892\ : InMux
    port map (
            O => \N__50295\,
            I => \N__50292\
        );

    \I__11891\ : LocalMux
    port map (
            O => \N__50292\,
            I => \N__50289\
        );

    \I__11890\ : Odrv12
    port map (
            O => \N__50289\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\
        );

    \I__11889\ : CEMux
    port map (
            O => \N__50286\,
            I => \N__50281\
        );

    \I__11888\ : CEMux
    port map (
            O => \N__50285\,
            I => \N__50273\
        );

    \I__11887\ : CEMux
    port map (
            O => \N__50284\,
            I => \N__50270\
        );

    \I__11886\ : LocalMux
    port map (
            O => \N__50281\,
            I => \N__50267\
        );

    \I__11885\ : CEMux
    port map (
            O => \N__50280\,
            I => \N__50264\
        );

    \I__11884\ : InMux
    port map (
            O => \N__50279\,
            I => \N__50252\
        );

    \I__11883\ : InMux
    port map (
            O => \N__50278\,
            I => \N__50252\
        );

    \I__11882\ : InMux
    port map (
            O => \N__50277\,
            I => \N__50252\
        );

    \I__11881\ : CEMux
    port map (
            O => \N__50276\,
            I => \N__50234\
        );

    \I__11880\ : LocalMux
    port map (
            O => \N__50273\,
            I => \N__50231\
        );

    \I__11879\ : LocalMux
    port map (
            O => \N__50270\,
            I => \N__50226\
        );

    \I__11878\ : Span4Mux_v
    port map (
            O => \N__50267\,
            I => \N__50226\
        );

    \I__11877\ : LocalMux
    port map (
            O => \N__50264\,
            I => \N__50223\
        );

    \I__11876\ : InMux
    port map (
            O => \N__50263\,
            I => \N__50214\
        );

    \I__11875\ : InMux
    port map (
            O => \N__50262\,
            I => \N__50214\
        );

    \I__11874\ : InMux
    port map (
            O => \N__50261\,
            I => \N__50214\
        );

    \I__11873\ : InMux
    port map (
            O => \N__50260\,
            I => \N__50214\
        );

    \I__11872\ : CEMux
    port map (
            O => \N__50259\,
            I => \N__50211\
        );

    \I__11871\ : LocalMux
    port map (
            O => \N__50252\,
            I => \N__50208\
        );

    \I__11870\ : InMux
    port map (
            O => \N__50251\,
            I => \N__50201\
        );

    \I__11869\ : InMux
    port map (
            O => \N__50250\,
            I => \N__50201\
        );

    \I__11868\ : InMux
    port map (
            O => \N__50249\,
            I => \N__50201\
        );

    \I__11867\ : InMux
    port map (
            O => \N__50248\,
            I => \N__50192\
        );

    \I__11866\ : InMux
    port map (
            O => \N__50247\,
            I => \N__50192\
        );

    \I__11865\ : InMux
    port map (
            O => \N__50246\,
            I => \N__50192\
        );

    \I__11864\ : InMux
    port map (
            O => \N__50245\,
            I => \N__50192\
        );

    \I__11863\ : InMux
    port map (
            O => \N__50244\,
            I => \N__50183\
        );

    \I__11862\ : InMux
    port map (
            O => \N__50243\,
            I => \N__50183\
        );

    \I__11861\ : InMux
    port map (
            O => \N__50242\,
            I => \N__50183\
        );

    \I__11860\ : InMux
    port map (
            O => \N__50241\,
            I => \N__50183\
        );

    \I__11859\ : InMux
    port map (
            O => \N__50240\,
            I => \N__50174\
        );

    \I__11858\ : InMux
    port map (
            O => \N__50239\,
            I => \N__50174\
        );

    \I__11857\ : InMux
    port map (
            O => \N__50238\,
            I => \N__50174\
        );

    \I__11856\ : InMux
    port map (
            O => \N__50237\,
            I => \N__50174\
        );

    \I__11855\ : LocalMux
    port map (
            O => \N__50234\,
            I => \N__50171\
        );

    \I__11854\ : Span4Mux_v
    port map (
            O => \N__50231\,
            I => \N__50167\
        );

    \I__11853\ : Span4Mux_h
    port map (
            O => \N__50226\,
            I => \N__50164\
        );

    \I__11852\ : Span4Mux_v
    port map (
            O => \N__50223\,
            I => \N__50153\
        );

    \I__11851\ : LocalMux
    port map (
            O => \N__50214\,
            I => \N__50150\
        );

    \I__11850\ : LocalMux
    port map (
            O => \N__50211\,
            I => \N__50137\
        );

    \I__11849\ : Span4Mux_v
    port map (
            O => \N__50208\,
            I => \N__50137\
        );

    \I__11848\ : LocalMux
    port map (
            O => \N__50201\,
            I => \N__50137\
        );

    \I__11847\ : LocalMux
    port map (
            O => \N__50192\,
            I => \N__50137\
        );

    \I__11846\ : LocalMux
    port map (
            O => \N__50183\,
            I => \N__50137\
        );

    \I__11845\ : LocalMux
    port map (
            O => \N__50174\,
            I => \N__50137\
        );

    \I__11844\ : Span4Mux_v
    port map (
            O => \N__50171\,
            I => \N__50134\
        );

    \I__11843\ : InMux
    port map (
            O => \N__50170\,
            I => \N__50131\
        );

    \I__11842\ : Span4Mux_h
    port map (
            O => \N__50167\,
            I => \N__50126\
        );

    \I__11841\ : Span4Mux_h
    port map (
            O => \N__50164\,
            I => \N__50126\
        );

    \I__11840\ : InMux
    port map (
            O => \N__50163\,
            I => \N__50117\
        );

    \I__11839\ : InMux
    port map (
            O => \N__50162\,
            I => \N__50117\
        );

    \I__11838\ : InMux
    port map (
            O => \N__50161\,
            I => \N__50117\
        );

    \I__11837\ : InMux
    port map (
            O => \N__50160\,
            I => \N__50117\
        );

    \I__11836\ : InMux
    port map (
            O => \N__50159\,
            I => \N__50108\
        );

    \I__11835\ : InMux
    port map (
            O => \N__50158\,
            I => \N__50108\
        );

    \I__11834\ : InMux
    port map (
            O => \N__50157\,
            I => \N__50108\
        );

    \I__11833\ : InMux
    port map (
            O => \N__50156\,
            I => \N__50108\
        );

    \I__11832\ : Span4Mux_h
    port map (
            O => \N__50153\,
            I => \N__50101\
        );

    \I__11831\ : Span4Mux_v
    port map (
            O => \N__50150\,
            I => \N__50101\
        );

    \I__11830\ : Span4Mux_v
    port map (
            O => \N__50137\,
            I => \N__50101\
        );

    \I__11829\ : Span4Mux_h
    port map (
            O => \N__50134\,
            I => \N__50098\
        );

    \I__11828\ : LocalMux
    port map (
            O => \N__50131\,
            I => \N__50087\
        );

    \I__11827\ : Sp12to4
    port map (
            O => \N__50126\,
            I => \N__50087\
        );

    \I__11826\ : LocalMux
    port map (
            O => \N__50117\,
            I => \N__50087\
        );

    \I__11825\ : LocalMux
    port map (
            O => \N__50108\,
            I => \N__50087\
        );

    \I__11824\ : Sp12to4
    port map (
            O => \N__50101\,
            I => \N__50087\
        );

    \I__11823\ : Odrv4
    port map (
            O => \N__50098\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__11822\ : Odrv12
    port map (
            O => \N__50087\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__11821\ : InMux
    port map (
            O => \N__50082\,
            I => \N__50078\
        );

    \I__11820\ : CascadeMux
    port map (
            O => \N__50081\,
            I => \N__50075\
        );

    \I__11819\ : LocalMux
    port map (
            O => \N__50078\,
            I => \N__50071\
        );

    \I__11818\ : InMux
    port map (
            O => \N__50075\,
            I => \N__50068\
        );

    \I__11817\ : InMux
    port map (
            O => \N__50074\,
            I => \N__50065\
        );

    \I__11816\ : Odrv4
    port map (
            O => \N__50071\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__11815\ : LocalMux
    port map (
            O => \N__50068\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__11814\ : LocalMux
    port map (
            O => \N__50065\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__11813\ : CascadeMux
    port map (
            O => \N__50058\,
            I => \N__50055\
        );

    \I__11812\ : InMux
    port map (
            O => \N__50055\,
            I => \N__50051\
        );

    \I__11811\ : InMux
    port map (
            O => \N__50054\,
            I => \N__50048\
        );

    \I__11810\ : LocalMux
    port map (
            O => \N__50051\,
            I => \N__50045\
        );

    \I__11809\ : LocalMux
    port map (
            O => \N__50048\,
            I => \N__50042\
        );

    \I__11808\ : Odrv4
    port map (
            O => \N__50045\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__11807\ : Odrv12
    port map (
            O => \N__50042\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__11806\ : InMux
    port map (
            O => \N__50037\,
            I => \N__50033\
        );

    \I__11805\ : CascadeMux
    port map (
            O => \N__50036\,
            I => \N__50030\
        );

    \I__11804\ : LocalMux
    port map (
            O => \N__50033\,
            I => \N__50026\
        );

    \I__11803\ : InMux
    port map (
            O => \N__50030\,
            I => \N__50023\
        );

    \I__11802\ : InMux
    port map (
            O => \N__50029\,
            I => \N__50020\
        );

    \I__11801\ : Odrv4
    port map (
            O => \N__50026\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__11800\ : LocalMux
    port map (
            O => \N__50023\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__11799\ : LocalMux
    port map (
            O => \N__50020\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__11798\ : InMux
    port map (
            O => \N__50013\,
            I => \N__50010\
        );

    \I__11797\ : LocalMux
    port map (
            O => \N__50010\,
            I => \N__50005\
        );

    \I__11796\ : InMux
    port map (
            O => \N__50009\,
            I => \N__50000\
        );

    \I__11795\ : InMux
    port map (
            O => \N__50008\,
            I => \N__50000\
        );

    \I__11794\ : Span4Mux_v
    port map (
            O => \N__50005\,
            I => \N__49997\
        );

    \I__11793\ : LocalMux
    port map (
            O => \N__50000\,
            I => \N__49994\
        );

    \I__11792\ : Odrv4
    port map (
            O => \N__49997\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__11791\ : Odrv12
    port map (
            O => \N__49994\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__11790\ : CEMux
    port map (
            O => \N__49989\,
            I => \N__49974\
        );

    \I__11789\ : CEMux
    port map (
            O => \N__49988\,
            I => \N__49974\
        );

    \I__11788\ : CEMux
    port map (
            O => \N__49987\,
            I => \N__49974\
        );

    \I__11787\ : CEMux
    port map (
            O => \N__49986\,
            I => \N__49974\
        );

    \I__11786\ : CEMux
    port map (
            O => \N__49985\,
            I => \N__49974\
        );

    \I__11785\ : GlobalMux
    port map (
            O => \N__49974\,
            I => \N__49971\
        );

    \I__11784\ : gio2CtrlBuf
    port map (
            O => \N__49971\,
            I => \delay_measurement_inst.delay_tr_timer.N_395_i_g\
        );

    \I__11783\ : InMux
    port map (
            O => \N__49968\,
            I => \N__49964\
        );

    \I__11782\ : CascadeMux
    port map (
            O => \N__49967\,
            I => \N__49958\
        );

    \I__11781\ : LocalMux
    port map (
            O => \N__49964\,
            I => \N__49955\
        );

    \I__11780\ : InMux
    port map (
            O => \N__49963\,
            I => \N__49952\
        );

    \I__11779\ : InMux
    port map (
            O => \N__49962\,
            I => \N__49948\
        );

    \I__11778\ : InMux
    port map (
            O => \N__49961\,
            I => \N__49943\
        );

    \I__11777\ : InMux
    port map (
            O => \N__49958\,
            I => \N__49943\
        );

    \I__11776\ : Span4Mux_h
    port map (
            O => \N__49955\,
            I => \N__49940\
        );

    \I__11775\ : LocalMux
    port map (
            O => \N__49952\,
            I => \N__49937\
        );

    \I__11774\ : InMux
    port map (
            O => \N__49951\,
            I => \N__49934\
        );

    \I__11773\ : LocalMux
    port map (
            O => \N__49948\,
            I => \N__49931\
        );

    \I__11772\ : LocalMux
    port map (
            O => \N__49943\,
            I => \N__49928\
        );

    \I__11771\ : Span4Mux_v
    port map (
            O => \N__49940\,
            I => \N__49925\
        );

    \I__11770\ : Span12Mux_v
    port map (
            O => \N__49937\,
            I => \N__49922\
        );

    \I__11769\ : LocalMux
    port map (
            O => \N__49934\,
            I => \N__49919\
        );

    \I__11768\ : Span4Mux_v
    port map (
            O => \N__49931\,
            I => \N__49912\
        );

    \I__11767\ : Span4Mux_v
    port map (
            O => \N__49928\,
            I => \N__49912\
        );

    \I__11766\ : Span4Mux_h
    port map (
            O => \N__49925\,
            I => \N__49912\
        );

    \I__11765\ : Odrv12
    port map (
            O => \N__49922\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__11764\ : Odrv12
    port map (
            O => \N__49919\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__11763\ : Odrv4
    port map (
            O => \N__49912\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__11762\ : CascadeMux
    port map (
            O => \N__49905\,
            I => \N__49901\
        );

    \I__11761\ : InMux
    port map (
            O => \N__49904\,
            I => \N__49897\
        );

    \I__11760\ : InMux
    port map (
            O => \N__49901\,
            I => \N__49894\
        );

    \I__11759\ : InMux
    port map (
            O => \N__49900\,
            I => \N__49890\
        );

    \I__11758\ : LocalMux
    port map (
            O => \N__49897\,
            I => \N__49883\
        );

    \I__11757\ : LocalMux
    port map (
            O => \N__49894\,
            I => \N__49880\
        );

    \I__11756\ : InMux
    port map (
            O => \N__49893\,
            I => \N__49877\
        );

    \I__11755\ : LocalMux
    port map (
            O => \N__49890\,
            I => \N__49871\
        );

    \I__11754\ : InMux
    port map (
            O => \N__49889\,
            I => \N__49866\
        );

    \I__11753\ : InMux
    port map (
            O => \N__49888\,
            I => \N__49866\
        );

    \I__11752\ : CascadeMux
    port map (
            O => \N__49887\,
            I => \N__49857\
        );

    \I__11751\ : CascadeMux
    port map (
            O => \N__49886\,
            I => \N__49854\
        );

    \I__11750\ : Span4Mux_v
    port map (
            O => \N__49883\,
            I => \N__49849\
        );

    \I__11749\ : Span4Mux_v
    port map (
            O => \N__49880\,
            I => \N__49849\
        );

    \I__11748\ : LocalMux
    port map (
            O => \N__49877\,
            I => \N__49846\
        );

    \I__11747\ : CascadeMux
    port map (
            O => \N__49876\,
            I => \N__49842\
        );

    \I__11746\ : CascadeMux
    port map (
            O => \N__49875\,
            I => \N__49836\
        );

    \I__11745\ : InMux
    port map (
            O => \N__49874\,
            I => \N__49833\
        );

    \I__11744\ : Span4Mux_h
    port map (
            O => \N__49871\,
            I => \N__49828\
        );

    \I__11743\ : LocalMux
    port map (
            O => \N__49866\,
            I => \N__49828\
        );

    \I__11742\ : CascadeMux
    port map (
            O => \N__49865\,
            I => \N__49825\
        );

    \I__11741\ : CascadeMux
    port map (
            O => \N__49864\,
            I => \N__49822\
        );

    \I__11740\ : InMux
    port map (
            O => \N__49863\,
            I => \N__49806\
        );

    \I__11739\ : InMux
    port map (
            O => \N__49862\,
            I => \N__49806\
        );

    \I__11738\ : InMux
    port map (
            O => \N__49861\,
            I => \N__49806\
        );

    \I__11737\ : InMux
    port map (
            O => \N__49860\,
            I => \N__49801\
        );

    \I__11736\ : InMux
    port map (
            O => \N__49857\,
            I => \N__49801\
        );

    \I__11735\ : InMux
    port map (
            O => \N__49854\,
            I => \N__49798\
        );

    \I__11734\ : Span4Mux_h
    port map (
            O => \N__49849\,
            I => \N__49795\
        );

    \I__11733\ : Span4Mux_h
    port map (
            O => \N__49846\,
            I => \N__49792\
        );

    \I__11732\ : InMux
    port map (
            O => \N__49845\,
            I => \N__49783\
        );

    \I__11731\ : InMux
    port map (
            O => \N__49842\,
            I => \N__49783\
        );

    \I__11730\ : InMux
    port map (
            O => \N__49841\,
            I => \N__49783\
        );

    \I__11729\ : InMux
    port map (
            O => \N__49840\,
            I => \N__49783\
        );

    \I__11728\ : InMux
    port map (
            O => \N__49839\,
            I => \N__49778\
        );

    \I__11727\ : InMux
    port map (
            O => \N__49836\,
            I => \N__49778\
        );

    \I__11726\ : LocalMux
    port map (
            O => \N__49833\,
            I => \N__49775\
        );

    \I__11725\ : Span4Mux_v
    port map (
            O => \N__49828\,
            I => \N__49772\
        );

    \I__11724\ : InMux
    port map (
            O => \N__49825\,
            I => \N__49761\
        );

    \I__11723\ : InMux
    port map (
            O => \N__49822\,
            I => \N__49761\
        );

    \I__11722\ : InMux
    port map (
            O => \N__49821\,
            I => \N__49761\
        );

    \I__11721\ : InMux
    port map (
            O => \N__49820\,
            I => \N__49761\
        );

    \I__11720\ : InMux
    port map (
            O => \N__49819\,
            I => \N__49761\
        );

    \I__11719\ : InMux
    port map (
            O => \N__49818\,
            I => \N__49758\
        );

    \I__11718\ : InMux
    port map (
            O => \N__49817\,
            I => \N__49755\
        );

    \I__11717\ : InMux
    port map (
            O => \N__49816\,
            I => \N__49746\
        );

    \I__11716\ : InMux
    port map (
            O => \N__49815\,
            I => \N__49746\
        );

    \I__11715\ : InMux
    port map (
            O => \N__49814\,
            I => \N__49746\
        );

    \I__11714\ : InMux
    port map (
            O => \N__49813\,
            I => \N__49746\
        );

    \I__11713\ : LocalMux
    port map (
            O => \N__49806\,
            I => \N__49743\
        );

    \I__11712\ : LocalMux
    port map (
            O => \N__49801\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__11711\ : LocalMux
    port map (
            O => \N__49798\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__11710\ : Odrv4
    port map (
            O => \N__49795\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__11709\ : Odrv4
    port map (
            O => \N__49792\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__11708\ : LocalMux
    port map (
            O => \N__49783\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__11707\ : LocalMux
    port map (
            O => \N__49778\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__11706\ : Odrv4
    port map (
            O => \N__49775\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__11705\ : Odrv4
    port map (
            O => \N__49772\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__11704\ : LocalMux
    port map (
            O => \N__49761\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__11703\ : LocalMux
    port map (
            O => \N__49758\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__11702\ : LocalMux
    port map (
            O => \N__49755\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__11701\ : LocalMux
    port map (
            O => \N__49746\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__11700\ : Odrv4
    port map (
            O => \N__49743\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__11699\ : InMux
    port map (
            O => \N__49716\,
            I => \N__49712\
        );

    \I__11698\ : InMux
    port map (
            O => \N__49715\,
            I => \N__49706\
        );

    \I__11697\ : LocalMux
    port map (
            O => \N__49712\,
            I => \N__49702\
        );

    \I__11696\ : CascadeMux
    port map (
            O => \N__49711\,
            I => \N__49697\
        );

    \I__11695\ : CascadeMux
    port map (
            O => \N__49710\,
            I => \N__49693\
        );

    \I__11694\ : CascadeMux
    port map (
            O => \N__49709\,
            I => \N__49687\
        );

    \I__11693\ : LocalMux
    port map (
            O => \N__49706\,
            I => \N__49675\
        );

    \I__11692\ : InMux
    port map (
            O => \N__49705\,
            I => \N__49672\
        );

    \I__11691\ : Span4Mux_h
    port map (
            O => \N__49702\,
            I => \N__49669\
        );

    \I__11690\ : InMux
    port map (
            O => \N__49701\,
            I => \N__49666\
        );

    \I__11689\ : InMux
    port map (
            O => \N__49700\,
            I => \N__49663\
        );

    \I__11688\ : InMux
    port map (
            O => \N__49697\,
            I => \N__49650\
        );

    \I__11687\ : InMux
    port map (
            O => \N__49696\,
            I => \N__49650\
        );

    \I__11686\ : InMux
    port map (
            O => \N__49693\,
            I => \N__49650\
        );

    \I__11685\ : InMux
    port map (
            O => \N__49692\,
            I => \N__49650\
        );

    \I__11684\ : InMux
    port map (
            O => \N__49691\,
            I => \N__49650\
        );

    \I__11683\ : InMux
    port map (
            O => \N__49690\,
            I => \N__49650\
        );

    \I__11682\ : InMux
    port map (
            O => \N__49687\,
            I => \N__49645\
        );

    \I__11681\ : InMux
    port map (
            O => \N__49686\,
            I => \N__49645\
        );

    \I__11680\ : InMux
    port map (
            O => \N__49685\,
            I => \N__49634\
        );

    \I__11679\ : InMux
    port map (
            O => \N__49684\,
            I => \N__49634\
        );

    \I__11678\ : InMux
    port map (
            O => \N__49683\,
            I => \N__49634\
        );

    \I__11677\ : InMux
    port map (
            O => \N__49682\,
            I => \N__49634\
        );

    \I__11676\ : InMux
    port map (
            O => \N__49681\,
            I => \N__49634\
        );

    \I__11675\ : InMux
    port map (
            O => \N__49680\,
            I => \N__49627\
        );

    \I__11674\ : InMux
    port map (
            O => \N__49679\,
            I => \N__49627\
        );

    \I__11673\ : InMux
    port map (
            O => \N__49678\,
            I => \N__49627\
        );

    \I__11672\ : Odrv12
    port map (
            O => \N__49675\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__11671\ : LocalMux
    port map (
            O => \N__49672\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__11670\ : Odrv4
    port map (
            O => \N__49669\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__11669\ : LocalMux
    port map (
            O => \N__49666\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__11668\ : LocalMux
    port map (
            O => \N__49663\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__11667\ : LocalMux
    port map (
            O => \N__49650\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__11666\ : LocalMux
    port map (
            O => \N__49645\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__11665\ : LocalMux
    port map (
            O => \N__49634\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__11664\ : LocalMux
    port map (
            O => \N__49627\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__11663\ : CascadeMux
    port map (
            O => \N__49608\,
            I => \N__49603\
        );

    \I__11662\ : CascadeMux
    port map (
            O => \N__49607\,
            I => \N__49600\
        );

    \I__11661\ : InMux
    port map (
            O => \N__49606\,
            I => \N__49589\
        );

    \I__11660\ : InMux
    port map (
            O => \N__49603\,
            I => \N__49589\
        );

    \I__11659\ : InMux
    port map (
            O => \N__49600\,
            I => \N__49589\
        );

    \I__11658\ : CascadeMux
    port map (
            O => \N__49599\,
            I => \N__49586\
        );

    \I__11657\ : CascadeMux
    port map (
            O => \N__49598\,
            I => \N__49571\
        );

    \I__11656\ : CascadeMux
    port map (
            O => \N__49597\,
            I => \N__49568\
        );

    \I__11655\ : InMux
    port map (
            O => \N__49596\,
            I => \N__49561\
        );

    \I__11654\ : LocalMux
    port map (
            O => \N__49589\,
            I => \N__49558\
        );

    \I__11653\ : InMux
    port map (
            O => \N__49586\,
            I => \N__49545\
        );

    \I__11652\ : InMux
    port map (
            O => \N__49585\,
            I => \N__49545\
        );

    \I__11651\ : InMux
    port map (
            O => \N__49584\,
            I => \N__49545\
        );

    \I__11650\ : InMux
    port map (
            O => \N__49583\,
            I => \N__49545\
        );

    \I__11649\ : InMux
    port map (
            O => \N__49582\,
            I => \N__49545\
        );

    \I__11648\ : InMux
    port map (
            O => \N__49581\,
            I => \N__49545\
        );

    \I__11647\ : InMux
    port map (
            O => \N__49580\,
            I => \N__49542\
        );

    \I__11646\ : CascadeMux
    port map (
            O => \N__49579\,
            I => \N__49539\
        );

    \I__11645\ : InMux
    port map (
            O => \N__49578\,
            I => \N__49534\
        );

    \I__11644\ : InMux
    port map (
            O => \N__49577\,
            I => \N__49527\
        );

    \I__11643\ : InMux
    port map (
            O => \N__49576\,
            I => \N__49527\
        );

    \I__11642\ : InMux
    port map (
            O => \N__49575\,
            I => \N__49527\
        );

    \I__11641\ : InMux
    port map (
            O => \N__49574\,
            I => \N__49524\
        );

    \I__11640\ : InMux
    port map (
            O => \N__49571\,
            I => \N__49517\
        );

    \I__11639\ : InMux
    port map (
            O => \N__49568\,
            I => \N__49517\
        );

    \I__11638\ : InMux
    port map (
            O => \N__49567\,
            I => \N__49517\
        );

    \I__11637\ : InMux
    port map (
            O => \N__49566\,
            I => \N__49510\
        );

    \I__11636\ : InMux
    port map (
            O => \N__49565\,
            I => \N__49510\
        );

    \I__11635\ : InMux
    port map (
            O => \N__49564\,
            I => \N__49510\
        );

    \I__11634\ : LocalMux
    port map (
            O => \N__49561\,
            I => \N__49507\
        );

    \I__11633\ : Span4Mux_v
    port map (
            O => \N__49558\,
            I => \N__49502\
        );

    \I__11632\ : LocalMux
    port map (
            O => \N__49545\,
            I => \N__49502\
        );

    \I__11631\ : LocalMux
    port map (
            O => \N__49542\,
            I => \N__49499\
        );

    \I__11630\ : InMux
    port map (
            O => \N__49539\,
            I => \N__49491\
        );

    \I__11629\ : InMux
    port map (
            O => \N__49538\,
            I => \N__49491\
        );

    \I__11628\ : InMux
    port map (
            O => \N__49537\,
            I => \N__49491\
        );

    \I__11627\ : LocalMux
    port map (
            O => \N__49534\,
            I => \N__49486\
        );

    \I__11626\ : LocalMux
    port map (
            O => \N__49527\,
            I => \N__49486\
        );

    \I__11625\ : LocalMux
    port map (
            O => \N__49524\,
            I => \N__49483\
        );

    \I__11624\ : LocalMux
    port map (
            O => \N__49517\,
            I => \N__49480\
        );

    \I__11623\ : LocalMux
    port map (
            O => \N__49510\,
            I => \N__49475\
        );

    \I__11622\ : Span4Mux_v
    port map (
            O => \N__49507\,
            I => \N__49475\
        );

    \I__11621\ : Span4Mux_h
    port map (
            O => \N__49502\,
            I => \N__49470\
        );

    \I__11620\ : Span4Mux_h
    port map (
            O => \N__49499\,
            I => \N__49470\
        );

    \I__11619\ : CascadeMux
    port map (
            O => \N__49498\,
            I => \N__49461\
        );

    \I__11618\ : LocalMux
    port map (
            O => \N__49491\,
            I => \N__49455\
        );

    \I__11617\ : Span4Mux_v
    port map (
            O => \N__49486\,
            I => \N__49452\
        );

    \I__11616\ : Span4Mux_v
    port map (
            O => \N__49483\,
            I => \N__49446\
        );

    \I__11615\ : Span4Mux_v
    port map (
            O => \N__49480\,
            I => \N__49446\
        );

    \I__11614\ : Sp12to4
    port map (
            O => \N__49475\,
            I => \N__49441\
        );

    \I__11613\ : Sp12to4
    port map (
            O => \N__49470\,
            I => \N__49441\
        );

    \I__11612\ : InMux
    port map (
            O => \N__49469\,
            I => \N__49432\
        );

    \I__11611\ : InMux
    port map (
            O => \N__49468\,
            I => \N__49432\
        );

    \I__11610\ : InMux
    port map (
            O => \N__49467\,
            I => \N__49432\
        );

    \I__11609\ : InMux
    port map (
            O => \N__49466\,
            I => \N__49432\
        );

    \I__11608\ : InMux
    port map (
            O => \N__49465\,
            I => \N__49427\
        );

    \I__11607\ : InMux
    port map (
            O => \N__49464\,
            I => \N__49427\
        );

    \I__11606\ : InMux
    port map (
            O => \N__49461\,
            I => \N__49424\
        );

    \I__11605\ : InMux
    port map (
            O => \N__49460\,
            I => \N__49421\
        );

    \I__11604\ : InMux
    port map (
            O => \N__49459\,
            I => \N__49416\
        );

    \I__11603\ : InMux
    port map (
            O => \N__49458\,
            I => \N__49416\
        );

    \I__11602\ : Span4Mux_h
    port map (
            O => \N__49455\,
            I => \N__49411\
        );

    \I__11601\ : Span4Mux_h
    port map (
            O => \N__49452\,
            I => \N__49411\
        );

    \I__11600\ : InMux
    port map (
            O => \N__49451\,
            I => \N__49408\
        );

    \I__11599\ : Sp12to4
    port map (
            O => \N__49446\,
            I => \N__49401\
        );

    \I__11598\ : Span12Mux_v
    port map (
            O => \N__49441\,
            I => \N__49401\
        );

    \I__11597\ : LocalMux
    port map (
            O => \N__49432\,
            I => \N__49401\
        );

    \I__11596\ : LocalMux
    port map (
            O => \N__49427\,
            I => \N__49398\
        );

    \I__11595\ : LocalMux
    port map (
            O => \N__49424\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__11594\ : LocalMux
    port map (
            O => \N__49421\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__11593\ : LocalMux
    port map (
            O => \N__49416\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__11592\ : Odrv4
    port map (
            O => \N__49411\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__11591\ : LocalMux
    port map (
            O => \N__49408\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__11590\ : Odrv12
    port map (
            O => \N__49401\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__11589\ : Odrv4
    port map (
            O => \N__49398\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__11588\ : InMux
    port map (
            O => \N__49383\,
            I => \N__49378\
        );

    \I__11587\ : InMux
    port map (
            O => \N__49382\,
            I => \N__49375\
        );

    \I__11586\ : InMux
    port map (
            O => \N__49381\,
            I => \N__49369\
        );

    \I__11585\ : LocalMux
    port map (
            O => \N__49378\,
            I => \N__49361\
        );

    \I__11584\ : LocalMux
    port map (
            O => \N__49375\,
            I => \N__49358\
        );

    \I__11583\ : InMux
    port map (
            O => \N__49374\,
            I => \N__49351\
        );

    \I__11582\ : InMux
    port map (
            O => \N__49373\,
            I => \N__49351\
        );

    \I__11581\ : InMux
    port map (
            O => \N__49372\,
            I => \N__49351\
        );

    \I__11580\ : LocalMux
    port map (
            O => \N__49369\,
            I => \N__49348\
        );

    \I__11579\ : InMux
    port map (
            O => \N__49368\,
            I => \N__49343\
        );

    \I__11578\ : InMux
    port map (
            O => \N__49367\,
            I => \N__49343\
        );

    \I__11577\ : InMux
    port map (
            O => \N__49366\,
            I => \N__49336\
        );

    \I__11576\ : InMux
    port map (
            O => \N__49365\,
            I => \N__49336\
        );

    \I__11575\ : InMux
    port map (
            O => \N__49364\,
            I => \N__49336\
        );

    \I__11574\ : Span4Mux_v
    port map (
            O => \N__49361\,
            I => \N__49331\
        );

    \I__11573\ : Span4Mux_h
    port map (
            O => \N__49358\,
            I => \N__49331\
        );

    \I__11572\ : LocalMux
    port map (
            O => \N__49351\,
            I => \N__49326\
        );

    \I__11571\ : Span4Mux_h
    port map (
            O => \N__49348\,
            I => \N__49326\
        );

    \I__11570\ : LocalMux
    port map (
            O => \N__49343\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\
        );

    \I__11569\ : LocalMux
    port map (
            O => \N__49336\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\
        );

    \I__11568\ : Odrv4
    port map (
            O => \N__49331\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\
        );

    \I__11567\ : Odrv4
    port map (
            O => \N__49326\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\
        );

    \I__11566\ : InMux
    port map (
            O => \N__49317\,
            I => \N__49312\
        );

    \I__11565\ : InMux
    port map (
            O => \N__49316\,
            I => \N__49309\
        );

    \I__11564\ : InMux
    port map (
            O => \N__49315\,
            I => \N__49306\
        );

    \I__11563\ : LocalMux
    port map (
            O => \N__49312\,
            I => \elapsed_time_ns_1_RNII6NQL1_0_1\
        );

    \I__11562\ : LocalMux
    port map (
            O => \N__49309\,
            I => \elapsed_time_ns_1_RNII6NQL1_0_1\
        );

    \I__11561\ : LocalMux
    port map (
            O => \N__49306\,
            I => \elapsed_time_ns_1_RNII6NQL1_0_1\
        );

    \I__11560\ : CascadeMux
    port map (
            O => \N__49299\,
            I => \N__49295\
        );

    \I__11559\ : InMux
    port map (
            O => \N__49298\,
            I => \N__49292\
        );

    \I__11558\ : InMux
    port map (
            O => \N__49295\,
            I => \N__49289\
        );

    \I__11557\ : LocalMux
    port map (
            O => \N__49292\,
            I => \N__49284\
        );

    \I__11556\ : LocalMux
    port map (
            O => \N__49289\,
            I => \N__49284\
        );

    \I__11555\ : Odrv4
    port map (
            O => \N__49284\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5Z0Z_1\
        );

    \I__11554\ : CascadeMux
    port map (
            O => \N__49281\,
            I => \N__49277\
        );

    \I__11553\ : InMux
    port map (
            O => \N__49280\,
            I => \N__49274\
        );

    \I__11552\ : InMux
    port map (
            O => \N__49277\,
            I => \N__49271\
        );

    \I__11551\ : LocalMux
    port map (
            O => \N__49274\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1\
        );

    \I__11550\ : LocalMux
    port map (
            O => \N__49271\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1\
        );

    \I__11549\ : InMux
    port map (
            O => \N__49266\,
            I => \N__49263\
        );

    \I__11548\ : LocalMux
    port map (
            O => \N__49263\,
            I => \N__49260\
        );

    \I__11547\ : Span4Mux_h
    port map (
            O => \N__49260\,
            I => \N__49257\
        );

    \I__11546\ : Span4Mux_v
    port map (
            O => \N__49257\,
            I => \N__49254\
        );

    \I__11545\ : Odrv4
    port map (
            O => \N__49254\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\
        );

    \I__11544\ : ClkMux
    port map (
            O => \N__49251\,
            I => \N__48825\
        );

    \I__11543\ : ClkMux
    port map (
            O => \N__49250\,
            I => \N__48825\
        );

    \I__11542\ : ClkMux
    port map (
            O => \N__49249\,
            I => \N__48825\
        );

    \I__11541\ : ClkMux
    port map (
            O => \N__49248\,
            I => \N__48825\
        );

    \I__11540\ : ClkMux
    port map (
            O => \N__49247\,
            I => \N__48825\
        );

    \I__11539\ : ClkMux
    port map (
            O => \N__49246\,
            I => \N__48825\
        );

    \I__11538\ : ClkMux
    port map (
            O => \N__49245\,
            I => \N__48825\
        );

    \I__11537\ : ClkMux
    port map (
            O => \N__49244\,
            I => \N__48825\
        );

    \I__11536\ : ClkMux
    port map (
            O => \N__49243\,
            I => \N__48825\
        );

    \I__11535\ : ClkMux
    port map (
            O => \N__49242\,
            I => \N__48825\
        );

    \I__11534\ : ClkMux
    port map (
            O => \N__49241\,
            I => \N__48825\
        );

    \I__11533\ : ClkMux
    port map (
            O => \N__49240\,
            I => \N__48825\
        );

    \I__11532\ : ClkMux
    port map (
            O => \N__49239\,
            I => \N__48825\
        );

    \I__11531\ : ClkMux
    port map (
            O => \N__49238\,
            I => \N__48825\
        );

    \I__11530\ : ClkMux
    port map (
            O => \N__49237\,
            I => \N__48825\
        );

    \I__11529\ : ClkMux
    port map (
            O => \N__49236\,
            I => \N__48825\
        );

    \I__11528\ : ClkMux
    port map (
            O => \N__49235\,
            I => \N__48825\
        );

    \I__11527\ : ClkMux
    port map (
            O => \N__49234\,
            I => \N__48825\
        );

    \I__11526\ : ClkMux
    port map (
            O => \N__49233\,
            I => \N__48825\
        );

    \I__11525\ : ClkMux
    port map (
            O => \N__49232\,
            I => \N__48825\
        );

    \I__11524\ : ClkMux
    port map (
            O => \N__49231\,
            I => \N__48825\
        );

    \I__11523\ : ClkMux
    port map (
            O => \N__49230\,
            I => \N__48825\
        );

    \I__11522\ : ClkMux
    port map (
            O => \N__49229\,
            I => \N__48825\
        );

    \I__11521\ : ClkMux
    port map (
            O => \N__49228\,
            I => \N__48825\
        );

    \I__11520\ : ClkMux
    port map (
            O => \N__49227\,
            I => \N__48825\
        );

    \I__11519\ : ClkMux
    port map (
            O => \N__49226\,
            I => \N__48825\
        );

    \I__11518\ : ClkMux
    port map (
            O => \N__49225\,
            I => \N__48825\
        );

    \I__11517\ : ClkMux
    port map (
            O => \N__49224\,
            I => \N__48825\
        );

    \I__11516\ : ClkMux
    port map (
            O => \N__49223\,
            I => \N__48825\
        );

    \I__11515\ : ClkMux
    port map (
            O => \N__49222\,
            I => \N__48825\
        );

    \I__11514\ : ClkMux
    port map (
            O => \N__49221\,
            I => \N__48825\
        );

    \I__11513\ : ClkMux
    port map (
            O => \N__49220\,
            I => \N__48825\
        );

    \I__11512\ : ClkMux
    port map (
            O => \N__49219\,
            I => \N__48825\
        );

    \I__11511\ : ClkMux
    port map (
            O => \N__49218\,
            I => \N__48825\
        );

    \I__11510\ : ClkMux
    port map (
            O => \N__49217\,
            I => \N__48825\
        );

    \I__11509\ : ClkMux
    port map (
            O => \N__49216\,
            I => \N__48825\
        );

    \I__11508\ : ClkMux
    port map (
            O => \N__49215\,
            I => \N__48825\
        );

    \I__11507\ : ClkMux
    port map (
            O => \N__49214\,
            I => \N__48825\
        );

    \I__11506\ : ClkMux
    port map (
            O => \N__49213\,
            I => \N__48825\
        );

    \I__11505\ : ClkMux
    port map (
            O => \N__49212\,
            I => \N__48825\
        );

    \I__11504\ : ClkMux
    port map (
            O => \N__49211\,
            I => \N__48825\
        );

    \I__11503\ : ClkMux
    port map (
            O => \N__49210\,
            I => \N__48825\
        );

    \I__11502\ : ClkMux
    port map (
            O => \N__49209\,
            I => \N__48825\
        );

    \I__11501\ : ClkMux
    port map (
            O => \N__49208\,
            I => \N__48825\
        );

    \I__11500\ : ClkMux
    port map (
            O => \N__49207\,
            I => \N__48825\
        );

    \I__11499\ : ClkMux
    port map (
            O => \N__49206\,
            I => \N__48825\
        );

    \I__11498\ : ClkMux
    port map (
            O => \N__49205\,
            I => \N__48825\
        );

    \I__11497\ : ClkMux
    port map (
            O => \N__49204\,
            I => \N__48825\
        );

    \I__11496\ : ClkMux
    port map (
            O => \N__49203\,
            I => \N__48825\
        );

    \I__11495\ : ClkMux
    port map (
            O => \N__49202\,
            I => \N__48825\
        );

    \I__11494\ : ClkMux
    port map (
            O => \N__49201\,
            I => \N__48825\
        );

    \I__11493\ : ClkMux
    port map (
            O => \N__49200\,
            I => \N__48825\
        );

    \I__11492\ : ClkMux
    port map (
            O => \N__49199\,
            I => \N__48825\
        );

    \I__11491\ : ClkMux
    port map (
            O => \N__49198\,
            I => \N__48825\
        );

    \I__11490\ : ClkMux
    port map (
            O => \N__49197\,
            I => \N__48825\
        );

    \I__11489\ : ClkMux
    port map (
            O => \N__49196\,
            I => \N__48825\
        );

    \I__11488\ : ClkMux
    port map (
            O => \N__49195\,
            I => \N__48825\
        );

    \I__11487\ : ClkMux
    port map (
            O => \N__49194\,
            I => \N__48825\
        );

    \I__11486\ : ClkMux
    port map (
            O => \N__49193\,
            I => \N__48825\
        );

    \I__11485\ : ClkMux
    port map (
            O => \N__49192\,
            I => \N__48825\
        );

    \I__11484\ : ClkMux
    port map (
            O => \N__49191\,
            I => \N__48825\
        );

    \I__11483\ : ClkMux
    port map (
            O => \N__49190\,
            I => \N__48825\
        );

    \I__11482\ : ClkMux
    port map (
            O => \N__49189\,
            I => \N__48825\
        );

    \I__11481\ : ClkMux
    port map (
            O => \N__49188\,
            I => \N__48825\
        );

    \I__11480\ : ClkMux
    port map (
            O => \N__49187\,
            I => \N__48825\
        );

    \I__11479\ : ClkMux
    port map (
            O => \N__49186\,
            I => \N__48825\
        );

    \I__11478\ : ClkMux
    port map (
            O => \N__49185\,
            I => \N__48825\
        );

    \I__11477\ : ClkMux
    port map (
            O => \N__49184\,
            I => \N__48825\
        );

    \I__11476\ : ClkMux
    port map (
            O => \N__49183\,
            I => \N__48825\
        );

    \I__11475\ : ClkMux
    port map (
            O => \N__49182\,
            I => \N__48825\
        );

    \I__11474\ : ClkMux
    port map (
            O => \N__49181\,
            I => \N__48825\
        );

    \I__11473\ : ClkMux
    port map (
            O => \N__49180\,
            I => \N__48825\
        );

    \I__11472\ : ClkMux
    port map (
            O => \N__49179\,
            I => \N__48825\
        );

    \I__11471\ : ClkMux
    port map (
            O => \N__49178\,
            I => \N__48825\
        );

    \I__11470\ : ClkMux
    port map (
            O => \N__49177\,
            I => \N__48825\
        );

    \I__11469\ : ClkMux
    port map (
            O => \N__49176\,
            I => \N__48825\
        );

    \I__11468\ : ClkMux
    port map (
            O => \N__49175\,
            I => \N__48825\
        );

    \I__11467\ : ClkMux
    port map (
            O => \N__49174\,
            I => \N__48825\
        );

    \I__11466\ : ClkMux
    port map (
            O => \N__49173\,
            I => \N__48825\
        );

    \I__11465\ : ClkMux
    port map (
            O => \N__49172\,
            I => \N__48825\
        );

    \I__11464\ : ClkMux
    port map (
            O => \N__49171\,
            I => \N__48825\
        );

    \I__11463\ : ClkMux
    port map (
            O => \N__49170\,
            I => \N__48825\
        );

    \I__11462\ : ClkMux
    port map (
            O => \N__49169\,
            I => \N__48825\
        );

    \I__11461\ : ClkMux
    port map (
            O => \N__49168\,
            I => \N__48825\
        );

    \I__11460\ : ClkMux
    port map (
            O => \N__49167\,
            I => \N__48825\
        );

    \I__11459\ : ClkMux
    port map (
            O => \N__49166\,
            I => \N__48825\
        );

    \I__11458\ : ClkMux
    port map (
            O => \N__49165\,
            I => \N__48825\
        );

    \I__11457\ : ClkMux
    port map (
            O => \N__49164\,
            I => \N__48825\
        );

    \I__11456\ : ClkMux
    port map (
            O => \N__49163\,
            I => \N__48825\
        );

    \I__11455\ : ClkMux
    port map (
            O => \N__49162\,
            I => \N__48825\
        );

    \I__11454\ : ClkMux
    port map (
            O => \N__49161\,
            I => \N__48825\
        );

    \I__11453\ : ClkMux
    port map (
            O => \N__49160\,
            I => \N__48825\
        );

    \I__11452\ : ClkMux
    port map (
            O => \N__49159\,
            I => \N__48825\
        );

    \I__11451\ : ClkMux
    port map (
            O => \N__49158\,
            I => \N__48825\
        );

    \I__11450\ : ClkMux
    port map (
            O => \N__49157\,
            I => \N__48825\
        );

    \I__11449\ : ClkMux
    port map (
            O => \N__49156\,
            I => \N__48825\
        );

    \I__11448\ : ClkMux
    port map (
            O => \N__49155\,
            I => \N__48825\
        );

    \I__11447\ : ClkMux
    port map (
            O => \N__49154\,
            I => \N__48825\
        );

    \I__11446\ : ClkMux
    port map (
            O => \N__49153\,
            I => \N__48825\
        );

    \I__11445\ : ClkMux
    port map (
            O => \N__49152\,
            I => \N__48825\
        );

    \I__11444\ : ClkMux
    port map (
            O => \N__49151\,
            I => \N__48825\
        );

    \I__11443\ : ClkMux
    port map (
            O => \N__49150\,
            I => \N__48825\
        );

    \I__11442\ : ClkMux
    port map (
            O => \N__49149\,
            I => \N__48825\
        );

    \I__11441\ : ClkMux
    port map (
            O => \N__49148\,
            I => \N__48825\
        );

    \I__11440\ : ClkMux
    port map (
            O => \N__49147\,
            I => \N__48825\
        );

    \I__11439\ : ClkMux
    port map (
            O => \N__49146\,
            I => \N__48825\
        );

    \I__11438\ : ClkMux
    port map (
            O => \N__49145\,
            I => \N__48825\
        );

    \I__11437\ : ClkMux
    port map (
            O => \N__49144\,
            I => \N__48825\
        );

    \I__11436\ : ClkMux
    port map (
            O => \N__49143\,
            I => \N__48825\
        );

    \I__11435\ : ClkMux
    port map (
            O => \N__49142\,
            I => \N__48825\
        );

    \I__11434\ : ClkMux
    port map (
            O => \N__49141\,
            I => \N__48825\
        );

    \I__11433\ : ClkMux
    port map (
            O => \N__49140\,
            I => \N__48825\
        );

    \I__11432\ : ClkMux
    port map (
            O => \N__49139\,
            I => \N__48825\
        );

    \I__11431\ : ClkMux
    port map (
            O => \N__49138\,
            I => \N__48825\
        );

    \I__11430\ : ClkMux
    port map (
            O => \N__49137\,
            I => \N__48825\
        );

    \I__11429\ : ClkMux
    port map (
            O => \N__49136\,
            I => \N__48825\
        );

    \I__11428\ : ClkMux
    port map (
            O => \N__49135\,
            I => \N__48825\
        );

    \I__11427\ : ClkMux
    port map (
            O => \N__49134\,
            I => \N__48825\
        );

    \I__11426\ : ClkMux
    port map (
            O => \N__49133\,
            I => \N__48825\
        );

    \I__11425\ : ClkMux
    port map (
            O => \N__49132\,
            I => \N__48825\
        );

    \I__11424\ : ClkMux
    port map (
            O => \N__49131\,
            I => \N__48825\
        );

    \I__11423\ : ClkMux
    port map (
            O => \N__49130\,
            I => \N__48825\
        );

    \I__11422\ : ClkMux
    port map (
            O => \N__49129\,
            I => \N__48825\
        );

    \I__11421\ : ClkMux
    port map (
            O => \N__49128\,
            I => \N__48825\
        );

    \I__11420\ : ClkMux
    port map (
            O => \N__49127\,
            I => \N__48825\
        );

    \I__11419\ : ClkMux
    port map (
            O => \N__49126\,
            I => \N__48825\
        );

    \I__11418\ : ClkMux
    port map (
            O => \N__49125\,
            I => \N__48825\
        );

    \I__11417\ : ClkMux
    port map (
            O => \N__49124\,
            I => \N__48825\
        );

    \I__11416\ : ClkMux
    port map (
            O => \N__49123\,
            I => \N__48825\
        );

    \I__11415\ : ClkMux
    port map (
            O => \N__49122\,
            I => \N__48825\
        );

    \I__11414\ : ClkMux
    port map (
            O => \N__49121\,
            I => \N__48825\
        );

    \I__11413\ : ClkMux
    port map (
            O => \N__49120\,
            I => \N__48825\
        );

    \I__11412\ : ClkMux
    port map (
            O => \N__49119\,
            I => \N__48825\
        );

    \I__11411\ : ClkMux
    port map (
            O => \N__49118\,
            I => \N__48825\
        );

    \I__11410\ : ClkMux
    port map (
            O => \N__49117\,
            I => \N__48825\
        );

    \I__11409\ : ClkMux
    port map (
            O => \N__49116\,
            I => \N__48825\
        );

    \I__11408\ : ClkMux
    port map (
            O => \N__49115\,
            I => \N__48825\
        );

    \I__11407\ : ClkMux
    port map (
            O => \N__49114\,
            I => \N__48825\
        );

    \I__11406\ : ClkMux
    port map (
            O => \N__49113\,
            I => \N__48825\
        );

    \I__11405\ : ClkMux
    port map (
            O => \N__49112\,
            I => \N__48825\
        );

    \I__11404\ : ClkMux
    port map (
            O => \N__49111\,
            I => \N__48825\
        );

    \I__11403\ : ClkMux
    port map (
            O => \N__49110\,
            I => \N__48825\
        );

    \I__11402\ : GlobalMux
    port map (
            O => \N__48825\,
            I => clk_100mhz_0
        );

    \I__11401\ : CEMux
    port map (
            O => \N__48822\,
            I => \N__48816\
        );

    \I__11400\ : CEMux
    port map (
            O => \N__48821\,
            I => \N__48808\
        );

    \I__11399\ : CEMux
    port map (
            O => \N__48820\,
            I => \N__48798\
        );

    \I__11398\ : CEMux
    port map (
            O => \N__48819\,
            I => \N__48795\
        );

    \I__11397\ : LocalMux
    port map (
            O => \N__48816\,
            I => \N__48792\
        );

    \I__11396\ : InMux
    port map (
            O => \N__48815\,
            I => \N__48783\
        );

    \I__11395\ : InMux
    port map (
            O => \N__48814\,
            I => \N__48783\
        );

    \I__11394\ : InMux
    port map (
            O => \N__48813\,
            I => \N__48783\
        );

    \I__11393\ : InMux
    port map (
            O => \N__48812\,
            I => \N__48783\
        );

    \I__11392\ : CEMux
    port map (
            O => \N__48811\,
            I => \N__48780\
        );

    \I__11391\ : LocalMux
    port map (
            O => \N__48808\,
            I => \N__48777\
        );

    \I__11390\ : InMux
    port map (
            O => \N__48807\,
            I => \N__48770\
        );

    \I__11389\ : InMux
    port map (
            O => \N__48806\,
            I => \N__48770\
        );

    \I__11388\ : InMux
    port map (
            O => \N__48805\,
            I => \N__48770\
        );

    \I__11387\ : CEMux
    port map (
            O => \N__48804\,
            I => \N__48767\
        );

    \I__11386\ : CEMux
    port map (
            O => \N__48803\,
            I => \N__48764\
        );

    \I__11385\ : CEMux
    port map (
            O => \N__48802\,
            I => \N__48742\
        );

    \I__11384\ : CEMux
    port map (
            O => \N__48801\,
            I => \N__48739\
        );

    \I__11383\ : LocalMux
    port map (
            O => \N__48798\,
            I => \N__48736\
        );

    \I__11382\ : LocalMux
    port map (
            O => \N__48795\,
            I => \N__48733\
        );

    \I__11381\ : Span4Mux_h
    port map (
            O => \N__48792\,
            I => \N__48730\
        );

    \I__11380\ : LocalMux
    port map (
            O => \N__48783\,
            I => \N__48727\
        );

    \I__11379\ : LocalMux
    port map (
            O => \N__48780\,
            I => \N__48722\
        );

    \I__11378\ : Span4Mux_v
    port map (
            O => \N__48777\,
            I => \N__48722\
        );

    \I__11377\ : LocalMux
    port map (
            O => \N__48770\,
            I => \N__48717\
        );

    \I__11376\ : LocalMux
    port map (
            O => \N__48767\,
            I => \N__48717\
        );

    \I__11375\ : LocalMux
    port map (
            O => \N__48764\,
            I => \N__48714\
        );

    \I__11374\ : InMux
    port map (
            O => \N__48763\,
            I => \N__48705\
        );

    \I__11373\ : InMux
    port map (
            O => \N__48762\,
            I => \N__48705\
        );

    \I__11372\ : InMux
    port map (
            O => \N__48761\,
            I => \N__48705\
        );

    \I__11371\ : InMux
    port map (
            O => \N__48760\,
            I => \N__48705\
        );

    \I__11370\ : InMux
    port map (
            O => \N__48759\,
            I => \N__48696\
        );

    \I__11369\ : InMux
    port map (
            O => \N__48758\,
            I => \N__48696\
        );

    \I__11368\ : InMux
    port map (
            O => \N__48757\,
            I => \N__48696\
        );

    \I__11367\ : InMux
    port map (
            O => \N__48756\,
            I => \N__48696\
        );

    \I__11366\ : InMux
    port map (
            O => \N__48755\,
            I => \N__48689\
        );

    \I__11365\ : InMux
    port map (
            O => \N__48754\,
            I => \N__48689\
        );

    \I__11364\ : InMux
    port map (
            O => \N__48753\,
            I => \N__48689\
        );

    \I__11363\ : InMux
    port map (
            O => \N__48752\,
            I => \N__48680\
        );

    \I__11362\ : InMux
    port map (
            O => \N__48751\,
            I => \N__48680\
        );

    \I__11361\ : InMux
    port map (
            O => \N__48750\,
            I => \N__48680\
        );

    \I__11360\ : InMux
    port map (
            O => \N__48749\,
            I => \N__48680\
        );

    \I__11359\ : InMux
    port map (
            O => \N__48748\,
            I => \N__48671\
        );

    \I__11358\ : InMux
    port map (
            O => \N__48747\,
            I => \N__48671\
        );

    \I__11357\ : InMux
    port map (
            O => \N__48746\,
            I => \N__48671\
        );

    \I__11356\ : InMux
    port map (
            O => \N__48745\,
            I => \N__48671\
        );

    \I__11355\ : LocalMux
    port map (
            O => \N__48742\,
            I => \N__48663\
        );

    \I__11354\ : LocalMux
    port map (
            O => \N__48739\,
            I => \N__48660\
        );

    \I__11353\ : Span4Mux_v
    port map (
            O => \N__48736\,
            I => \N__48655\
        );

    \I__11352\ : Span4Mux_v
    port map (
            O => \N__48733\,
            I => \N__48655\
        );

    \I__11351\ : Span4Mux_v
    port map (
            O => \N__48730\,
            I => \N__48652\
        );

    \I__11350\ : Span4Mux_v
    port map (
            O => \N__48727\,
            I => \N__48645\
        );

    \I__11349\ : Span4Mux_v
    port map (
            O => \N__48722\,
            I => \N__48645\
        );

    \I__11348\ : Span4Mux_v
    port map (
            O => \N__48717\,
            I => \N__48645\
        );

    \I__11347\ : Span4Mux_v
    port map (
            O => \N__48714\,
            I => \N__48638\
        );

    \I__11346\ : LocalMux
    port map (
            O => \N__48705\,
            I => \N__48638\
        );

    \I__11345\ : LocalMux
    port map (
            O => \N__48696\,
            I => \N__48638\
        );

    \I__11344\ : LocalMux
    port map (
            O => \N__48689\,
            I => \N__48631\
        );

    \I__11343\ : LocalMux
    port map (
            O => \N__48680\,
            I => \N__48631\
        );

    \I__11342\ : LocalMux
    port map (
            O => \N__48671\,
            I => \N__48631\
        );

    \I__11341\ : InMux
    port map (
            O => \N__48670\,
            I => \N__48622\
        );

    \I__11340\ : InMux
    port map (
            O => \N__48669\,
            I => \N__48622\
        );

    \I__11339\ : InMux
    port map (
            O => \N__48668\,
            I => \N__48622\
        );

    \I__11338\ : InMux
    port map (
            O => \N__48667\,
            I => \N__48622\
        );

    \I__11337\ : InMux
    port map (
            O => \N__48666\,
            I => \N__48619\
        );

    \I__11336\ : Sp12to4
    port map (
            O => \N__48663\,
            I => \N__48616\
        );

    \I__11335\ : Span4Mux_v
    port map (
            O => \N__48660\,
            I => \N__48611\
        );

    \I__11334\ : Span4Mux_v
    port map (
            O => \N__48655\,
            I => \N__48611\
        );

    \I__11333\ : Span4Mux_h
    port map (
            O => \N__48652\,
            I => \N__48602\
        );

    \I__11332\ : Span4Mux_h
    port map (
            O => \N__48645\,
            I => \N__48602\
        );

    \I__11331\ : Span4Mux_v
    port map (
            O => \N__48638\,
            I => \N__48602\
        );

    \I__11330\ : Span4Mux_v
    port map (
            O => \N__48631\,
            I => \N__48602\
        );

    \I__11329\ : LocalMux
    port map (
            O => \N__48622\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__11328\ : LocalMux
    port map (
            O => \N__48619\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__11327\ : Odrv12
    port map (
            O => \N__48616\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__11326\ : Odrv4
    port map (
            O => \N__48611\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__11325\ : Odrv4
    port map (
            O => \N__48602\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__11324\ : InMux
    port map (
            O => \N__48591\,
            I => \N__48580\
        );

    \I__11323\ : InMux
    port map (
            O => \N__48590\,
            I => \N__48577\
        );

    \I__11322\ : InMux
    port map (
            O => \N__48589\,
            I => \N__48574\
        );

    \I__11321\ : InMux
    port map (
            O => \N__48588\,
            I => \N__48571\
        );

    \I__11320\ : InMux
    port map (
            O => \N__48587\,
            I => \N__48568\
        );

    \I__11319\ : InMux
    port map (
            O => \N__48586\,
            I => \N__48565\
        );

    \I__11318\ : InMux
    port map (
            O => \N__48585\,
            I => \N__48562\
        );

    \I__11317\ : InMux
    port map (
            O => \N__48584\,
            I => \N__48559\
        );

    \I__11316\ : InMux
    port map (
            O => \N__48583\,
            I => \N__48556\
        );

    \I__11315\ : LocalMux
    port map (
            O => \N__48580\,
            I => \N__48553\
        );

    \I__11314\ : LocalMux
    port map (
            O => \N__48577\,
            I => \N__48550\
        );

    \I__11313\ : LocalMux
    port map (
            O => \N__48574\,
            I => \N__48547\
        );

    \I__11312\ : LocalMux
    port map (
            O => \N__48571\,
            I => \N__48501\
        );

    \I__11311\ : LocalMux
    port map (
            O => \N__48568\,
            I => \N__48489\
        );

    \I__11310\ : LocalMux
    port map (
            O => \N__48565\,
            I => \N__48450\
        );

    \I__11309\ : LocalMux
    port map (
            O => \N__48562\,
            I => \N__48438\
        );

    \I__11308\ : LocalMux
    port map (
            O => \N__48559\,
            I => \N__48423\
        );

    \I__11307\ : LocalMux
    port map (
            O => \N__48556\,
            I => \N__48409\
        );

    \I__11306\ : Glb2LocalMux
    port map (
            O => \N__48553\,
            I => \N__48096\
        );

    \I__11305\ : Glb2LocalMux
    port map (
            O => \N__48550\,
            I => \N__48096\
        );

    \I__11304\ : Glb2LocalMux
    port map (
            O => \N__48547\,
            I => \N__48096\
        );

    \I__11303\ : SRMux
    port map (
            O => \N__48546\,
            I => \N__48096\
        );

    \I__11302\ : SRMux
    port map (
            O => \N__48545\,
            I => \N__48096\
        );

    \I__11301\ : SRMux
    port map (
            O => \N__48544\,
            I => \N__48096\
        );

    \I__11300\ : SRMux
    port map (
            O => \N__48543\,
            I => \N__48096\
        );

    \I__11299\ : SRMux
    port map (
            O => \N__48542\,
            I => \N__48096\
        );

    \I__11298\ : SRMux
    port map (
            O => \N__48541\,
            I => \N__48096\
        );

    \I__11297\ : SRMux
    port map (
            O => \N__48540\,
            I => \N__48096\
        );

    \I__11296\ : SRMux
    port map (
            O => \N__48539\,
            I => \N__48096\
        );

    \I__11295\ : SRMux
    port map (
            O => \N__48538\,
            I => \N__48096\
        );

    \I__11294\ : SRMux
    port map (
            O => \N__48537\,
            I => \N__48096\
        );

    \I__11293\ : SRMux
    port map (
            O => \N__48536\,
            I => \N__48096\
        );

    \I__11292\ : SRMux
    port map (
            O => \N__48535\,
            I => \N__48096\
        );

    \I__11291\ : SRMux
    port map (
            O => \N__48534\,
            I => \N__48096\
        );

    \I__11290\ : SRMux
    port map (
            O => \N__48533\,
            I => \N__48096\
        );

    \I__11289\ : SRMux
    port map (
            O => \N__48532\,
            I => \N__48096\
        );

    \I__11288\ : SRMux
    port map (
            O => \N__48531\,
            I => \N__48096\
        );

    \I__11287\ : SRMux
    port map (
            O => \N__48530\,
            I => \N__48096\
        );

    \I__11286\ : SRMux
    port map (
            O => \N__48529\,
            I => \N__48096\
        );

    \I__11285\ : SRMux
    port map (
            O => \N__48528\,
            I => \N__48096\
        );

    \I__11284\ : SRMux
    port map (
            O => \N__48527\,
            I => \N__48096\
        );

    \I__11283\ : SRMux
    port map (
            O => \N__48526\,
            I => \N__48096\
        );

    \I__11282\ : SRMux
    port map (
            O => \N__48525\,
            I => \N__48096\
        );

    \I__11281\ : SRMux
    port map (
            O => \N__48524\,
            I => \N__48096\
        );

    \I__11280\ : SRMux
    port map (
            O => \N__48523\,
            I => \N__48096\
        );

    \I__11279\ : SRMux
    port map (
            O => \N__48522\,
            I => \N__48096\
        );

    \I__11278\ : SRMux
    port map (
            O => \N__48521\,
            I => \N__48096\
        );

    \I__11277\ : SRMux
    port map (
            O => \N__48520\,
            I => \N__48096\
        );

    \I__11276\ : SRMux
    port map (
            O => \N__48519\,
            I => \N__48096\
        );

    \I__11275\ : SRMux
    port map (
            O => \N__48518\,
            I => \N__48096\
        );

    \I__11274\ : SRMux
    port map (
            O => \N__48517\,
            I => \N__48096\
        );

    \I__11273\ : SRMux
    port map (
            O => \N__48516\,
            I => \N__48096\
        );

    \I__11272\ : SRMux
    port map (
            O => \N__48515\,
            I => \N__48096\
        );

    \I__11271\ : SRMux
    port map (
            O => \N__48514\,
            I => \N__48096\
        );

    \I__11270\ : SRMux
    port map (
            O => \N__48513\,
            I => \N__48096\
        );

    \I__11269\ : SRMux
    port map (
            O => \N__48512\,
            I => \N__48096\
        );

    \I__11268\ : SRMux
    port map (
            O => \N__48511\,
            I => \N__48096\
        );

    \I__11267\ : SRMux
    port map (
            O => \N__48510\,
            I => \N__48096\
        );

    \I__11266\ : SRMux
    port map (
            O => \N__48509\,
            I => \N__48096\
        );

    \I__11265\ : SRMux
    port map (
            O => \N__48508\,
            I => \N__48096\
        );

    \I__11264\ : SRMux
    port map (
            O => \N__48507\,
            I => \N__48096\
        );

    \I__11263\ : SRMux
    port map (
            O => \N__48506\,
            I => \N__48096\
        );

    \I__11262\ : SRMux
    port map (
            O => \N__48505\,
            I => \N__48096\
        );

    \I__11261\ : SRMux
    port map (
            O => \N__48504\,
            I => \N__48096\
        );

    \I__11260\ : Glb2LocalMux
    port map (
            O => \N__48501\,
            I => \N__48096\
        );

    \I__11259\ : SRMux
    port map (
            O => \N__48500\,
            I => \N__48096\
        );

    \I__11258\ : SRMux
    port map (
            O => \N__48499\,
            I => \N__48096\
        );

    \I__11257\ : SRMux
    port map (
            O => \N__48498\,
            I => \N__48096\
        );

    \I__11256\ : SRMux
    port map (
            O => \N__48497\,
            I => \N__48096\
        );

    \I__11255\ : SRMux
    port map (
            O => \N__48496\,
            I => \N__48096\
        );

    \I__11254\ : SRMux
    port map (
            O => \N__48495\,
            I => \N__48096\
        );

    \I__11253\ : SRMux
    port map (
            O => \N__48494\,
            I => \N__48096\
        );

    \I__11252\ : SRMux
    port map (
            O => \N__48493\,
            I => \N__48096\
        );

    \I__11251\ : SRMux
    port map (
            O => \N__48492\,
            I => \N__48096\
        );

    \I__11250\ : Glb2LocalMux
    port map (
            O => \N__48489\,
            I => \N__48096\
        );

    \I__11249\ : SRMux
    port map (
            O => \N__48488\,
            I => \N__48096\
        );

    \I__11248\ : SRMux
    port map (
            O => \N__48487\,
            I => \N__48096\
        );

    \I__11247\ : SRMux
    port map (
            O => \N__48486\,
            I => \N__48096\
        );

    \I__11246\ : SRMux
    port map (
            O => \N__48485\,
            I => \N__48096\
        );

    \I__11245\ : SRMux
    port map (
            O => \N__48484\,
            I => \N__48096\
        );

    \I__11244\ : SRMux
    port map (
            O => \N__48483\,
            I => \N__48096\
        );

    \I__11243\ : SRMux
    port map (
            O => \N__48482\,
            I => \N__48096\
        );

    \I__11242\ : SRMux
    port map (
            O => \N__48481\,
            I => \N__48096\
        );

    \I__11241\ : SRMux
    port map (
            O => \N__48480\,
            I => \N__48096\
        );

    \I__11240\ : SRMux
    port map (
            O => \N__48479\,
            I => \N__48096\
        );

    \I__11239\ : SRMux
    port map (
            O => \N__48478\,
            I => \N__48096\
        );

    \I__11238\ : SRMux
    port map (
            O => \N__48477\,
            I => \N__48096\
        );

    \I__11237\ : SRMux
    port map (
            O => \N__48476\,
            I => \N__48096\
        );

    \I__11236\ : SRMux
    port map (
            O => \N__48475\,
            I => \N__48096\
        );

    \I__11235\ : SRMux
    port map (
            O => \N__48474\,
            I => \N__48096\
        );

    \I__11234\ : SRMux
    port map (
            O => \N__48473\,
            I => \N__48096\
        );

    \I__11233\ : SRMux
    port map (
            O => \N__48472\,
            I => \N__48096\
        );

    \I__11232\ : SRMux
    port map (
            O => \N__48471\,
            I => \N__48096\
        );

    \I__11231\ : SRMux
    port map (
            O => \N__48470\,
            I => \N__48096\
        );

    \I__11230\ : SRMux
    port map (
            O => \N__48469\,
            I => \N__48096\
        );

    \I__11229\ : SRMux
    port map (
            O => \N__48468\,
            I => \N__48096\
        );

    \I__11228\ : SRMux
    port map (
            O => \N__48467\,
            I => \N__48096\
        );

    \I__11227\ : SRMux
    port map (
            O => \N__48466\,
            I => \N__48096\
        );

    \I__11226\ : SRMux
    port map (
            O => \N__48465\,
            I => \N__48096\
        );

    \I__11225\ : SRMux
    port map (
            O => \N__48464\,
            I => \N__48096\
        );

    \I__11224\ : SRMux
    port map (
            O => \N__48463\,
            I => \N__48096\
        );

    \I__11223\ : SRMux
    port map (
            O => \N__48462\,
            I => \N__48096\
        );

    \I__11222\ : SRMux
    port map (
            O => \N__48461\,
            I => \N__48096\
        );

    \I__11221\ : SRMux
    port map (
            O => \N__48460\,
            I => \N__48096\
        );

    \I__11220\ : SRMux
    port map (
            O => \N__48459\,
            I => \N__48096\
        );

    \I__11219\ : SRMux
    port map (
            O => \N__48458\,
            I => \N__48096\
        );

    \I__11218\ : SRMux
    port map (
            O => \N__48457\,
            I => \N__48096\
        );

    \I__11217\ : SRMux
    port map (
            O => \N__48456\,
            I => \N__48096\
        );

    \I__11216\ : SRMux
    port map (
            O => \N__48455\,
            I => \N__48096\
        );

    \I__11215\ : SRMux
    port map (
            O => \N__48454\,
            I => \N__48096\
        );

    \I__11214\ : SRMux
    port map (
            O => \N__48453\,
            I => \N__48096\
        );

    \I__11213\ : Glb2LocalMux
    port map (
            O => \N__48450\,
            I => \N__48096\
        );

    \I__11212\ : SRMux
    port map (
            O => \N__48449\,
            I => \N__48096\
        );

    \I__11211\ : SRMux
    port map (
            O => \N__48448\,
            I => \N__48096\
        );

    \I__11210\ : SRMux
    port map (
            O => \N__48447\,
            I => \N__48096\
        );

    \I__11209\ : SRMux
    port map (
            O => \N__48446\,
            I => \N__48096\
        );

    \I__11208\ : SRMux
    port map (
            O => \N__48445\,
            I => \N__48096\
        );

    \I__11207\ : SRMux
    port map (
            O => \N__48444\,
            I => \N__48096\
        );

    \I__11206\ : SRMux
    port map (
            O => \N__48443\,
            I => \N__48096\
        );

    \I__11205\ : SRMux
    port map (
            O => \N__48442\,
            I => \N__48096\
        );

    \I__11204\ : SRMux
    port map (
            O => \N__48441\,
            I => \N__48096\
        );

    \I__11203\ : Glb2LocalMux
    port map (
            O => \N__48438\,
            I => \N__48096\
        );

    \I__11202\ : SRMux
    port map (
            O => \N__48437\,
            I => \N__48096\
        );

    \I__11201\ : SRMux
    port map (
            O => \N__48436\,
            I => \N__48096\
        );

    \I__11200\ : SRMux
    port map (
            O => \N__48435\,
            I => \N__48096\
        );

    \I__11199\ : SRMux
    port map (
            O => \N__48434\,
            I => \N__48096\
        );

    \I__11198\ : SRMux
    port map (
            O => \N__48433\,
            I => \N__48096\
        );

    \I__11197\ : SRMux
    port map (
            O => \N__48432\,
            I => \N__48096\
        );

    \I__11196\ : SRMux
    port map (
            O => \N__48431\,
            I => \N__48096\
        );

    \I__11195\ : SRMux
    port map (
            O => \N__48430\,
            I => \N__48096\
        );

    \I__11194\ : SRMux
    port map (
            O => \N__48429\,
            I => \N__48096\
        );

    \I__11193\ : SRMux
    port map (
            O => \N__48428\,
            I => \N__48096\
        );

    \I__11192\ : SRMux
    port map (
            O => \N__48427\,
            I => \N__48096\
        );

    \I__11191\ : SRMux
    port map (
            O => \N__48426\,
            I => \N__48096\
        );

    \I__11190\ : Glb2LocalMux
    port map (
            O => \N__48423\,
            I => \N__48096\
        );

    \I__11189\ : SRMux
    port map (
            O => \N__48422\,
            I => \N__48096\
        );

    \I__11188\ : SRMux
    port map (
            O => \N__48421\,
            I => \N__48096\
        );

    \I__11187\ : SRMux
    port map (
            O => \N__48420\,
            I => \N__48096\
        );

    \I__11186\ : SRMux
    port map (
            O => \N__48419\,
            I => \N__48096\
        );

    \I__11185\ : SRMux
    port map (
            O => \N__48418\,
            I => \N__48096\
        );

    \I__11184\ : SRMux
    port map (
            O => \N__48417\,
            I => \N__48096\
        );

    \I__11183\ : SRMux
    port map (
            O => \N__48416\,
            I => \N__48096\
        );

    \I__11182\ : SRMux
    port map (
            O => \N__48415\,
            I => \N__48096\
        );

    \I__11181\ : SRMux
    port map (
            O => \N__48414\,
            I => \N__48096\
        );

    \I__11180\ : SRMux
    port map (
            O => \N__48413\,
            I => \N__48096\
        );

    \I__11179\ : SRMux
    port map (
            O => \N__48412\,
            I => \N__48096\
        );

    \I__11178\ : Glb2LocalMux
    port map (
            O => \N__48409\,
            I => \N__48096\
        );

    \I__11177\ : SRMux
    port map (
            O => \N__48408\,
            I => \N__48096\
        );

    \I__11176\ : SRMux
    port map (
            O => \N__48407\,
            I => \N__48096\
        );

    \I__11175\ : SRMux
    port map (
            O => \N__48406\,
            I => \N__48096\
        );

    \I__11174\ : SRMux
    port map (
            O => \N__48405\,
            I => \N__48096\
        );

    \I__11173\ : SRMux
    port map (
            O => \N__48404\,
            I => \N__48096\
        );

    \I__11172\ : SRMux
    port map (
            O => \N__48403\,
            I => \N__48096\
        );

    \I__11171\ : SRMux
    port map (
            O => \N__48402\,
            I => \N__48096\
        );

    \I__11170\ : SRMux
    port map (
            O => \N__48401\,
            I => \N__48096\
        );

    \I__11169\ : SRMux
    port map (
            O => \N__48400\,
            I => \N__48096\
        );

    \I__11168\ : SRMux
    port map (
            O => \N__48399\,
            I => \N__48096\
        );

    \I__11167\ : SRMux
    port map (
            O => \N__48398\,
            I => \N__48096\
        );

    \I__11166\ : SRMux
    port map (
            O => \N__48397\,
            I => \N__48096\
        );

    \I__11165\ : SRMux
    port map (
            O => \N__48396\,
            I => \N__48096\
        );

    \I__11164\ : SRMux
    port map (
            O => \N__48395\,
            I => \N__48096\
        );

    \I__11163\ : SRMux
    port map (
            O => \N__48394\,
            I => \N__48096\
        );

    \I__11162\ : SRMux
    port map (
            O => \N__48393\,
            I => \N__48096\
        );

    \I__11161\ : SRMux
    port map (
            O => \N__48392\,
            I => \N__48096\
        );

    \I__11160\ : SRMux
    port map (
            O => \N__48391\,
            I => \N__48096\
        );

    \I__11159\ : GlobalMux
    port map (
            O => \N__48096\,
            I => \N__48093\
        );

    \I__11158\ : gio2CtrlBuf
    port map (
            O => \N__48093\,
            I => red_c_g
        );

    \I__11157\ : InMux
    port map (
            O => \N__48090\,
            I => \N__48052\
        );

    \I__11156\ : InMux
    port map (
            O => \N__48089\,
            I => \N__48052\
        );

    \I__11155\ : InMux
    port map (
            O => \N__48088\,
            I => \N__48052\
        );

    \I__11154\ : InMux
    port map (
            O => \N__48087\,
            I => \N__48052\
        );

    \I__11153\ : InMux
    port map (
            O => \N__48086\,
            I => \N__48043\
        );

    \I__11152\ : InMux
    port map (
            O => \N__48085\,
            I => \N__48043\
        );

    \I__11151\ : InMux
    port map (
            O => \N__48084\,
            I => \N__48043\
        );

    \I__11150\ : InMux
    port map (
            O => \N__48083\,
            I => \N__48043\
        );

    \I__11149\ : InMux
    port map (
            O => \N__48082\,
            I => \N__48038\
        );

    \I__11148\ : InMux
    port map (
            O => \N__48081\,
            I => \N__48038\
        );

    \I__11147\ : InMux
    port map (
            O => \N__48080\,
            I => \N__48029\
        );

    \I__11146\ : InMux
    port map (
            O => \N__48079\,
            I => \N__48029\
        );

    \I__11145\ : InMux
    port map (
            O => \N__48078\,
            I => \N__48029\
        );

    \I__11144\ : InMux
    port map (
            O => \N__48077\,
            I => \N__48029\
        );

    \I__11143\ : InMux
    port map (
            O => \N__48076\,
            I => \N__48020\
        );

    \I__11142\ : InMux
    port map (
            O => \N__48075\,
            I => \N__48020\
        );

    \I__11141\ : InMux
    port map (
            O => \N__48074\,
            I => \N__48020\
        );

    \I__11140\ : InMux
    port map (
            O => \N__48073\,
            I => \N__48020\
        );

    \I__11139\ : InMux
    port map (
            O => \N__48072\,
            I => \N__48011\
        );

    \I__11138\ : InMux
    port map (
            O => \N__48071\,
            I => \N__48011\
        );

    \I__11137\ : InMux
    port map (
            O => \N__48070\,
            I => \N__48011\
        );

    \I__11136\ : InMux
    port map (
            O => \N__48069\,
            I => \N__48011\
        );

    \I__11135\ : InMux
    port map (
            O => \N__48068\,
            I => \N__48002\
        );

    \I__11134\ : InMux
    port map (
            O => \N__48067\,
            I => \N__48002\
        );

    \I__11133\ : InMux
    port map (
            O => \N__48066\,
            I => \N__48002\
        );

    \I__11132\ : InMux
    port map (
            O => \N__48065\,
            I => \N__48002\
        );

    \I__11131\ : InMux
    port map (
            O => \N__48064\,
            I => \N__47993\
        );

    \I__11130\ : InMux
    port map (
            O => \N__48063\,
            I => \N__47993\
        );

    \I__11129\ : InMux
    port map (
            O => \N__48062\,
            I => \N__47993\
        );

    \I__11128\ : InMux
    port map (
            O => \N__48061\,
            I => \N__47993\
        );

    \I__11127\ : LocalMux
    port map (
            O => \N__48052\,
            I => \N__47990\
        );

    \I__11126\ : LocalMux
    port map (
            O => \N__48043\,
            I => \N__47987\
        );

    \I__11125\ : LocalMux
    port map (
            O => \N__48038\,
            I => \N__47974\
        );

    \I__11124\ : LocalMux
    port map (
            O => \N__48029\,
            I => \N__47974\
        );

    \I__11123\ : LocalMux
    port map (
            O => \N__48020\,
            I => \N__47974\
        );

    \I__11122\ : LocalMux
    port map (
            O => \N__48011\,
            I => \N__47974\
        );

    \I__11121\ : LocalMux
    port map (
            O => \N__48002\,
            I => \N__47974\
        );

    \I__11120\ : LocalMux
    port map (
            O => \N__47993\,
            I => \N__47974\
        );

    \I__11119\ : Span4Mux_h
    port map (
            O => \N__47990\,
            I => \N__47971\
        );

    \I__11118\ : Span4Mux_v
    port map (
            O => \N__47987\,
            I => \N__47966\
        );

    \I__11117\ : Span4Mux_v
    port map (
            O => \N__47974\,
            I => \N__47966\
        );

    \I__11116\ : Odrv4
    port map (
            O => \N__47971\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__11115\ : Odrv4
    port map (
            O => \N__47966\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__11114\ : InMux
    port map (
            O => \N__47961\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__11113\ : InMux
    port map (
            O => \N__47958\,
            I => \N__47954\
        );

    \I__11112\ : InMux
    port map (
            O => \N__47957\,
            I => \N__47951\
        );

    \I__11111\ : LocalMux
    port map (
            O => \N__47954\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__11110\ : LocalMux
    port map (
            O => \N__47951\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__11109\ : CEMux
    port map (
            O => \N__47946\,
            I => \N__47941\
        );

    \I__11108\ : CEMux
    port map (
            O => \N__47945\,
            I => \N__47938\
        );

    \I__11107\ : CEMux
    port map (
            O => \N__47944\,
            I => \N__47935\
        );

    \I__11106\ : LocalMux
    port map (
            O => \N__47941\,
            I => \N__47929\
        );

    \I__11105\ : LocalMux
    port map (
            O => \N__47938\,
            I => \N__47929\
        );

    \I__11104\ : LocalMux
    port map (
            O => \N__47935\,
            I => \N__47926\
        );

    \I__11103\ : CEMux
    port map (
            O => \N__47934\,
            I => \N__47923\
        );

    \I__11102\ : Span4Mux_v
    port map (
            O => \N__47929\,
            I => \N__47920\
        );

    \I__11101\ : Span4Mux_v
    port map (
            O => \N__47926\,
            I => \N__47915\
        );

    \I__11100\ : LocalMux
    port map (
            O => \N__47923\,
            I => \N__47915\
        );

    \I__11099\ : Span4Mux_h
    port map (
            O => \N__47920\,
            I => \N__47910\
        );

    \I__11098\ : Span4Mux_h
    port map (
            O => \N__47915\,
            I => \N__47910\
        );

    \I__11097\ : Odrv4
    port map (
            O => \N__47910\,
            I => \delay_measurement_inst.delay_tr_timer.N_396_i\
        );

    \I__11096\ : CascadeMux
    port map (
            O => \N__47907\,
            I => \N__47904\
        );

    \I__11095\ : InMux
    port map (
            O => \N__47904\,
            I => \N__47901\
        );

    \I__11094\ : LocalMux
    port map (
            O => \N__47901\,
            I => \N__47898\
        );

    \I__11093\ : Span12Mux_v
    port map (
            O => \N__47898\,
            I => \N__47894\
        );

    \I__11092\ : InMux
    port map (
            O => \N__47897\,
            I => \N__47891\
        );

    \I__11091\ : Odrv12
    port map (
            O => \N__47894\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__11090\ : LocalMux
    port map (
            O => \N__47891\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__11089\ : InMux
    port map (
            O => \N__47886\,
            I => \N__47882\
        );

    \I__11088\ : InMux
    port map (
            O => \N__47885\,
            I => \N__47878\
        );

    \I__11087\ : LocalMux
    port map (
            O => \N__47882\,
            I => \N__47875\
        );

    \I__11086\ : InMux
    port map (
            O => \N__47881\,
            I => \N__47872\
        );

    \I__11085\ : LocalMux
    port map (
            O => \N__47878\,
            I => \N__47868\
        );

    \I__11084\ : Span4Mux_v
    port map (
            O => \N__47875\,
            I => \N__47863\
        );

    \I__11083\ : LocalMux
    port map (
            O => \N__47872\,
            I => \N__47863\
        );

    \I__11082\ : InMux
    port map (
            O => \N__47871\,
            I => \N__47860\
        );

    \I__11081\ : Span4Mux_h
    port map (
            O => \N__47868\,
            I => \N__47857\
        );

    \I__11080\ : Span4Mux_h
    port map (
            O => \N__47863\,
            I => \N__47854\
        );

    \I__11079\ : LocalMux
    port map (
            O => \N__47860\,
            I => \elapsed_time_ns_1_RNIGK2591_0_8\
        );

    \I__11078\ : Odrv4
    port map (
            O => \N__47857\,
            I => \elapsed_time_ns_1_RNIGK2591_0_8\
        );

    \I__11077\ : Odrv4
    port map (
            O => \N__47854\,
            I => \elapsed_time_ns_1_RNIGK2591_0_8\
        );

    \I__11076\ : InMux
    port map (
            O => \N__47847\,
            I => \N__47843\
        );

    \I__11075\ : InMux
    port map (
            O => \N__47846\,
            I => \N__47838\
        );

    \I__11074\ : LocalMux
    port map (
            O => \N__47843\,
            I => \N__47835\
        );

    \I__11073\ : InMux
    port map (
            O => \N__47842\,
            I => \N__47832\
        );

    \I__11072\ : InMux
    port map (
            O => \N__47841\,
            I => \N__47829\
        );

    \I__11071\ : LocalMux
    port map (
            O => \N__47838\,
            I => \N__47823\
        );

    \I__11070\ : Span4Mux_v
    port map (
            O => \N__47835\,
            I => \N__47819\
        );

    \I__11069\ : LocalMux
    port map (
            O => \N__47832\,
            I => \N__47814\
        );

    \I__11068\ : LocalMux
    port map (
            O => \N__47829\,
            I => \N__47814\
        );

    \I__11067\ : InMux
    port map (
            O => \N__47828\,
            I => \N__47807\
        );

    \I__11066\ : InMux
    port map (
            O => \N__47827\,
            I => \N__47807\
        );

    \I__11065\ : InMux
    port map (
            O => \N__47826\,
            I => \N__47807\
        );

    \I__11064\ : Span4Mux_v
    port map (
            O => \N__47823\,
            I => \N__47804\
        );

    \I__11063\ : InMux
    port map (
            O => \N__47822\,
            I => \N__47801\
        );

    \I__11062\ : Span4Mux_h
    port map (
            O => \N__47819\,
            I => \N__47796\
        );

    \I__11061\ : Span4Mux_v
    port map (
            O => \N__47814\,
            I => \N__47796\
        );

    \I__11060\ : LocalMux
    port map (
            O => \N__47807\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\
        );

    \I__11059\ : Odrv4
    port map (
            O => \N__47804\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\
        );

    \I__11058\ : LocalMux
    port map (
            O => \N__47801\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\
        );

    \I__11057\ : Odrv4
    port map (
            O => \N__47796\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\
        );

    \I__11056\ : CascadeMux
    port map (
            O => \N__47787\,
            I => \elapsed_time_ns_1_RNII6NQL1_0_1_cascade_\
        );

    \I__11055\ : InMux
    port map (
            O => \N__47784\,
            I => \N__47779\
        );

    \I__11054\ : InMux
    port map (
            O => \N__47783\,
            I => \N__47776\
        );

    \I__11053\ : InMux
    port map (
            O => \N__47782\,
            I => \N__47773\
        );

    \I__11052\ : LocalMux
    port map (
            O => \N__47779\,
            I => \N__47770\
        );

    \I__11051\ : LocalMux
    port map (
            O => \N__47776\,
            I => \N__47767\
        );

    \I__11050\ : LocalMux
    port map (
            O => \N__47773\,
            I => \N__47763\
        );

    \I__11049\ : Span4Mux_h
    port map (
            O => \N__47770\,
            I => \N__47760\
        );

    \I__11048\ : Sp12to4
    port map (
            O => \N__47767\,
            I => \N__47757\
        );

    \I__11047\ : InMux
    port map (
            O => \N__47766\,
            I => \N__47754\
        );

    \I__11046\ : Span4Mux_h
    port map (
            O => \N__47763\,
            I => \N__47751\
        );

    \I__11045\ : Odrv4
    port map (
            O => \N__47760\,
            I => \elapsed_time_ns_1_RNIBA65M1_0_19\
        );

    \I__11044\ : Odrv12
    port map (
            O => \N__47757\,
            I => \elapsed_time_ns_1_RNIBA65M1_0_19\
        );

    \I__11043\ : LocalMux
    port map (
            O => \N__47754\,
            I => \elapsed_time_ns_1_RNIBA65M1_0_19\
        );

    \I__11042\ : Odrv4
    port map (
            O => \N__47751\,
            I => \elapsed_time_ns_1_RNIBA65M1_0_19\
        );

    \I__11041\ : InMux
    port map (
            O => \N__47742\,
            I => \N__47739\
        );

    \I__11040\ : LocalMux
    port map (
            O => \N__47739\,
            I => \N__47736\
        );

    \I__11039\ : Span4Mux_v
    port map (
            O => \N__47736\,
            I => \N__47732\
        );

    \I__11038\ : InMux
    port map (
            O => \N__47735\,
            I => \N__47729\
        );

    \I__11037\ : Span4Mux_h
    port map (
            O => \N__47732\,
            I => \N__47723\
        );

    \I__11036\ : LocalMux
    port map (
            O => \N__47729\,
            I => \N__47723\
        );

    \I__11035\ : InMux
    port map (
            O => \N__47728\,
            I => \N__47720\
        );

    \I__11034\ : Odrv4
    port map (
            O => \N__47723\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__11033\ : LocalMux
    port map (
            O => \N__47720\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__11032\ : InMux
    port map (
            O => \N__47715\,
            I => \N__47712\
        );

    \I__11031\ : LocalMux
    port map (
            O => \N__47712\,
            I => \N__47709\
        );

    \I__11030\ : Span4Mux_h
    port map (
            O => \N__47709\,
            I => \N__47706\
        );

    \I__11029\ : Odrv4
    port map (
            O => \N__47706\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19\
        );

    \I__11028\ : InMux
    port map (
            O => \N__47703\,
            I => \N__47695\
        );

    \I__11027\ : InMux
    port map (
            O => \N__47702\,
            I => \N__47692\
        );

    \I__11026\ : CascadeMux
    port map (
            O => \N__47701\,
            I => \N__47687\
        );

    \I__11025\ : InMux
    port map (
            O => \N__47700\,
            I => \N__47684\
        );

    \I__11024\ : InMux
    port map (
            O => \N__47699\,
            I => \N__47681\
        );

    \I__11023\ : InMux
    port map (
            O => \N__47698\,
            I => \N__47678\
        );

    \I__11022\ : LocalMux
    port map (
            O => \N__47695\,
            I => \N__47672\
        );

    \I__11021\ : LocalMux
    port map (
            O => \N__47692\,
            I => \N__47672\
        );

    \I__11020\ : InMux
    port map (
            O => \N__47691\,
            I => \N__47669\
        );

    \I__11019\ : InMux
    port map (
            O => \N__47690\,
            I => \N__47663\
        );

    \I__11018\ : InMux
    port map (
            O => \N__47687\,
            I => \N__47663\
        );

    \I__11017\ : LocalMux
    port map (
            O => \N__47684\,
            I => \N__47659\
        );

    \I__11016\ : LocalMux
    port map (
            O => \N__47681\,
            I => \N__47656\
        );

    \I__11015\ : LocalMux
    port map (
            O => \N__47678\,
            I => \N__47653\
        );

    \I__11014\ : InMux
    port map (
            O => \N__47677\,
            I => \N__47650\
        );

    \I__11013\ : Span4Mux_v
    port map (
            O => \N__47672\,
            I => \N__47645\
        );

    \I__11012\ : LocalMux
    port map (
            O => \N__47669\,
            I => \N__47645\
        );

    \I__11011\ : InMux
    port map (
            O => \N__47668\,
            I => \N__47641\
        );

    \I__11010\ : LocalMux
    port map (
            O => \N__47663\,
            I => \N__47638\
        );

    \I__11009\ : InMux
    port map (
            O => \N__47662\,
            I => \N__47635\
        );

    \I__11008\ : Span4Mux_v
    port map (
            O => \N__47659\,
            I => \N__47627\
        );

    \I__11007\ : Span4Mux_v
    port map (
            O => \N__47656\,
            I => \N__47619\
        );

    \I__11006\ : Span4Mux_v
    port map (
            O => \N__47653\,
            I => \N__47619\
        );

    \I__11005\ : LocalMux
    port map (
            O => \N__47650\,
            I => \N__47619\
        );

    \I__11004\ : Span4Mux_h
    port map (
            O => \N__47645\,
            I => \N__47616\
        );

    \I__11003\ : CascadeMux
    port map (
            O => \N__47644\,
            I => \N__47612\
        );

    \I__11002\ : LocalMux
    port map (
            O => \N__47641\,
            I => \N__47605\
        );

    \I__11001\ : Span4Mux_h
    port map (
            O => \N__47638\,
            I => \N__47605\
        );

    \I__11000\ : LocalMux
    port map (
            O => \N__47635\,
            I => \N__47602\
        );

    \I__10999\ : InMux
    port map (
            O => \N__47634\,
            I => \N__47597\
        );

    \I__10998\ : InMux
    port map (
            O => \N__47633\,
            I => \N__47597\
        );

    \I__10997\ : InMux
    port map (
            O => \N__47632\,
            I => \N__47590\
        );

    \I__10996\ : InMux
    port map (
            O => \N__47631\,
            I => \N__47590\
        );

    \I__10995\ : InMux
    port map (
            O => \N__47630\,
            I => \N__47590\
        );

    \I__10994\ : Span4Mux_h
    port map (
            O => \N__47627\,
            I => \N__47587\
        );

    \I__10993\ : InMux
    port map (
            O => \N__47626\,
            I => \N__47584\
        );

    \I__10992\ : Span4Mux_h
    port map (
            O => \N__47619\,
            I => \N__47579\
        );

    \I__10991\ : Span4Mux_v
    port map (
            O => \N__47616\,
            I => \N__47579\
        );

    \I__10990\ : InMux
    port map (
            O => \N__47615\,
            I => \N__47576\
        );

    \I__10989\ : InMux
    port map (
            O => \N__47612\,
            I => \N__47569\
        );

    \I__10988\ : InMux
    port map (
            O => \N__47611\,
            I => \N__47569\
        );

    \I__10987\ : InMux
    port map (
            O => \N__47610\,
            I => \N__47569\
        );

    \I__10986\ : Span4Mux_h
    port map (
            O => \N__47605\,
            I => \N__47566\
        );

    \I__10985\ : Span12Mux_v
    port map (
            O => \N__47602\,
            I => \N__47559\
        );

    \I__10984\ : LocalMux
    port map (
            O => \N__47597\,
            I => \N__47559\
        );

    \I__10983\ : LocalMux
    port map (
            O => \N__47590\,
            I => \N__47559\
        );

    \I__10982\ : Odrv4
    port map (
            O => \N__47587\,
            I => \delay_measurement_inst.delay_tr9\
        );

    \I__10981\ : LocalMux
    port map (
            O => \N__47584\,
            I => \delay_measurement_inst.delay_tr9\
        );

    \I__10980\ : Odrv4
    port map (
            O => \N__47579\,
            I => \delay_measurement_inst.delay_tr9\
        );

    \I__10979\ : LocalMux
    port map (
            O => \N__47576\,
            I => \delay_measurement_inst.delay_tr9\
        );

    \I__10978\ : LocalMux
    port map (
            O => \N__47569\,
            I => \delay_measurement_inst.delay_tr9\
        );

    \I__10977\ : Odrv4
    port map (
            O => \N__47566\,
            I => \delay_measurement_inst.delay_tr9\
        );

    \I__10976\ : Odrv12
    port map (
            O => \N__47559\,
            I => \delay_measurement_inst.delay_tr9\
        );

    \I__10975\ : InMux
    port map (
            O => \N__47544\,
            I => \N__47541\
        );

    \I__10974\ : LocalMux
    port map (
            O => \N__47541\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1\
        );

    \I__10973\ : CascadeMux
    port map (
            O => \N__47538\,
            I => \N__47534\
        );

    \I__10972\ : InMux
    port map (
            O => \N__47537\,
            I => \N__47531\
        );

    \I__10971\ : InMux
    port map (
            O => \N__47534\,
            I => \N__47528\
        );

    \I__10970\ : LocalMux
    port map (
            O => \N__47531\,
            I => \N__47524\
        );

    \I__10969\ : LocalMux
    port map (
            O => \N__47528\,
            I => \N__47521\
        );

    \I__10968\ : InMux
    port map (
            O => \N__47527\,
            I => \N__47517\
        );

    \I__10967\ : Span4Mux_v
    port map (
            O => \N__47524\,
            I => \N__47512\
        );

    \I__10966\ : Span4Mux_v
    port map (
            O => \N__47521\,
            I => \N__47512\
        );

    \I__10965\ : InMux
    port map (
            O => \N__47520\,
            I => \N__47509\
        );

    \I__10964\ : LocalMux
    port map (
            O => \N__47517\,
            I => \elapsed_time_ns_1_RNIFJ2591_0_7\
        );

    \I__10963\ : Odrv4
    port map (
            O => \N__47512\,
            I => \elapsed_time_ns_1_RNIFJ2591_0_7\
        );

    \I__10962\ : LocalMux
    port map (
            O => \N__47509\,
            I => \elapsed_time_ns_1_RNIFJ2591_0_7\
        );

    \I__10961\ : InMux
    port map (
            O => \N__47502\,
            I => \N__47499\
        );

    \I__10960\ : LocalMux
    port map (
            O => \N__47499\,
            I => \N__47496\
        );

    \I__10959\ : Span12Mux_h
    port map (
            O => \N__47496\,
            I => \N__47493\
        );

    \I__10958\ : Odrv12
    port map (
            O => \N__47493\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\
        );

    \I__10957\ : InMux
    port map (
            O => \N__47490\,
            I => \N__47487\
        );

    \I__10956\ : LocalMux
    port map (
            O => \N__47487\,
            I => \N__47484\
        );

    \I__10955\ : Odrv12
    port map (
            O => \N__47484\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\
        );

    \I__10954\ : CascadeMux
    port map (
            O => \N__47481\,
            I => \N__47478\
        );

    \I__10953\ : InMux
    port map (
            O => \N__47478\,
            I => \N__47473\
        );

    \I__10952\ : InMux
    port map (
            O => \N__47477\,
            I => \N__47470\
        );

    \I__10951\ : InMux
    port map (
            O => \N__47476\,
            I => \N__47467\
        );

    \I__10950\ : LocalMux
    port map (
            O => \N__47473\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__10949\ : LocalMux
    port map (
            O => \N__47470\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__10948\ : LocalMux
    port map (
            O => \N__47467\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__10947\ : InMux
    port map (
            O => \N__47460\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__10946\ : CascadeMux
    port map (
            O => \N__47457\,
            I => \N__47454\
        );

    \I__10945\ : InMux
    port map (
            O => \N__47454\,
            I => \N__47449\
        );

    \I__10944\ : InMux
    port map (
            O => \N__47453\,
            I => \N__47446\
        );

    \I__10943\ : InMux
    port map (
            O => \N__47452\,
            I => \N__47443\
        );

    \I__10942\ : LocalMux
    port map (
            O => \N__47449\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__10941\ : LocalMux
    port map (
            O => \N__47446\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__10940\ : LocalMux
    port map (
            O => \N__47443\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__10939\ : InMux
    port map (
            O => \N__47436\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__10938\ : CascadeMux
    port map (
            O => \N__47433\,
            I => \N__47430\
        );

    \I__10937\ : InMux
    port map (
            O => \N__47430\,
            I => \N__47425\
        );

    \I__10936\ : InMux
    port map (
            O => \N__47429\,
            I => \N__47422\
        );

    \I__10935\ : InMux
    port map (
            O => \N__47428\,
            I => \N__47419\
        );

    \I__10934\ : LocalMux
    port map (
            O => \N__47425\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__10933\ : LocalMux
    port map (
            O => \N__47422\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__10932\ : LocalMux
    port map (
            O => \N__47419\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__10931\ : InMux
    port map (
            O => \N__47412\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__10930\ : CascadeMux
    port map (
            O => \N__47409\,
            I => \N__47406\
        );

    \I__10929\ : InMux
    port map (
            O => \N__47406\,
            I => \N__47401\
        );

    \I__10928\ : InMux
    port map (
            O => \N__47405\,
            I => \N__47398\
        );

    \I__10927\ : InMux
    port map (
            O => \N__47404\,
            I => \N__47395\
        );

    \I__10926\ : LocalMux
    port map (
            O => \N__47401\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__10925\ : LocalMux
    port map (
            O => \N__47398\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__10924\ : LocalMux
    port map (
            O => \N__47395\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__10923\ : InMux
    port map (
            O => \N__47388\,
            I => \bfn_18_21_0_\
        );

    \I__10922\ : CascadeMux
    port map (
            O => \N__47385\,
            I => \N__47382\
        );

    \I__10921\ : InMux
    port map (
            O => \N__47382\,
            I => \N__47377\
        );

    \I__10920\ : InMux
    port map (
            O => \N__47381\,
            I => \N__47374\
        );

    \I__10919\ : InMux
    port map (
            O => \N__47380\,
            I => \N__47371\
        );

    \I__10918\ : LocalMux
    port map (
            O => \N__47377\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__10917\ : LocalMux
    port map (
            O => \N__47374\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__10916\ : LocalMux
    port map (
            O => \N__47371\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__10915\ : InMux
    port map (
            O => \N__47364\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__10914\ : CascadeMux
    port map (
            O => \N__47361\,
            I => \N__47358\
        );

    \I__10913\ : InMux
    port map (
            O => \N__47358\,
            I => \N__47353\
        );

    \I__10912\ : InMux
    port map (
            O => \N__47357\,
            I => \N__47350\
        );

    \I__10911\ : InMux
    port map (
            O => \N__47356\,
            I => \N__47347\
        );

    \I__10910\ : LocalMux
    port map (
            O => \N__47353\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__10909\ : LocalMux
    port map (
            O => \N__47350\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__10908\ : LocalMux
    port map (
            O => \N__47347\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__10907\ : InMux
    port map (
            O => \N__47340\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__10906\ : CascadeMux
    port map (
            O => \N__47337\,
            I => \N__47334\
        );

    \I__10905\ : InMux
    port map (
            O => \N__47334\,
            I => \N__47329\
        );

    \I__10904\ : InMux
    port map (
            O => \N__47333\,
            I => \N__47326\
        );

    \I__10903\ : InMux
    port map (
            O => \N__47332\,
            I => \N__47323\
        );

    \I__10902\ : LocalMux
    port map (
            O => \N__47329\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__10901\ : LocalMux
    port map (
            O => \N__47326\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__10900\ : LocalMux
    port map (
            O => \N__47323\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__10899\ : InMux
    port map (
            O => \N__47316\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__10898\ : InMux
    port map (
            O => \N__47313\,
            I => \N__47309\
        );

    \I__10897\ : InMux
    port map (
            O => \N__47312\,
            I => \N__47306\
        );

    \I__10896\ : LocalMux
    port map (
            O => \N__47309\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__10895\ : LocalMux
    port map (
            O => \N__47306\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__10894\ : InMux
    port map (
            O => \N__47301\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__10893\ : CascadeMux
    port map (
            O => \N__47298\,
            I => \N__47295\
        );

    \I__10892\ : InMux
    port map (
            O => \N__47295\,
            I => \N__47290\
        );

    \I__10891\ : InMux
    port map (
            O => \N__47294\,
            I => \N__47287\
        );

    \I__10890\ : InMux
    port map (
            O => \N__47293\,
            I => \N__47284\
        );

    \I__10889\ : LocalMux
    port map (
            O => \N__47290\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__10888\ : LocalMux
    port map (
            O => \N__47287\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__10887\ : LocalMux
    port map (
            O => \N__47284\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__10886\ : InMux
    port map (
            O => \N__47277\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__10885\ : CascadeMux
    port map (
            O => \N__47274\,
            I => \N__47271\
        );

    \I__10884\ : InMux
    port map (
            O => \N__47271\,
            I => \N__47266\
        );

    \I__10883\ : InMux
    port map (
            O => \N__47270\,
            I => \N__47263\
        );

    \I__10882\ : InMux
    port map (
            O => \N__47269\,
            I => \N__47260\
        );

    \I__10881\ : LocalMux
    port map (
            O => \N__47266\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__10880\ : LocalMux
    port map (
            O => \N__47263\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__10879\ : LocalMux
    port map (
            O => \N__47260\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__10878\ : InMux
    port map (
            O => \N__47253\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__10877\ : CascadeMux
    port map (
            O => \N__47250\,
            I => \N__47247\
        );

    \I__10876\ : InMux
    port map (
            O => \N__47247\,
            I => \N__47242\
        );

    \I__10875\ : InMux
    port map (
            O => \N__47246\,
            I => \N__47239\
        );

    \I__10874\ : InMux
    port map (
            O => \N__47245\,
            I => \N__47236\
        );

    \I__10873\ : LocalMux
    port map (
            O => \N__47242\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__10872\ : LocalMux
    port map (
            O => \N__47239\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__10871\ : LocalMux
    port map (
            O => \N__47236\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__10870\ : InMux
    port map (
            O => \N__47229\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__10869\ : CascadeMux
    port map (
            O => \N__47226\,
            I => \N__47223\
        );

    \I__10868\ : InMux
    port map (
            O => \N__47223\,
            I => \N__47218\
        );

    \I__10867\ : InMux
    port map (
            O => \N__47222\,
            I => \N__47215\
        );

    \I__10866\ : InMux
    port map (
            O => \N__47221\,
            I => \N__47212\
        );

    \I__10865\ : LocalMux
    port map (
            O => \N__47218\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__10864\ : LocalMux
    port map (
            O => \N__47215\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__10863\ : LocalMux
    port map (
            O => \N__47212\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__10862\ : InMux
    port map (
            O => \N__47205\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__10861\ : CascadeMux
    port map (
            O => \N__47202\,
            I => \N__47199\
        );

    \I__10860\ : InMux
    port map (
            O => \N__47199\,
            I => \N__47194\
        );

    \I__10859\ : InMux
    port map (
            O => \N__47198\,
            I => \N__47191\
        );

    \I__10858\ : InMux
    port map (
            O => \N__47197\,
            I => \N__47188\
        );

    \I__10857\ : LocalMux
    port map (
            O => \N__47194\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__10856\ : LocalMux
    port map (
            O => \N__47191\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__10855\ : LocalMux
    port map (
            O => \N__47188\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__10854\ : InMux
    port map (
            O => \N__47181\,
            I => \bfn_18_20_0_\
        );

    \I__10853\ : CascadeMux
    port map (
            O => \N__47178\,
            I => \N__47175\
        );

    \I__10852\ : InMux
    port map (
            O => \N__47175\,
            I => \N__47170\
        );

    \I__10851\ : InMux
    port map (
            O => \N__47174\,
            I => \N__47167\
        );

    \I__10850\ : InMux
    port map (
            O => \N__47173\,
            I => \N__47164\
        );

    \I__10849\ : LocalMux
    port map (
            O => \N__47170\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__10848\ : LocalMux
    port map (
            O => \N__47167\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__10847\ : LocalMux
    port map (
            O => \N__47164\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__10846\ : InMux
    port map (
            O => \N__47157\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__10845\ : CascadeMux
    port map (
            O => \N__47154\,
            I => \N__47151\
        );

    \I__10844\ : InMux
    port map (
            O => \N__47151\,
            I => \N__47146\
        );

    \I__10843\ : InMux
    port map (
            O => \N__47150\,
            I => \N__47143\
        );

    \I__10842\ : InMux
    port map (
            O => \N__47149\,
            I => \N__47140\
        );

    \I__10841\ : LocalMux
    port map (
            O => \N__47146\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__10840\ : LocalMux
    port map (
            O => \N__47143\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__10839\ : LocalMux
    port map (
            O => \N__47140\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__10838\ : InMux
    port map (
            O => \N__47133\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__10837\ : CascadeMux
    port map (
            O => \N__47130\,
            I => \N__47127\
        );

    \I__10836\ : InMux
    port map (
            O => \N__47127\,
            I => \N__47122\
        );

    \I__10835\ : InMux
    port map (
            O => \N__47126\,
            I => \N__47119\
        );

    \I__10834\ : InMux
    port map (
            O => \N__47125\,
            I => \N__47116\
        );

    \I__10833\ : LocalMux
    port map (
            O => \N__47122\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__10832\ : LocalMux
    port map (
            O => \N__47119\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__10831\ : LocalMux
    port map (
            O => \N__47116\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__10830\ : InMux
    port map (
            O => \N__47109\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__10829\ : CascadeMux
    port map (
            O => \N__47106\,
            I => \N__47103\
        );

    \I__10828\ : InMux
    port map (
            O => \N__47103\,
            I => \N__47098\
        );

    \I__10827\ : InMux
    port map (
            O => \N__47102\,
            I => \N__47095\
        );

    \I__10826\ : InMux
    port map (
            O => \N__47101\,
            I => \N__47092\
        );

    \I__10825\ : LocalMux
    port map (
            O => \N__47098\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__10824\ : LocalMux
    port map (
            O => \N__47095\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__10823\ : LocalMux
    port map (
            O => \N__47092\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__10822\ : InMux
    port map (
            O => \N__47085\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__10821\ : CascadeMux
    port map (
            O => \N__47082\,
            I => \N__47079\
        );

    \I__10820\ : InMux
    port map (
            O => \N__47079\,
            I => \N__47074\
        );

    \I__10819\ : InMux
    port map (
            O => \N__47078\,
            I => \N__47071\
        );

    \I__10818\ : InMux
    port map (
            O => \N__47077\,
            I => \N__47068\
        );

    \I__10817\ : LocalMux
    port map (
            O => \N__47074\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__10816\ : LocalMux
    port map (
            O => \N__47071\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__10815\ : LocalMux
    port map (
            O => \N__47068\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__10814\ : InMux
    port map (
            O => \N__47061\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__10813\ : CascadeMux
    port map (
            O => \N__47058\,
            I => \N__47055\
        );

    \I__10812\ : InMux
    port map (
            O => \N__47055\,
            I => \N__47050\
        );

    \I__10811\ : InMux
    port map (
            O => \N__47054\,
            I => \N__47047\
        );

    \I__10810\ : InMux
    port map (
            O => \N__47053\,
            I => \N__47044\
        );

    \I__10809\ : LocalMux
    port map (
            O => \N__47050\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__10808\ : LocalMux
    port map (
            O => \N__47047\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__10807\ : LocalMux
    port map (
            O => \N__47044\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__10806\ : InMux
    port map (
            O => \N__47037\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__10805\ : CascadeMux
    port map (
            O => \N__47034\,
            I => \N__47031\
        );

    \I__10804\ : InMux
    port map (
            O => \N__47031\,
            I => \N__47026\
        );

    \I__10803\ : InMux
    port map (
            O => \N__47030\,
            I => \N__47023\
        );

    \I__10802\ : InMux
    port map (
            O => \N__47029\,
            I => \N__47020\
        );

    \I__10801\ : LocalMux
    port map (
            O => \N__47026\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__10800\ : LocalMux
    port map (
            O => \N__47023\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__10799\ : LocalMux
    port map (
            O => \N__47020\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__10798\ : InMux
    port map (
            O => \N__47013\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__10797\ : CascadeMux
    port map (
            O => \N__47010\,
            I => \N__47007\
        );

    \I__10796\ : InMux
    port map (
            O => \N__47007\,
            I => \N__47002\
        );

    \I__10795\ : InMux
    port map (
            O => \N__47006\,
            I => \N__46999\
        );

    \I__10794\ : InMux
    port map (
            O => \N__47005\,
            I => \N__46996\
        );

    \I__10793\ : LocalMux
    port map (
            O => \N__47002\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__10792\ : LocalMux
    port map (
            O => \N__46999\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__10791\ : LocalMux
    port map (
            O => \N__46996\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__10790\ : InMux
    port map (
            O => \N__46989\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__10789\ : CascadeMux
    port map (
            O => \N__46986\,
            I => \N__46983\
        );

    \I__10788\ : InMux
    port map (
            O => \N__46983\,
            I => \N__46978\
        );

    \I__10787\ : InMux
    port map (
            O => \N__46982\,
            I => \N__46975\
        );

    \I__10786\ : InMux
    port map (
            O => \N__46981\,
            I => \N__46972\
        );

    \I__10785\ : LocalMux
    port map (
            O => \N__46978\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__10784\ : LocalMux
    port map (
            O => \N__46975\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__10783\ : LocalMux
    port map (
            O => \N__46972\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__10782\ : InMux
    port map (
            O => \N__46965\,
            I => \bfn_18_19_0_\
        );

    \I__10781\ : CascadeMux
    port map (
            O => \N__46962\,
            I => \N__46959\
        );

    \I__10780\ : InMux
    port map (
            O => \N__46959\,
            I => \N__46954\
        );

    \I__10779\ : InMux
    port map (
            O => \N__46958\,
            I => \N__46951\
        );

    \I__10778\ : InMux
    port map (
            O => \N__46957\,
            I => \N__46948\
        );

    \I__10777\ : LocalMux
    port map (
            O => \N__46954\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__10776\ : LocalMux
    port map (
            O => \N__46951\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__10775\ : LocalMux
    port map (
            O => \N__46948\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__10774\ : InMux
    port map (
            O => \N__46941\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__10773\ : CascadeMux
    port map (
            O => \N__46938\,
            I => \N__46935\
        );

    \I__10772\ : InMux
    port map (
            O => \N__46935\,
            I => \N__46930\
        );

    \I__10771\ : InMux
    port map (
            O => \N__46934\,
            I => \N__46927\
        );

    \I__10770\ : InMux
    port map (
            O => \N__46933\,
            I => \N__46924\
        );

    \I__10769\ : LocalMux
    port map (
            O => \N__46930\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__10768\ : LocalMux
    port map (
            O => \N__46927\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__10767\ : LocalMux
    port map (
            O => \N__46924\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__10766\ : InMux
    port map (
            O => \N__46917\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__10765\ : CascadeMux
    port map (
            O => \N__46914\,
            I => \N__46911\
        );

    \I__10764\ : InMux
    port map (
            O => \N__46911\,
            I => \N__46906\
        );

    \I__10763\ : InMux
    port map (
            O => \N__46910\,
            I => \N__46903\
        );

    \I__10762\ : InMux
    port map (
            O => \N__46909\,
            I => \N__46900\
        );

    \I__10761\ : LocalMux
    port map (
            O => \N__46906\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__10760\ : LocalMux
    port map (
            O => \N__46903\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__46900\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__10758\ : InMux
    port map (
            O => \N__46893\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__10757\ : CascadeMux
    port map (
            O => \N__46890\,
            I => \N__46887\
        );

    \I__10756\ : InMux
    port map (
            O => \N__46887\,
            I => \N__46882\
        );

    \I__10755\ : InMux
    port map (
            O => \N__46886\,
            I => \N__46879\
        );

    \I__10754\ : InMux
    port map (
            O => \N__46885\,
            I => \N__46875\
        );

    \I__10753\ : LocalMux
    port map (
            O => \N__46882\,
            I => \N__46869\
        );

    \I__10752\ : LocalMux
    port map (
            O => \N__46879\,
            I => \N__46869\
        );

    \I__10751\ : InMux
    port map (
            O => \N__46878\,
            I => \N__46864\
        );

    \I__10750\ : LocalMux
    port map (
            O => \N__46875\,
            I => \N__46861\
        );

    \I__10749\ : InMux
    port map (
            O => \N__46874\,
            I => \N__46857\
        );

    \I__10748\ : Span4Mux_h
    port map (
            O => \N__46869\,
            I => \N__46854\
        );

    \I__10747\ : InMux
    port map (
            O => \N__46868\,
            I => \N__46851\
        );

    \I__10746\ : InMux
    port map (
            O => \N__46867\,
            I => \N__46848\
        );

    \I__10745\ : LocalMux
    port map (
            O => \N__46864\,
            I => \N__46843\
        );

    \I__10744\ : Span12Mux_v
    port map (
            O => \N__46861\,
            I => \N__46843\
        );

    \I__10743\ : InMux
    port map (
            O => \N__46860\,
            I => \N__46840\
        );

    \I__10742\ : LocalMux
    port map (
            O => \N__46857\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__10741\ : Odrv4
    port map (
            O => \N__46854\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__10740\ : LocalMux
    port map (
            O => \N__46851\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__10739\ : LocalMux
    port map (
            O => \N__46848\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__10738\ : Odrv12
    port map (
            O => \N__46843\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__10737\ : LocalMux
    port map (
            O => \N__46840\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__10736\ : CascadeMux
    port map (
            O => \N__46827\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2_cascade_\
        );

    \I__10735\ : InMux
    port map (
            O => \N__46824\,
            I => \N__46809\
        );

    \I__10734\ : InMux
    port map (
            O => \N__46823\,
            I => \N__46804\
        );

    \I__10733\ : InMux
    port map (
            O => \N__46822\,
            I => \N__46797\
        );

    \I__10732\ : InMux
    port map (
            O => \N__46821\,
            I => \N__46797\
        );

    \I__10731\ : InMux
    port map (
            O => \N__46820\,
            I => \N__46797\
        );

    \I__10730\ : InMux
    port map (
            O => \N__46819\,
            I => \N__46794\
        );

    \I__10729\ : InMux
    port map (
            O => \N__46818\,
            I => \N__46791\
        );

    \I__10728\ : InMux
    port map (
            O => \N__46817\,
            I => \N__46784\
        );

    \I__10727\ : InMux
    port map (
            O => \N__46816\,
            I => \N__46784\
        );

    \I__10726\ : InMux
    port map (
            O => \N__46815\,
            I => \N__46784\
        );

    \I__10725\ : InMux
    port map (
            O => \N__46814\,
            I => \N__46779\
        );

    \I__10724\ : InMux
    port map (
            O => \N__46813\,
            I => \N__46779\
        );

    \I__10723\ : InMux
    port map (
            O => \N__46812\,
            I => \N__46776\
        );

    \I__10722\ : LocalMux
    port map (
            O => \N__46809\,
            I => \N__46773\
        );

    \I__10721\ : CascadeMux
    port map (
            O => \N__46808\,
            I => \N__46769\
        );

    \I__10720\ : CascadeMux
    port map (
            O => \N__46807\,
            I => \N__46761\
        );

    \I__10719\ : LocalMux
    port map (
            O => \N__46804\,
            I => \N__46758\
        );

    \I__10718\ : LocalMux
    port map (
            O => \N__46797\,
            I => \N__46753\
        );

    \I__10717\ : LocalMux
    port map (
            O => \N__46794\,
            I => \N__46753\
        );

    \I__10716\ : LocalMux
    port map (
            O => \N__46791\,
            I => \N__46745\
        );

    \I__10715\ : LocalMux
    port map (
            O => \N__46784\,
            I => \N__46738\
        );

    \I__10714\ : LocalMux
    port map (
            O => \N__46779\,
            I => \N__46738\
        );

    \I__10713\ : LocalMux
    port map (
            O => \N__46776\,
            I => \N__46738\
        );

    \I__10712\ : Span4Mux_v
    port map (
            O => \N__46773\,
            I => \N__46735\
        );

    \I__10711\ : InMux
    port map (
            O => \N__46772\,
            I => \N__46728\
        );

    \I__10710\ : InMux
    port map (
            O => \N__46769\,
            I => \N__46728\
        );

    \I__10709\ : InMux
    port map (
            O => \N__46768\,
            I => \N__46728\
        );

    \I__10708\ : InMux
    port map (
            O => \N__46767\,
            I => \N__46722\
        );

    \I__10707\ : InMux
    port map (
            O => \N__46766\,
            I => \N__46722\
        );

    \I__10706\ : InMux
    port map (
            O => \N__46765\,
            I => \N__46715\
        );

    \I__10705\ : InMux
    port map (
            O => \N__46764\,
            I => \N__46715\
        );

    \I__10704\ : InMux
    port map (
            O => \N__46761\,
            I => \N__46715\
        );

    \I__10703\ : Span4Mux_h
    port map (
            O => \N__46758\,
            I => \N__46712\
        );

    \I__10702\ : Span4Mux_v
    port map (
            O => \N__46753\,
            I => \N__46709\
        );

    \I__10701\ : InMux
    port map (
            O => \N__46752\,
            I => \N__46698\
        );

    \I__10700\ : InMux
    port map (
            O => \N__46751\,
            I => \N__46698\
        );

    \I__10699\ : InMux
    port map (
            O => \N__46750\,
            I => \N__46698\
        );

    \I__10698\ : InMux
    port map (
            O => \N__46749\,
            I => \N__46698\
        );

    \I__10697\ : InMux
    port map (
            O => \N__46748\,
            I => \N__46698\
        );

    \I__10696\ : Span4Mux_v
    port map (
            O => \N__46745\,
            I => \N__46689\
        );

    \I__10695\ : Span4Mux_v
    port map (
            O => \N__46738\,
            I => \N__46689\
        );

    \I__10694\ : Span4Mux_v
    port map (
            O => \N__46735\,
            I => \N__46689\
        );

    \I__10693\ : LocalMux
    port map (
            O => \N__46728\,
            I => \N__46689\
        );

    \I__10692\ : InMux
    port map (
            O => \N__46727\,
            I => \N__46686\
        );

    \I__10691\ : LocalMux
    port map (
            O => \N__46722\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__10690\ : LocalMux
    port map (
            O => \N__46715\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__10689\ : Odrv4
    port map (
            O => \N__46712\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__10688\ : Odrv4
    port map (
            O => \N__46709\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__10687\ : LocalMux
    port map (
            O => \N__46698\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__10686\ : Odrv4
    port map (
            O => \N__46689\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__10685\ : LocalMux
    port map (
            O => \N__46686\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__10684\ : CascadeMux
    port map (
            O => \N__46671\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6_cascade_\
        );

    \I__10683\ : CascadeMux
    port map (
            O => \N__46668\,
            I => \N__46665\
        );

    \I__10682\ : InMux
    port map (
            O => \N__46665\,
            I => \N__46662\
        );

    \I__10681\ : LocalMux
    port map (
            O => \N__46662\,
            I => \N__46659\
        );

    \I__10680\ : Odrv12
    port map (
            O => \N__46659\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\
        );

    \I__10679\ : InMux
    port map (
            O => \N__46656\,
            I => \N__46653\
        );

    \I__10678\ : LocalMux
    port map (
            O => \N__46653\,
            I => \N__46650\
        );

    \I__10677\ : Span4Mux_v
    port map (
            O => \N__46650\,
            I => \N__46647\
        );

    \I__10676\ : Odrv4
    port map (
            O => \N__46647\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\
        );

    \I__10675\ : InMux
    port map (
            O => \N__46644\,
            I => \N__46641\
        );

    \I__10674\ : LocalMux
    port map (
            O => \N__46641\,
            I => \N__46638\
        );

    \I__10673\ : Span4Mux_h
    port map (
            O => \N__46638\,
            I => \N__46635\
        );

    \I__10672\ : Odrv4
    port map (
            O => \N__46635\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\
        );

    \I__10671\ : InMux
    port map (
            O => \N__46632\,
            I => \N__46627\
        );

    \I__10670\ : InMux
    port map (
            O => \N__46631\,
            I => \N__46622\
        );

    \I__10669\ : InMux
    port map (
            O => \N__46630\,
            I => \N__46622\
        );

    \I__10668\ : LocalMux
    port map (
            O => \N__46627\,
            I => \elapsed_time_ns_1_RNINBNQL1_0_6\
        );

    \I__10667\ : LocalMux
    port map (
            O => \N__46622\,
            I => \elapsed_time_ns_1_RNINBNQL1_0_6\
        );

    \I__10666\ : InMux
    port map (
            O => \N__46617\,
            I => \N__46614\
        );

    \I__10665\ : LocalMux
    port map (
            O => \N__46614\,
            I => \N__46611\
        );

    \I__10664\ : Span4Mux_h
    port map (
            O => \N__46611\,
            I => \N__46608\
        );

    \I__10663\ : Odrv4
    port map (
            O => \N__46608\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\
        );

    \I__10662\ : InMux
    port map (
            O => \N__46605\,
            I => \bfn_18_18_0_\
        );

    \I__10661\ : InMux
    port map (
            O => \N__46602\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__10660\ : CascadeMux
    port map (
            O => \N__46599\,
            I => \N__46596\
        );

    \I__10659\ : InMux
    port map (
            O => \N__46596\,
            I => \N__46591\
        );

    \I__10658\ : InMux
    port map (
            O => \N__46595\,
            I => \N__46588\
        );

    \I__10657\ : InMux
    port map (
            O => \N__46594\,
            I => \N__46585\
        );

    \I__10656\ : LocalMux
    port map (
            O => \N__46591\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__10655\ : LocalMux
    port map (
            O => \N__46588\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__10654\ : LocalMux
    port map (
            O => \N__46585\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__10653\ : InMux
    port map (
            O => \N__46578\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__10652\ : CascadeMux
    port map (
            O => \N__46575\,
            I => \N__46572\
        );

    \I__10651\ : InMux
    port map (
            O => \N__46572\,
            I => \N__46567\
        );

    \I__10650\ : InMux
    port map (
            O => \N__46571\,
            I => \N__46564\
        );

    \I__10649\ : InMux
    port map (
            O => \N__46570\,
            I => \N__46561\
        );

    \I__10648\ : LocalMux
    port map (
            O => \N__46567\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__10647\ : LocalMux
    port map (
            O => \N__46564\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__10646\ : LocalMux
    port map (
            O => \N__46561\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__10645\ : InMux
    port map (
            O => \N__46554\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__10644\ : CascadeMux
    port map (
            O => \N__46551\,
            I => \N__46548\
        );

    \I__10643\ : InMux
    port map (
            O => \N__46548\,
            I => \N__46544\
        );

    \I__10642\ : InMux
    port map (
            O => \N__46547\,
            I => \N__46541\
        );

    \I__10641\ : LocalMux
    port map (
            O => \N__46544\,
            I => \N__46538\
        );

    \I__10640\ : LocalMux
    port map (
            O => \N__46541\,
            I => \N__46533\
        );

    \I__10639\ : Span4Mux_v
    port map (
            O => \N__46538\,
            I => \N__46530\
        );

    \I__10638\ : InMux
    port map (
            O => \N__46537\,
            I => \N__46525\
        );

    \I__10637\ : InMux
    port map (
            O => \N__46536\,
            I => \N__46525\
        );

    \I__10636\ : Odrv4
    port map (
            O => \N__46533\,
            I => \elapsed_time_ns_1_RNIDH2591_0_5\
        );

    \I__10635\ : Odrv4
    port map (
            O => \N__46530\,
            I => \elapsed_time_ns_1_RNIDH2591_0_5\
        );

    \I__10634\ : LocalMux
    port map (
            O => \N__46525\,
            I => \elapsed_time_ns_1_RNIDH2591_0_5\
        );

    \I__10633\ : InMux
    port map (
            O => \N__46518\,
            I => \N__46515\
        );

    \I__10632\ : LocalMux
    port map (
            O => \N__46515\,
            I => \N__46512\
        );

    \I__10631\ : Span4Mux_v
    port map (
            O => \N__46512\,
            I => \N__46509\
        );

    \I__10630\ : Span4Mux_h
    port map (
            O => \N__46509\,
            I => \N__46506\
        );

    \I__10629\ : Odrv4
    port map (
            O => \N__46506\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\
        );

    \I__10628\ : InMux
    port map (
            O => \N__46503\,
            I => \N__46500\
        );

    \I__10627\ : LocalMux
    port map (
            O => \N__46500\,
            I => \N__46497\
        );

    \I__10626\ : Span4Mux_v
    port map (
            O => \N__46497\,
            I => \N__46494\
        );

    \I__10625\ : Span4Mux_h
    port map (
            O => \N__46494\,
            I => \N__46491\
        );

    \I__10624\ : Span4Mux_h
    port map (
            O => \N__46491\,
            I => \N__46488\
        );

    \I__10623\ : Odrv4
    port map (
            O => \N__46488\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\
        );

    \I__10622\ : InMux
    port map (
            O => \N__46485\,
            I => \N__46481\
        );

    \I__10621\ : InMux
    port map (
            O => \N__46484\,
            I => \N__46477\
        );

    \I__10620\ : LocalMux
    port map (
            O => \N__46481\,
            I => \N__46474\
        );

    \I__10619\ : InMux
    port map (
            O => \N__46480\,
            I => \N__46469\
        );

    \I__10618\ : LocalMux
    port map (
            O => \N__46477\,
            I => \N__46466\
        );

    \I__10617\ : Span4Mux_v
    port map (
            O => \N__46474\,
            I => \N__46463\
        );

    \I__10616\ : InMux
    port map (
            O => \N__46473\,
            I => \N__46460\
        );

    \I__10615\ : InMux
    port map (
            O => \N__46472\,
            I => \N__46457\
        );

    \I__10614\ : LocalMux
    port map (
            O => \N__46469\,
            I => \elapsed_time_ns_1_RNI8765M1_0_16\
        );

    \I__10613\ : Odrv12
    port map (
            O => \N__46466\,
            I => \elapsed_time_ns_1_RNI8765M1_0_16\
        );

    \I__10612\ : Odrv4
    port map (
            O => \N__46463\,
            I => \elapsed_time_ns_1_RNI8765M1_0_16\
        );

    \I__10611\ : LocalMux
    port map (
            O => \N__46460\,
            I => \elapsed_time_ns_1_RNI8765M1_0_16\
        );

    \I__10610\ : LocalMux
    port map (
            O => \N__46457\,
            I => \elapsed_time_ns_1_RNI8765M1_0_16\
        );

    \I__10609\ : CascadeMux
    port map (
            O => \N__46446\,
            I => \N__46442\
        );

    \I__10608\ : InMux
    port map (
            O => \N__46445\,
            I => \N__46437\
        );

    \I__10607\ : InMux
    port map (
            O => \N__46442\,
            I => \N__46437\
        );

    \I__10606\ : LocalMux
    port map (
            O => \N__46437\,
            I => \N__46434\
        );

    \I__10605\ : Span4Mux_h
    port map (
            O => \N__46434\,
            I => \N__46431\
        );

    \I__10604\ : Odrv4
    port map (
            O => \N__46431\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\
        );

    \I__10603\ : InMux
    port map (
            O => \N__46428\,
            I => \N__46424\
        );

    \I__10602\ : InMux
    port map (
            O => \N__46427\,
            I => \N__46419\
        );

    \I__10601\ : LocalMux
    port map (
            O => \N__46424\,
            I => \N__46416\
        );

    \I__10600\ : InMux
    port map (
            O => \N__46423\,
            I => \N__46413\
        );

    \I__10599\ : InMux
    port map (
            O => \N__46422\,
            I => \N__46410\
        );

    \I__10598\ : LocalMux
    port map (
            O => \N__46419\,
            I => \elapsed_time_ns_1_RNIK8NQL1_0_3\
        );

    \I__10597\ : Odrv4
    port map (
            O => \N__46416\,
            I => \elapsed_time_ns_1_RNIK8NQL1_0_3\
        );

    \I__10596\ : LocalMux
    port map (
            O => \N__46413\,
            I => \elapsed_time_ns_1_RNIK8NQL1_0_3\
        );

    \I__10595\ : LocalMux
    port map (
            O => \N__46410\,
            I => \elapsed_time_ns_1_RNIK8NQL1_0_3\
        );

    \I__10594\ : InMux
    port map (
            O => \N__46401\,
            I => \N__46396\
        );

    \I__10593\ : InMux
    port map (
            O => \N__46400\,
            I => \N__46391\
        );

    \I__10592\ : InMux
    port map (
            O => \N__46399\,
            I => \N__46391\
        );

    \I__10591\ : LocalMux
    port map (
            O => \N__46396\,
            I => \elapsed_time_ns_1_RNIAE2591_0_2\
        );

    \I__10590\ : LocalMux
    port map (
            O => \N__46391\,
            I => \elapsed_time_ns_1_RNIAE2591_0_2\
        );

    \I__10589\ : CascadeMux
    port map (
            O => \N__46386\,
            I => \N__46383\
        );

    \I__10588\ : InMux
    port map (
            O => \N__46383\,
            I => \N__46379\
        );

    \I__10587\ : InMux
    port map (
            O => \N__46382\,
            I => \N__46376\
        );

    \I__10586\ : LocalMux
    port map (
            O => \N__46379\,
            I => \N__46373\
        );

    \I__10585\ : LocalMux
    port map (
            O => \N__46376\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3\
        );

    \I__10584\ : Odrv4
    port map (
            O => \N__46373\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3\
        );

    \I__10583\ : InMux
    port map (
            O => \N__46368\,
            I => \N__46359\
        );

    \I__10582\ : InMux
    port map (
            O => \N__46367\,
            I => \N__46359\
        );

    \I__10581\ : InMux
    port map (
            O => \N__46366\,
            I => \N__46359\
        );

    \I__10580\ : LocalMux
    port map (
            O => \N__46359\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_0_2\
        );

    \I__10579\ : InMux
    port map (
            O => \N__46356\,
            I => \N__46353\
        );

    \I__10578\ : LocalMux
    port map (
            O => \N__46353\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2Z0Z_1\
        );

    \I__10577\ : InMux
    port map (
            O => \N__46350\,
            I => \N__46347\
        );

    \I__10576\ : LocalMux
    port map (
            O => \N__46347\,
            I => \N__46341\
        );

    \I__10575\ : InMux
    port map (
            O => \N__46346\,
            I => \N__46338\
        );

    \I__10574\ : InMux
    port map (
            O => \N__46345\,
            I => \N__46333\
        );

    \I__10573\ : InMux
    port map (
            O => \N__46344\,
            I => \N__46333\
        );

    \I__10572\ : Odrv4
    port map (
            O => \N__46341\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\
        );

    \I__10571\ : LocalMux
    port map (
            O => \N__46338\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\
        );

    \I__10570\ : LocalMux
    port map (
            O => \N__46333\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\
        );

    \I__10569\ : CascadeMux
    port map (
            O => \N__46326\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6_cascade_\
        );

    \I__10568\ : CascadeMux
    port map (
            O => \N__46323\,
            I => \elapsed_time_ns_1_RNINBNQL1_0_6_cascade_\
        );

    \I__10567\ : InMux
    port map (
            O => \N__46320\,
            I => \N__46317\
        );

    \I__10566\ : LocalMux
    port map (
            O => \N__46317\,
            I => \N__46314\
        );

    \I__10565\ : Span4Mux_v
    port map (
            O => \N__46314\,
            I => \N__46311\
        );

    \I__10564\ : Span4Mux_h
    port map (
            O => \N__46311\,
            I => \N__46307\
        );

    \I__10563\ : InMux
    port map (
            O => \N__46310\,
            I => \N__46304\
        );

    \I__10562\ : Odrv4
    port map (
            O => \N__46307\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2\
        );

    \I__10561\ : LocalMux
    port map (
            O => \N__46304\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2\
        );

    \I__10560\ : CascadeMux
    port map (
            O => \N__46299\,
            I => \N__46295\
        );

    \I__10559\ : CascadeMux
    port map (
            O => \N__46298\,
            I => \N__46291\
        );

    \I__10558\ : InMux
    port map (
            O => \N__46295\,
            I => \N__46284\
        );

    \I__10557\ : InMux
    port map (
            O => \N__46294\,
            I => \N__46284\
        );

    \I__10556\ : InMux
    port map (
            O => \N__46291\,
            I => \N__46284\
        );

    \I__10555\ : LocalMux
    port map (
            O => \N__46284\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2\
        );

    \I__10554\ : CascadeMux
    port map (
            O => \N__46281\,
            I => \N__46278\
        );

    \I__10553\ : InMux
    port map (
            O => \N__46278\,
            I => \N__46274\
        );

    \I__10552\ : CascadeMux
    port map (
            O => \N__46277\,
            I => \N__46270\
        );

    \I__10551\ : LocalMux
    port map (
            O => \N__46274\,
            I => \N__46266\
        );

    \I__10550\ : CascadeMux
    port map (
            O => \N__46273\,
            I => \N__46263\
        );

    \I__10549\ : InMux
    port map (
            O => \N__46270\,
            I => \N__46258\
        );

    \I__10548\ : InMux
    port map (
            O => \N__46269\,
            I => \N__46258\
        );

    \I__10547\ : Span4Mux_v
    port map (
            O => \N__46266\,
            I => \N__46255\
        );

    \I__10546\ : InMux
    port map (
            O => \N__46263\,
            I => \N__46252\
        );

    \I__10545\ : LocalMux
    port map (
            O => \N__46258\,
            I => \N__46249\
        );

    \I__10544\ : Span4Mux_h
    port map (
            O => \N__46255\,
            I => \N__46246\
        );

    \I__10543\ : LocalMux
    port map (
            O => \N__46252\,
            I => \N__46241\
        );

    \I__10542\ : Span4Mux_v
    port map (
            O => \N__46249\,
            I => \N__46241\
        );

    \I__10541\ : Odrv4
    port map (
            O => \N__46246\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__10540\ : Odrv4
    port map (
            O => \N__46241\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__10539\ : InMux
    port map (
            O => \N__46236\,
            I => \N__46233\
        );

    \I__10538\ : LocalMux
    port map (
            O => \N__46233\,
            I => \N__46228\
        );

    \I__10537\ : InMux
    port map (
            O => \N__46232\,
            I => \N__46225\
        );

    \I__10536\ : InMux
    port map (
            O => \N__46231\,
            I => \N__46222\
        );

    \I__10535\ : Odrv4
    port map (
            O => \N__46228\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__10534\ : LocalMux
    port map (
            O => \N__46225\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__10533\ : LocalMux
    port map (
            O => \N__46222\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__10532\ : CascadeMux
    port map (
            O => \N__46215\,
            I => \N__46212\
        );

    \I__10531\ : InMux
    port map (
            O => \N__46212\,
            I => \N__46209\
        );

    \I__10530\ : LocalMux
    port map (
            O => \N__46209\,
            I => \N__46206\
        );

    \I__10529\ : Span4Mux_v
    port map (
            O => \N__46206\,
            I => \N__46203\
        );

    \I__10528\ : Odrv4
    port map (
            O => \N__46203\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\
        );

    \I__10527\ : InMux
    port map (
            O => \N__46200\,
            I => \N__46197\
        );

    \I__10526\ : LocalMux
    port map (
            O => \N__46197\,
            I => \current_shift_inst.un4_control_input_1_axb_20\
        );

    \I__10525\ : CascadeMux
    port map (
            O => \N__46194\,
            I => \N__46190\
        );

    \I__10524\ : InMux
    port map (
            O => \N__46193\,
            I => \N__46186\
        );

    \I__10523\ : InMux
    port map (
            O => \N__46190\,
            I => \N__46183\
        );

    \I__10522\ : InMux
    port map (
            O => \N__46189\,
            I => \N__46180\
        );

    \I__10521\ : LocalMux
    port map (
            O => \N__46186\,
            I => \N__46177\
        );

    \I__10520\ : LocalMux
    port map (
            O => \N__46183\,
            I => \N__46174\
        );

    \I__10519\ : LocalMux
    port map (
            O => \N__46180\,
            I => \N__46171\
        );

    \I__10518\ : Span4Mux_v
    port map (
            O => \N__46177\,
            I => \N__46166\
        );

    \I__10517\ : Span4Mux_h
    port map (
            O => \N__46174\,
            I => \N__46166\
        );

    \I__10516\ : Span4Mux_v
    port map (
            O => \N__46171\,
            I => \N__46163\
        );

    \I__10515\ : Span4Mux_h
    port map (
            O => \N__46166\,
            I => \N__46159\
        );

    \I__10514\ : Span4Mux_h
    port map (
            O => \N__46163\,
            I => \N__46156\
        );

    \I__10513\ : InMux
    port map (
            O => \N__46162\,
            I => \N__46153\
        );

    \I__10512\ : Odrv4
    port map (
            O => \N__46159\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__10511\ : Odrv4
    port map (
            O => \N__46156\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__10510\ : LocalMux
    port map (
            O => \N__46153\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__10509\ : InMux
    port map (
            O => \N__46146\,
            I => \N__46143\
        );

    \I__10508\ : LocalMux
    port map (
            O => \N__46143\,
            I => \N__46140\
        );

    \I__10507\ : Span4Mux_v
    port map (
            O => \N__46140\,
            I => \N__46135\
        );

    \I__10506\ : InMux
    port map (
            O => \N__46139\,
            I => \N__46132\
        );

    \I__10505\ : InMux
    port map (
            O => \N__46138\,
            I => \N__46129\
        );

    \I__10504\ : Odrv4
    port map (
            O => \N__46135\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__10503\ : LocalMux
    port map (
            O => \N__46132\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__10502\ : LocalMux
    port map (
            O => \N__46129\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__10501\ : InMux
    port map (
            O => \N__46122\,
            I => \N__46119\
        );

    \I__10500\ : LocalMux
    port map (
            O => \N__46119\,
            I => \N__46116\
        );

    \I__10499\ : Odrv4
    port map (
            O => \N__46116\,
            I => \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\
        );

    \I__10498\ : CascadeMux
    port map (
            O => \N__46113\,
            I => \N__46109\
        );

    \I__10497\ : CascadeMux
    port map (
            O => \N__46112\,
            I => \N__46106\
        );

    \I__10496\ : InMux
    port map (
            O => \N__46109\,
            I => \N__46102\
        );

    \I__10495\ : InMux
    port map (
            O => \N__46106\,
            I => \N__46099\
        );

    \I__10494\ : InMux
    port map (
            O => \N__46105\,
            I => \N__46096\
        );

    \I__10493\ : LocalMux
    port map (
            O => \N__46102\,
            I => \N__46092\
        );

    \I__10492\ : LocalMux
    port map (
            O => \N__46099\,
            I => \N__46089\
        );

    \I__10491\ : LocalMux
    port map (
            O => \N__46096\,
            I => \N__46086\
        );

    \I__10490\ : InMux
    port map (
            O => \N__46095\,
            I => \N__46083\
        );

    \I__10489\ : Span4Mux_h
    port map (
            O => \N__46092\,
            I => \N__46080\
        );

    \I__10488\ : Span4Mux_v
    port map (
            O => \N__46089\,
            I => \N__46077\
        );

    \I__10487\ : Span4Mux_h
    port map (
            O => \N__46086\,
            I => \N__46074\
        );

    \I__10486\ : LocalMux
    port map (
            O => \N__46083\,
            I => \N__46071\
        );

    \I__10485\ : Span4Mux_h
    port map (
            O => \N__46080\,
            I => \N__46068\
        );

    \I__10484\ : Span4Mux_h
    port map (
            O => \N__46077\,
            I => \N__46063\
        );

    \I__10483\ : Span4Mux_h
    port map (
            O => \N__46074\,
            I => \N__46063\
        );

    \I__10482\ : Odrv12
    port map (
            O => \N__46071\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__10481\ : Odrv4
    port map (
            O => \N__46068\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__10480\ : Odrv4
    port map (
            O => \N__46063\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__10479\ : InMux
    port map (
            O => \N__46056\,
            I => \N__46053\
        );

    \I__10478\ : LocalMux
    port map (
            O => \N__46053\,
            I => \N__46049\
        );

    \I__10477\ : InMux
    port map (
            O => \N__46052\,
            I => \N__46046\
        );

    \I__10476\ : Span4Mux_v
    port map (
            O => \N__46049\,
            I => \N__46042\
        );

    \I__10475\ : LocalMux
    port map (
            O => \N__46046\,
            I => \N__46039\
        );

    \I__10474\ : InMux
    port map (
            O => \N__46045\,
            I => \N__46036\
        );

    \I__10473\ : Odrv4
    port map (
            O => \N__46042\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__10472\ : Odrv4
    port map (
            O => \N__46039\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__10471\ : LocalMux
    port map (
            O => \N__46036\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__10470\ : CascadeMux
    port map (
            O => \N__46029\,
            I => \N__46026\
        );

    \I__10469\ : InMux
    port map (
            O => \N__46026\,
            I => \N__46023\
        );

    \I__10468\ : LocalMux
    port map (
            O => \N__46023\,
            I => \N__46020\
        );

    \I__10467\ : Span4Mux_h
    port map (
            O => \N__46020\,
            I => \N__46017\
        );

    \I__10466\ : Odrv4
    port map (
            O => \N__46017\,
            I => \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\
        );

    \I__10465\ : CascadeMux
    port map (
            O => \N__46014\,
            I => \N__45989\
        );

    \I__10464\ : CascadeMux
    port map (
            O => \N__46013\,
            I => \N__45983\
        );

    \I__10463\ : CascadeMux
    port map (
            O => \N__46012\,
            I => \N__45977\
        );

    \I__10462\ : InMux
    port map (
            O => \N__46011\,
            I => \N__45965\
        );

    \I__10461\ : InMux
    port map (
            O => \N__46010\,
            I => \N__45965\
        );

    \I__10460\ : InMux
    port map (
            O => \N__46009\,
            I => \N__45965\
        );

    \I__10459\ : InMux
    port map (
            O => \N__46008\,
            I => \N__45965\
        );

    \I__10458\ : InMux
    port map (
            O => \N__46007\,
            I => \N__45956\
        );

    \I__10457\ : InMux
    port map (
            O => \N__46006\,
            I => \N__45956\
        );

    \I__10456\ : InMux
    port map (
            O => \N__46005\,
            I => \N__45956\
        );

    \I__10455\ : InMux
    port map (
            O => \N__46004\,
            I => \N__45956\
        );

    \I__10454\ : CascadeMux
    port map (
            O => \N__46003\,
            I => \N__45949\
        );

    \I__10453\ : CascadeMux
    port map (
            O => \N__46002\,
            I => \N__45936\
        );

    \I__10452\ : CascadeMux
    port map (
            O => \N__46001\,
            I => \N__45932\
        );

    \I__10451\ : CascadeMux
    port map (
            O => \N__46000\,
            I => \N__45928\
        );

    \I__10450\ : CascadeMux
    port map (
            O => \N__45999\,
            I => \N__45924\
        );

    \I__10449\ : CascadeMux
    port map (
            O => \N__45998\,
            I => \N__45920\
        );

    \I__10448\ : CascadeMux
    port map (
            O => \N__45997\,
            I => \N__45916\
        );

    \I__10447\ : CascadeMux
    port map (
            O => \N__45996\,
            I => \N__45912\
        );

    \I__10446\ : CascadeMux
    port map (
            O => \N__45995\,
            I => \N__45897\
        );

    \I__10445\ : CascadeMux
    port map (
            O => \N__45994\,
            I => \N__45893\
        );

    \I__10444\ : CascadeMux
    port map (
            O => \N__45993\,
            I => \N__45889\
        );

    \I__10443\ : InMux
    port map (
            O => \N__45992\,
            I => \N__45877\
        );

    \I__10442\ : InMux
    port map (
            O => \N__45989\,
            I => \N__45877\
        );

    \I__10441\ : InMux
    port map (
            O => \N__45988\,
            I => \N__45871\
        );

    \I__10440\ : InMux
    port map (
            O => \N__45987\,
            I => \N__45864\
        );

    \I__10439\ : InMux
    port map (
            O => \N__45986\,
            I => \N__45864\
        );

    \I__10438\ : InMux
    port map (
            O => \N__45983\,
            I => \N__45864\
        );

    \I__10437\ : InMux
    port map (
            O => \N__45982\,
            I => \N__45853\
        );

    \I__10436\ : InMux
    port map (
            O => \N__45981\,
            I => \N__45853\
        );

    \I__10435\ : InMux
    port map (
            O => \N__45980\,
            I => \N__45853\
        );

    \I__10434\ : InMux
    port map (
            O => \N__45977\,
            I => \N__45853\
        );

    \I__10433\ : InMux
    port map (
            O => \N__45976\,
            I => \N__45853\
        );

    \I__10432\ : CascadeMux
    port map (
            O => \N__45975\,
            I => \N__45849\
        );

    \I__10431\ : CascadeMux
    port map (
            O => \N__45974\,
            I => \N__45845\
        );

    \I__10430\ : LocalMux
    port map (
            O => \N__45965\,
            I => \N__45835\
        );

    \I__10429\ : LocalMux
    port map (
            O => \N__45956\,
            I => \N__45835\
        );

    \I__10428\ : InMux
    port map (
            O => \N__45955\,
            I => \N__45822\
        );

    \I__10427\ : InMux
    port map (
            O => \N__45954\,
            I => \N__45822\
        );

    \I__10426\ : InMux
    port map (
            O => \N__45953\,
            I => \N__45822\
        );

    \I__10425\ : InMux
    port map (
            O => \N__45952\,
            I => \N__45822\
        );

    \I__10424\ : InMux
    port map (
            O => \N__45949\,
            I => \N__45822\
        );

    \I__10423\ : InMux
    port map (
            O => \N__45948\,
            I => \N__45822\
        );

    \I__10422\ : InMux
    port map (
            O => \N__45947\,
            I => \N__45811\
        );

    \I__10421\ : InMux
    port map (
            O => \N__45946\,
            I => \N__45811\
        );

    \I__10420\ : InMux
    port map (
            O => \N__45945\,
            I => \N__45811\
        );

    \I__10419\ : InMux
    port map (
            O => \N__45944\,
            I => \N__45811\
        );

    \I__10418\ : InMux
    port map (
            O => \N__45943\,
            I => \N__45811\
        );

    \I__10417\ : InMux
    port map (
            O => \N__45942\,
            I => \N__45806\
        );

    \I__10416\ : InMux
    port map (
            O => \N__45941\,
            I => \N__45806\
        );

    \I__10415\ : InMux
    port map (
            O => \N__45940\,
            I => \N__45784\
        );

    \I__10414\ : InMux
    port map (
            O => \N__45939\,
            I => \N__45784\
        );

    \I__10413\ : InMux
    port map (
            O => \N__45936\,
            I => \N__45784\
        );

    \I__10412\ : InMux
    port map (
            O => \N__45935\,
            I => \N__45784\
        );

    \I__10411\ : InMux
    port map (
            O => \N__45932\,
            I => \N__45784\
        );

    \I__10410\ : InMux
    port map (
            O => \N__45931\,
            I => \N__45784\
        );

    \I__10409\ : InMux
    port map (
            O => \N__45928\,
            I => \N__45784\
        );

    \I__10408\ : InMux
    port map (
            O => \N__45927\,
            I => \N__45784\
        );

    \I__10407\ : InMux
    port map (
            O => \N__45924\,
            I => \N__45767\
        );

    \I__10406\ : InMux
    port map (
            O => \N__45923\,
            I => \N__45767\
        );

    \I__10405\ : InMux
    port map (
            O => \N__45920\,
            I => \N__45767\
        );

    \I__10404\ : InMux
    port map (
            O => \N__45919\,
            I => \N__45767\
        );

    \I__10403\ : InMux
    port map (
            O => \N__45916\,
            I => \N__45767\
        );

    \I__10402\ : InMux
    port map (
            O => \N__45915\,
            I => \N__45767\
        );

    \I__10401\ : InMux
    port map (
            O => \N__45912\,
            I => \N__45767\
        );

    \I__10400\ : InMux
    port map (
            O => \N__45911\,
            I => \N__45767\
        );

    \I__10399\ : CascadeMux
    port map (
            O => \N__45910\,
            I => \N__45764\
        );

    \I__10398\ : CascadeMux
    port map (
            O => \N__45909\,
            I => \N__45760\
        );

    \I__10397\ : CascadeMux
    port map (
            O => \N__45908\,
            I => \N__45756\
        );

    \I__10396\ : CascadeMux
    port map (
            O => \N__45907\,
            I => \N__45752\
        );

    \I__10395\ : CascadeMux
    port map (
            O => \N__45906\,
            I => \N__45744\
        );

    \I__10394\ : CascadeMux
    port map (
            O => \N__45905\,
            I => \N__45740\
        );

    \I__10393\ : CascadeMux
    port map (
            O => \N__45904\,
            I => \N__45736\
        );

    \I__10392\ : CascadeMux
    port map (
            O => \N__45903\,
            I => \N__45732\
        );

    \I__10391\ : CascadeMux
    port map (
            O => \N__45902\,
            I => \N__45728\
        );

    \I__10390\ : CascadeMux
    port map (
            O => \N__45901\,
            I => \N__45724\
        );

    \I__10389\ : CascadeMux
    port map (
            O => \N__45900\,
            I => \N__45720\
        );

    \I__10388\ : InMux
    port map (
            O => \N__45897\,
            I => \N__45706\
        );

    \I__10387\ : InMux
    port map (
            O => \N__45896\,
            I => \N__45706\
        );

    \I__10386\ : InMux
    port map (
            O => \N__45893\,
            I => \N__45706\
        );

    \I__10385\ : InMux
    port map (
            O => \N__45892\,
            I => \N__45706\
        );

    \I__10384\ : InMux
    port map (
            O => \N__45889\,
            I => \N__45706\
        );

    \I__10383\ : InMux
    port map (
            O => \N__45888\,
            I => \N__45706\
        );

    \I__10382\ : InMux
    port map (
            O => \N__45887\,
            I => \N__45697\
        );

    \I__10381\ : InMux
    port map (
            O => \N__45886\,
            I => \N__45697\
        );

    \I__10380\ : InMux
    port map (
            O => \N__45885\,
            I => \N__45697\
        );

    \I__10379\ : InMux
    port map (
            O => \N__45884\,
            I => \N__45697\
        );

    \I__10378\ : InMux
    port map (
            O => \N__45883\,
            I => \N__45692\
        );

    \I__10377\ : InMux
    port map (
            O => \N__45882\,
            I => \N__45692\
        );

    \I__10376\ : LocalMux
    port map (
            O => \N__45877\,
            I => \N__45689\
        );

    \I__10375\ : InMux
    port map (
            O => \N__45876\,
            I => \N__45686\
        );

    \I__10374\ : CascadeMux
    port map (
            O => \N__45875\,
            I => \N__45682\
        );

    \I__10373\ : CascadeMux
    port map (
            O => \N__45874\,
            I => \N__45676\
        );

    \I__10372\ : LocalMux
    port map (
            O => \N__45871\,
            I => \N__45667\
        );

    \I__10371\ : LocalMux
    port map (
            O => \N__45864\,
            I => \N__45667\
        );

    \I__10370\ : LocalMux
    port map (
            O => \N__45853\,
            I => \N__45664\
        );

    \I__10369\ : InMux
    port map (
            O => \N__45852\,
            I => \N__45653\
        );

    \I__10368\ : InMux
    port map (
            O => \N__45849\,
            I => \N__45653\
        );

    \I__10367\ : InMux
    port map (
            O => \N__45848\,
            I => \N__45653\
        );

    \I__10366\ : InMux
    port map (
            O => \N__45845\,
            I => \N__45653\
        );

    \I__10365\ : InMux
    port map (
            O => \N__45844\,
            I => \N__45653\
        );

    \I__10364\ : CascadeMux
    port map (
            O => \N__45843\,
            I => \N__45650\
        );

    \I__10363\ : CascadeMux
    port map (
            O => \N__45842\,
            I => \N__45646\
        );

    \I__10362\ : CascadeMux
    port map (
            O => \N__45841\,
            I => \N__45642\
        );

    \I__10361\ : CascadeMux
    port map (
            O => \N__45840\,
            I => \N__45638\
        );

    \I__10360\ : Span4Mux_v
    port map (
            O => \N__45835\,
            I => \N__45628\
        );

    \I__10359\ : LocalMux
    port map (
            O => \N__45822\,
            I => \N__45628\
        );

    \I__10358\ : LocalMux
    port map (
            O => \N__45811\,
            I => \N__45628\
        );

    \I__10357\ : LocalMux
    port map (
            O => \N__45806\,
            I => \N__45628\
        );

    \I__10356\ : InMux
    port map (
            O => \N__45805\,
            I => \N__45617\
        );

    \I__10355\ : InMux
    port map (
            O => \N__45804\,
            I => \N__45617\
        );

    \I__10354\ : InMux
    port map (
            O => \N__45803\,
            I => \N__45617\
        );

    \I__10353\ : InMux
    port map (
            O => \N__45802\,
            I => \N__45617\
        );

    \I__10352\ : InMux
    port map (
            O => \N__45801\,
            I => \N__45617\
        );

    \I__10351\ : LocalMux
    port map (
            O => \N__45784\,
            I => \N__45612\
        );

    \I__10350\ : LocalMux
    port map (
            O => \N__45767\,
            I => \N__45612\
        );

    \I__10349\ : InMux
    port map (
            O => \N__45764\,
            I => \N__45595\
        );

    \I__10348\ : InMux
    port map (
            O => \N__45763\,
            I => \N__45595\
        );

    \I__10347\ : InMux
    port map (
            O => \N__45760\,
            I => \N__45595\
        );

    \I__10346\ : InMux
    port map (
            O => \N__45759\,
            I => \N__45595\
        );

    \I__10345\ : InMux
    port map (
            O => \N__45756\,
            I => \N__45595\
        );

    \I__10344\ : InMux
    port map (
            O => \N__45755\,
            I => \N__45595\
        );

    \I__10343\ : InMux
    port map (
            O => \N__45752\,
            I => \N__45595\
        );

    \I__10342\ : InMux
    port map (
            O => \N__45751\,
            I => \N__45595\
        );

    \I__10341\ : CascadeMux
    port map (
            O => \N__45750\,
            I => \N__45592\
        );

    \I__10340\ : CascadeMux
    port map (
            O => \N__45749\,
            I => \N__45588\
        );

    \I__10339\ : CascadeMux
    port map (
            O => \N__45748\,
            I => \N__45584\
        );

    \I__10338\ : InMux
    port map (
            O => \N__45747\,
            I => \N__45568\
        );

    \I__10337\ : InMux
    port map (
            O => \N__45744\,
            I => \N__45568\
        );

    \I__10336\ : InMux
    port map (
            O => \N__45743\,
            I => \N__45568\
        );

    \I__10335\ : InMux
    port map (
            O => \N__45740\,
            I => \N__45568\
        );

    \I__10334\ : InMux
    port map (
            O => \N__45739\,
            I => \N__45568\
        );

    \I__10333\ : InMux
    port map (
            O => \N__45736\,
            I => \N__45568\
        );

    \I__10332\ : InMux
    port map (
            O => \N__45735\,
            I => \N__45568\
        );

    \I__10331\ : InMux
    port map (
            O => \N__45732\,
            I => \N__45551\
        );

    \I__10330\ : InMux
    port map (
            O => \N__45731\,
            I => \N__45551\
        );

    \I__10329\ : InMux
    port map (
            O => \N__45728\,
            I => \N__45551\
        );

    \I__10328\ : InMux
    port map (
            O => \N__45727\,
            I => \N__45551\
        );

    \I__10327\ : InMux
    port map (
            O => \N__45724\,
            I => \N__45551\
        );

    \I__10326\ : InMux
    port map (
            O => \N__45723\,
            I => \N__45551\
        );

    \I__10325\ : InMux
    port map (
            O => \N__45720\,
            I => \N__45551\
        );

    \I__10324\ : InMux
    port map (
            O => \N__45719\,
            I => \N__45551\
        );

    \I__10323\ : LocalMux
    port map (
            O => \N__45706\,
            I => \N__45548\
        );

    \I__10322\ : LocalMux
    port map (
            O => \N__45697\,
            I => \N__45543\
        );

    \I__10321\ : LocalMux
    port map (
            O => \N__45692\,
            I => \N__45543\
        );

    \I__10320\ : Span4Mux_h
    port map (
            O => \N__45689\,
            I => \N__45538\
        );

    \I__10319\ : LocalMux
    port map (
            O => \N__45686\,
            I => \N__45538\
        );

    \I__10318\ : InMux
    port map (
            O => \N__45685\,
            I => \N__45523\
        );

    \I__10317\ : InMux
    port map (
            O => \N__45682\,
            I => \N__45523\
        );

    \I__10316\ : InMux
    port map (
            O => \N__45681\,
            I => \N__45523\
        );

    \I__10315\ : InMux
    port map (
            O => \N__45680\,
            I => \N__45523\
        );

    \I__10314\ : InMux
    port map (
            O => \N__45679\,
            I => \N__45523\
        );

    \I__10313\ : InMux
    port map (
            O => \N__45676\,
            I => \N__45523\
        );

    \I__10312\ : InMux
    port map (
            O => \N__45675\,
            I => \N__45523\
        );

    \I__10311\ : InMux
    port map (
            O => \N__45674\,
            I => \N__45516\
        );

    \I__10310\ : InMux
    port map (
            O => \N__45673\,
            I => \N__45516\
        );

    \I__10309\ : InMux
    port map (
            O => \N__45672\,
            I => \N__45516\
        );

    \I__10308\ : Span4Mux_v
    port map (
            O => \N__45667\,
            I => \N__45509\
        );

    \I__10307\ : Span4Mux_v
    port map (
            O => \N__45664\,
            I => \N__45509\
        );

    \I__10306\ : LocalMux
    port map (
            O => \N__45653\,
            I => \N__45509\
        );

    \I__10305\ : InMux
    port map (
            O => \N__45650\,
            I => \N__45492\
        );

    \I__10304\ : InMux
    port map (
            O => \N__45649\,
            I => \N__45492\
        );

    \I__10303\ : InMux
    port map (
            O => \N__45646\,
            I => \N__45492\
        );

    \I__10302\ : InMux
    port map (
            O => \N__45645\,
            I => \N__45492\
        );

    \I__10301\ : InMux
    port map (
            O => \N__45642\,
            I => \N__45492\
        );

    \I__10300\ : InMux
    port map (
            O => \N__45641\,
            I => \N__45492\
        );

    \I__10299\ : InMux
    port map (
            O => \N__45638\,
            I => \N__45492\
        );

    \I__10298\ : InMux
    port map (
            O => \N__45637\,
            I => \N__45492\
        );

    \I__10297\ : Span4Mux_v
    port map (
            O => \N__45628\,
            I => \N__45483\
        );

    \I__10296\ : LocalMux
    port map (
            O => \N__45617\,
            I => \N__45483\
        );

    \I__10295\ : Span4Mux_v
    port map (
            O => \N__45612\,
            I => \N__45483\
        );

    \I__10294\ : LocalMux
    port map (
            O => \N__45595\,
            I => \N__45483\
        );

    \I__10293\ : InMux
    port map (
            O => \N__45592\,
            I => \N__45470\
        );

    \I__10292\ : InMux
    port map (
            O => \N__45591\,
            I => \N__45470\
        );

    \I__10291\ : InMux
    port map (
            O => \N__45588\,
            I => \N__45470\
        );

    \I__10290\ : InMux
    port map (
            O => \N__45587\,
            I => \N__45470\
        );

    \I__10289\ : InMux
    port map (
            O => \N__45584\,
            I => \N__45470\
        );

    \I__10288\ : InMux
    port map (
            O => \N__45583\,
            I => \N__45470\
        );

    \I__10287\ : LocalMux
    port map (
            O => \N__45568\,
            I => \N__45463\
        );

    \I__10286\ : LocalMux
    port map (
            O => \N__45551\,
            I => \N__45463\
        );

    \I__10285\ : Span4Mux_h
    port map (
            O => \N__45548\,
            I => \N__45463\
        );

    \I__10284\ : Odrv12
    port map (
            O => \N__45543\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10283\ : Odrv4
    port map (
            O => \N__45538\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10282\ : LocalMux
    port map (
            O => \N__45523\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10281\ : LocalMux
    port map (
            O => \N__45516\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10280\ : Odrv4
    port map (
            O => \N__45509\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10279\ : LocalMux
    port map (
            O => \N__45492\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10278\ : Odrv4
    port map (
            O => \N__45483\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10277\ : LocalMux
    port map (
            O => \N__45470\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10276\ : Odrv4
    port map (
            O => \N__45463\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10275\ : CascadeMux
    port map (
            O => \N__45444\,
            I => \N__45400\
        );

    \I__10274\ : InMux
    port map (
            O => \N__45443\,
            I => \N__45389\
        );

    \I__10273\ : InMux
    port map (
            O => \N__45442\,
            I => \N__45378\
        );

    \I__10272\ : InMux
    port map (
            O => \N__45441\,
            I => \N__45378\
        );

    \I__10271\ : InMux
    port map (
            O => \N__45440\,
            I => \N__45378\
        );

    \I__10270\ : InMux
    port map (
            O => \N__45439\,
            I => \N__45378\
        );

    \I__10269\ : InMux
    port map (
            O => \N__45438\,
            I => \N__45378\
        );

    \I__10268\ : InMux
    port map (
            O => \N__45437\,
            I => \N__45365\
        );

    \I__10267\ : InMux
    port map (
            O => \N__45436\,
            I => \N__45365\
        );

    \I__10266\ : InMux
    port map (
            O => \N__45435\,
            I => \N__45365\
        );

    \I__10265\ : InMux
    port map (
            O => \N__45434\,
            I => \N__45365\
        );

    \I__10264\ : InMux
    port map (
            O => \N__45433\,
            I => \N__45365\
        );

    \I__10263\ : InMux
    port map (
            O => \N__45432\,
            I => \N__45365\
        );

    \I__10262\ : InMux
    port map (
            O => \N__45431\,
            I => \N__45355\
        );

    \I__10261\ : InMux
    port map (
            O => \N__45430\,
            I => \N__45355\
        );

    \I__10260\ : InMux
    port map (
            O => \N__45429\,
            I => \N__45355\
        );

    \I__10259\ : InMux
    port map (
            O => \N__45428\,
            I => \N__45355\
        );

    \I__10258\ : InMux
    port map (
            O => \N__45427\,
            I => \N__45346\
        );

    \I__10257\ : InMux
    port map (
            O => \N__45426\,
            I => \N__45346\
        );

    \I__10256\ : InMux
    port map (
            O => \N__45425\,
            I => \N__45346\
        );

    \I__10255\ : InMux
    port map (
            O => \N__45424\,
            I => \N__45346\
        );

    \I__10254\ : InMux
    port map (
            O => \N__45423\,
            I => \N__45333\
        );

    \I__10253\ : InMux
    port map (
            O => \N__45422\,
            I => \N__45333\
        );

    \I__10252\ : InMux
    port map (
            O => \N__45421\,
            I => \N__45324\
        );

    \I__10251\ : InMux
    port map (
            O => \N__45420\,
            I => \N__45324\
        );

    \I__10250\ : InMux
    port map (
            O => \N__45419\,
            I => \N__45324\
        );

    \I__10249\ : InMux
    port map (
            O => \N__45418\,
            I => \N__45324\
        );

    \I__10248\ : InMux
    port map (
            O => \N__45417\,
            I => \N__45313\
        );

    \I__10247\ : InMux
    port map (
            O => \N__45416\,
            I => \N__45313\
        );

    \I__10246\ : InMux
    port map (
            O => \N__45415\,
            I => \N__45313\
        );

    \I__10245\ : InMux
    port map (
            O => \N__45414\,
            I => \N__45313\
        );

    \I__10244\ : InMux
    port map (
            O => \N__45413\,
            I => \N__45313\
        );

    \I__10243\ : InMux
    port map (
            O => \N__45412\,
            I => \N__45306\
        );

    \I__10242\ : InMux
    port map (
            O => \N__45411\,
            I => \N__45306\
        );

    \I__10241\ : InMux
    port map (
            O => \N__45410\,
            I => \N__45306\
        );

    \I__10240\ : InMux
    port map (
            O => \N__45409\,
            I => \N__45303\
        );

    \I__10239\ : InMux
    port map (
            O => \N__45408\,
            I => \N__45286\
        );

    \I__10238\ : InMux
    port map (
            O => \N__45407\,
            I => \N__45286\
        );

    \I__10237\ : InMux
    port map (
            O => \N__45406\,
            I => \N__45286\
        );

    \I__10236\ : InMux
    port map (
            O => \N__45405\,
            I => \N__45286\
        );

    \I__10235\ : InMux
    port map (
            O => \N__45404\,
            I => \N__45286\
        );

    \I__10234\ : InMux
    port map (
            O => \N__45403\,
            I => \N__45283\
        );

    \I__10233\ : InMux
    port map (
            O => \N__45400\,
            I => \N__45268\
        );

    \I__10232\ : InMux
    port map (
            O => \N__45399\,
            I => \N__45268\
        );

    \I__10231\ : InMux
    port map (
            O => \N__45398\,
            I => \N__45268\
        );

    \I__10230\ : InMux
    port map (
            O => \N__45397\,
            I => \N__45268\
        );

    \I__10229\ : InMux
    port map (
            O => \N__45396\,
            I => \N__45268\
        );

    \I__10228\ : InMux
    port map (
            O => \N__45395\,
            I => \N__45268\
        );

    \I__10227\ : InMux
    port map (
            O => \N__45394\,
            I => \N__45268\
        );

    \I__10226\ : InMux
    port map (
            O => \N__45393\,
            I => \N__45263\
        );

    \I__10225\ : InMux
    port map (
            O => \N__45392\,
            I => \N__45260\
        );

    \I__10224\ : LocalMux
    port map (
            O => \N__45389\,
            I => \N__45257\
        );

    \I__10223\ : LocalMux
    port map (
            O => \N__45378\,
            I => \N__45252\
        );

    \I__10222\ : LocalMux
    port map (
            O => \N__45365\,
            I => \N__45252\
        );

    \I__10221\ : CascadeMux
    port map (
            O => \N__45364\,
            I => \N__45246\
        );

    \I__10220\ : LocalMux
    port map (
            O => \N__45355\,
            I => \N__45242\
        );

    \I__10219\ : LocalMux
    port map (
            O => \N__45346\,
            I => \N__45239\
        );

    \I__10218\ : InMux
    port map (
            O => \N__45345\,
            I => \N__45236\
        );

    \I__10217\ : InMux
    port map (
            O => \N__45344\,
            I => \N__45221\
        );

    \I__10216\ : InMux
    port map (
            O => \N__45343\,
            I => \N__45221\
        );

    \I__10215\ : InMux
    port map (
            O => \N__45342\,
            I => \N__45221\
        );

    \I__10214\ : InMux
    port map (
            O => \N__45341\,
            I => \N__45221\
        );

    \I__10213\ : InMux
    port map (
            O => \N__45340\,
            I => \N__45221\
        );

    \I__10212\ : InMux
    port map (
            O => \N__45339\,
            I => \N__45221\
        );

    \I__10211\ : InMux
    port map (
            O => \N__45338\,
            I => \N__45221\
        );

    \I__10210\ : LocalMux
    port map (
            O => \N__45333\,
            I => \N__45216\
        );

    \I__10209\ : LocalMux
    port map (
            O => \N__45324\,
            I => \N__45216\
        );

    \I__10208\ : LocalMux
    port map (
            O => \N__45313\,
            I => \N__45213\
        );

    \I__10207\ : LocalMux
    port map (
            O => \N__45306\,
            I => \N__45208\
        );

    \I__10206\ : LocalMux
    port map (
            O => \N__45303\,
            I => \N__45208\
        );

    \I__10205\ : InMux
    port map (
            O => \N__45302\,
            I => \N__45195\
        );

    \I__10204\ : InMux
    port map (
            O => \N__45301\,
            I => \N__45195\
        );

    \I__10203\ : InMux
    port map (
            O => \N__45300\,
            I => \N__45195\
        );

    \I__10202\ : InMux
    port map (
            O => \N__45299\,
            I => \N__45195\
        );

    \I__10201\ : InMux
    port map (
            O => \N__45298\,
            I => \N__45195\
        );

    \I__10200\ : InMux
    port map (
            O => \N__45297\,
            I => \N__45195\
        );

    \I__10199\ : LocalMux
    port map (
            O => \N__45286\,
            I => \N__45192\
        );

    \I__10198\ : LocalMux
    port map (
            O => \N__45283\,
            I => \N__45187\
        );

    \I__10197\ : LocalMux
    port map (
            O => \N__45268\,
            I => \N__45187\
        );

    \I__10196\ : InMux
    port map (
            O => \N__45267\,
            I => \N__45182\
        );

    \I__10195\ : InMux
    port map (
            O => \N__45266\,
            I => \N__45182\
        );

    \I__10194\ : LocalMux
    port map (
            O => \N__45263\,
            I => \N__45173\
        );

    \I__10193\ : LocalMux
    port map (
            O => \N__45260\,
            I => \N__45173\
        );

    \I__10192\ : Span4Mux_v
    port map (
            O => \N__45257\,
            I => \N__45173\
        );

    \I__10191\ : Span4Mux_v
    port map (
            O => \N__45252\,
            I => \N__45173\
        );

    \I__10190\ : InMux
    port map (
            O => \N__45251\,
            I => \N__45162\
        );

    \I__10189\ : InMux
    port map (
            O => \N__45250\,
            I => \N__45162\
        );

    \I__10188\ : InMux
    port map (
            O => \N__45249\,
            I => \N__45162\
        );

    \I__10187\ : InMux
    port map (
            O => \N__45246\,
            I => \N__45162\
        );

    \I__10186\ : InMux
    port map (
            O => \N__45245\,
            I => \N__45162\
        );

    \I__10185\ : Span4Mux_h
    port map (
            O => \N__45242\,
            I => \N__45159\
        );

    \I__10184\ : Span4Mux_v
    port map (
            O => \N__45239\,
            I => \N__45156\
        );

    \I__10183\ : LocalMux
    port map (
            O => \N__45236\,
            I => \N__45145\
        );

    \I__10182\ : LocalMux
    port map (
            O => \N__45221\,
            I => \N__45145\
        );

    \I__10181\ : Span4Mux_v
    port map (
            O => \N__45216\,
            I => \N__45145\
        );

    \I__10180\ : Span4Mux_h
    port map (
            O => \N__45213\,
            I => \N__45145\
        );

    \I__10179\ : Span4Mux_v
    port map (
            O => \N__45208\,
            I => \N__45145\
        );

    \I__10178\ : LocalMux
    port map (
            O => \N__45195\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10177\ : Odrv4
    port map (
            O => \N__45192\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10176\ : Odrv4
    port map (
            O => \N__45187\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10175\ : LocalMux
    port map (
            O => \N__45182\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10174\ : Odrv4
    port map (
            O => \N__45173\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10173\ : LocalMux
    port map (
            O => \N__45162\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10172\ : Odrv4
    port map (
            O => \N__45159\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10171\ : Odrv4
    port map (
            O => \N__45156\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10170\ : Odrv4
    port map (
            O => \N__45145\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10169\ : CascadeMux
    port map (
            O => \N__45126\,
            I => \N__45123\
        );

    \I__10168\ : InMux
    port map (
            O => \N__45123\,
            I => \N__45119\
        );

    \I__10167\ : CascadeMux
    port map (
            O => \N__45122\,
            I => \N__45116\
        );

    \I__10166\ : LocalMux
    port map (
            O => \N__45119\,
            I => \N__45112\
        );

    \I__10165\ : InMux
    port map (
            O => \N__45116\,
            I => \N__45107\
        );

    \I__10164\ : InMux
    port map (
            O => \N__45115\,
            I => \N__45107\
        );

    \I__10163\ : Odrv4
    port map (
            O => \N__45112\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__10162\ : LocalMux
    port map (
            O => \N__45107\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__10161\ : InMux
    port map (
            O => \N__45102\,
            I => \N__45096\
        );

    \I__10160\ : InMux
    port map (
            O => \N__45101\,
            I => \N__45096\
        );

    \I__10159\ : LocalMux
    port map (
            O => \N__45096\,
            I => \N__45091\
        );

    \I__10158\ : InMux
    port map (
            O => \N__45095\,
            I => \N__45086\
        );

    \I__10157\ : InMux
    port map (
            O => \N__45094\,
            I => \N__45086\
        );

    \I__10156\ : Span4Mux_h
    port map (
            O => \N__45091\,
            I => \N__45083\
        );

    \I__10155\ : LocalMux
    port map (
            O => \N__45086\,
            I => \N__45080\
        );

    \I__10154\ : Span4Mux_h
    port map (
            O => \N__45083\,
            I => \N__45077\
        );

    \I__10153\ : Odrv4
    port map (
            O => \N__45080\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__10152\ : Odrv4
    port map (
            O => \N__45077\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__10151\ : CascadeMux
    port map (
            O => \N__45072\,
            I => \N__45069\
        );

    \I__10150\ : InMux
    port map (
            O => \N__45069\,
            I => \N__45066\
        );

    \I__10149\ : LocalMux
    port map (
            O => \N__45066\,
            I => \N__45063\
        );

    \I__10148\ : Span4Mux_h
    port map (
            O => \N__45063\,
            I => \N__45060\
        );

    \I__10147\ : Odrv4
    port map (
            O => \N__45060\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\
        );

    \I__10146\ : InMux
    port map (
            O => \N__45057\,
            I => \N__45054\
        );

    \I__10145\ : LocalMux
    port map (
            O => \N__45054\,
            I => \N__45051\
        );

    \I__10144\ : Span4Mux_h
    port map (
            O => \N__45051\,
            I => \N__45048\
        );

    \I__10143\ : Span4Mux_v
    port map (
            O => \N__45048\,
            I => \N__45045\
        );

    \I__10142\ : Odrv4
    port map (
            O => \N__45045\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\
        );

    \I__10141\ : CascadeMux
    port map (
            O => \N__45042\,
            I => \N__45039\
        );

    \I__10140\ : InMux
    port map (
            O => \N__45039\,
            I => \N__45036\
        );

    \I__10139\ : LocalMux
    port map (
            O => \N__45036\,
            I => \N__45033\
        );

    \I__10138\ : Span4Mux_v
    port map (
            O => \N__45033\,
            I => \N__45029\
        );

    \I__10137\ : InMux
    port map (
            O => \N__45032\,
            I => \N__45026\
        );

    \I__10136\ : Odrv4
    port map (
            O => \N__45029\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__10135\ : LocalMux
    port map (
            O => \N__45026\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__10134\ : InMux
    port map (
            O => \N__45021\,
            I => \N__45018\
        );

    \I__10133\ : LocalMux
    port map (
            O => \N__45018\,
            I => \N__45015\
        );

    \I__10132\ : Span4Mux_h
    port map (
            O => \N__45015\,
            I => \N__45012\
        );

    \I__10131\ : Span4Mux_h
    port map (
            O => \N__45012\,
            I => \N__45009\
        );

    \I__10130\ : Odrv4
    port map (
            O => \N__45009\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\
        );

    \I__10129\ : CascadeMux
    port map (
            O => \N__45006\,
            I => \N__45003\
        );

    \I__10128\ : InMux
    port map (
            O => \N__45003\,
            I => \N__44999\
        );

    \I__10127\ : CascadeMux
    port map (
            O => \N__45002\,
            I => \N__44995\
        );

    \I__10126\ : LocalMux
    port map (
            O => \N__44999\,
            I => \N__44991\
        );

    \I__10125\ : InMux
    port map (
            O => \N__44998\,
            I => \N__44988\
        );

    \I__10124\ : InMux
    port map (
            O => \N__44995\,
            I => \N__44985\
        );

    \I__10123\ : InMux
    port map (
            O => \N__44994\,
            I => \N__44982\
        );

    \I__10122\ : Span4Mux_v
    port map (
            O => \N__44991\,
            I => \N__44977\
        );

    \I__10121\ : LocalMux
    port map (
            O => \N__44988\,
            I => \N__44977\
        );

    \I__10120\ : LocalMux
    port map (
            O => \N__44985\,
            I => \N__44974\
        );

    \I__10119\ : LocalMux
    port map (
            O => \N__44982\,
            I => \N__44969\
        );

    \I__10118\ : Span4Mux_v
    port map (
            O => \N__44977\,
            I => \N__44969\
        );

    \I__10117\ : Odrv12
    port map (
            O => \N__44974\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10116\ : Odrv4
    port map (
            O => \N__44969\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10115\ : InMux
    port map (
            O => \N__44964\,
            I => \N__44961\
        );

    \I__10114\ : LocalMux
    port map (
            O => \N__44961\,
            I => \N__44958\
        );

    \I__10113\ : Span4Mux_v
    port map (
            O => \N__44958\,
            I => \N__44953\
        );

    \I__10112\ : InMux
    port map (
            O => \N__44957\,
            I => \N__44950\
        );

    \I__10111\ : InMux
    port map (
            O => \N__44956\,
            I => \N__44947\
        );

    \I__10110\ : Odrv4
    port map (
            O => \N__44953\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__10109\ : LocalMux
    port map (
            O => \N__44950\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__10108\ : LocalMux
    port map (
            O => \N__44947\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__10107\ : InMux
    port map (
            O => \N__44940\,
            I => \N__44937\
        );

    \I__10106\ : LocalMux
    port map (
            O => \N__44937\,
            I => \N__44934\
        );

    \I__10105\ : Span4Mux_v
    port map (
            O => \N__44934\,
            I => \N__44931\
        );

    \I__10104\ : Odrv4
    port map (
            O => \N__44931\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\
        );

    \I__10103\ : InMux
    port map (
            O => \N__44928\,
            I => \N__44925\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__44925\,
            I => \N__44921\
        );

    \I__10101\ : InMux
    port map (
            O => \N__44924\,
            I => \N__44918\
        );

    \I__10100\ : Sp12to4
    port map (
            O => \N__44921\,
            I => \N__44912\
        );

    \I__10099\ : LocalMux
    port map (
            O => \N__44918\,
            I => \N__44912\
        );

    \I__10098\ : InMux
    port map (
            O => \N__44917\,
            I => \N__44909\
        );

    \I__10097\ : Span12Mux_v
    port map (
            O => \N__44912\,
            I => \N__44906\
        );

    \I__10096\ : LocalMux
    port map (
            O => \N__44909\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\
        );

    \I__10095\ : Odrv12
    port map (
            O => \N__44906\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\
        );

    \I__10094\ : InMux
    port map (
            O => \N__44901\,
            I => \N__44893\
        );

    \I__10093\ : InMux
    port map (
            O => \N__44900\,
            I => \N__44893\
        );

    \I__10092\ : InMux
    port map (
            O => \N__44899\,
            I => \N__44890\
        );

    \I__10091\ : InMux
    port map (
            O => \N__44898\,
            I => \N__44887\
        );

    \I__10090\ : LocalMux
    port map (
            O => \N__44893\,
            I => \N__44884\
        );

    \I__10089\ : LocalMux
    port map (
            O => \N__44890\,
            I => \N__44881\
        );

    \I__10088\ : LocalMux
    port map (
            O => \N__44887\,
            I => \N__44878\
        );

    \I__10087\ : Span4Mux_v
    port map (
            O => \N__44884\,
            I => \N__44875\
        );

    \I__10086\ : Span12Mux_s9_v
    port map (
            O => \N__44881\,
            I => \N__44872\
        );

    \I__10085\ : Span4Mux_h
    port map (
            O => \N__44878\,
            I => \N__44869\
        );

    \I__10084\ : Odrv4
    port map (
            O => \N__44875\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__10083\ : Odrv12
    port map (
            O => \N__44872\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__10082\ : Odrv4
    port map (
            O => \N__44869\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__10081\ : CascadeMux
    port map (
            O => \N__44862\,
            I => \N__44859\
        );

    \I__10080\ : InMux
    port map (
            O => \N__44859\,
            I => \N__44852\
        );

    \I__10079\ : InMux
    port map (
            O => \N__44858\,
            I => \N__44852\
        );

    \I__10078\ : InMux
    port map (
            O => \N__44857\,
            I => \N__44849\
        );

    \I__10077\ : LocalMux
    port map (
            O => \N__44852\,
            I => \N__44846\
        );

    \I__10076\ : LocalMux
    port map (
            O => \N__44849\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__10075\ : Odrv4
    port map (
            O => \N__44846\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__10074\ : InMux
    port map (
            O => \N__44841\,
            I => \N__44838\
        );

    \I__10073\ : LocalMux
    port map (
            O => \N__44838\,
            I => \N__44835\
        );

    \I__10072\ : Span4Mux_v
    port map (
            O => \N__44835\,
            I => \N__44832\
        );

    \I__10071\ : Odrv4
    port map (
            O => \N__44832\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\
        );

    \I__10070\ : CascadeMux
    port map (
            O => \N__44829\,
            I => \N__44826\
        );

    \I__10069\ : InMux
    port map (
            O => \N__44826\,
            I => \N__44822\
        );

    \I__10068\ : CascadeMux
    port map (
            O => \N__44825\,
            I => \N__44819\
        );

    \I__10067\ : LocalMux
    port map (
            O => \N__44822\,
            I => \N__44816\
        );

    \I__10066\ : InMux
    port map (
            O => \N__44819\,
            I => \N__44813\
        );

    \I__10065\ : Span4Mux_h
    port map (
            O => \N__44816\,
            I => \N__44809\
        );

    \I__10064\ : LocalMux
    port map (
            O => \N__44813\,
            I => \N__44806\
        );

    \I__10063\ : CascadeMux
    port map (
            O => \N__44812\,
            I => \N__44803\
        );

    \I__10062\ : Span4Mux_v
    port map (
            O => \N__44809\,
            I => \N__44797\
        );

    \I__10061\ : Span4Mux_h
    port map (
            O => \N__44806\,
            I => \N__44797\
        );

    \I__10060\ : InMux
    port map (
            O => \N__44803\,
            I => \N__44792\
        );

    \I__10059\ : InMux
    port map (
            O => \N__44802\,
            I => \N__44792\
        );

    \I__10058\ : Span4Mux_h
    port map (
            O => \N__44797\,
            I => \N__44789\
        );

    \I__10057\ : LocalMux
    port map (
            O => \N__44792\,
            I => \N__44786\
        );

    \I__10056\ : Odrv4
    port map (
            O => \N__44789\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__10055\ : Odrv4
    port map (
            O => \N__44786\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__10054\ : InMux
    port map (
            O => \N__44781\,
            I => \N__44778\
        );

    \I__10053\ : LocalMux
    port map (
            O => \N__44778\,
            I => \N__44775\
        );

    \I__10052\ : Span4Mux_v
    port map (
            O => \N__44775\,
            I => \N__44770\
        );

    \I__10051\ : InMux
    port map (
            O => \N__44774\,
            I => \N__44767\
        );

    \I__10050\ : InMux
    port map (
            O => \N__44773\,
            I => \N__44764\
        );

    \I__10049\ : Odrv4
    port map (
            O => \N__44770\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__10048\ : LocalMux
    port map (
            O => \N__44767\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__10047\ : LocalMux
    port map (
            O => \N__44764\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__10046\ : CascadeMux
    port map (
            O => \N__44757\,
            I => \N__44754\
        );

    \I__10045\ : InMux
    port map (
            O => \N__44754\,
            I => \N__44751\
        );

    \I__10044\ : LocalMux
    port map (
            O => \N__44751\,
            I => \N__44748\
        );

    \I__10043\ : Odrv4
    port map (
            O => \N__44748\,
            I => \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\
        );

    \I__10042\ : InMux
    port map (
            O => \N__44745\,
            I => \N__44742\
        );

    \I__10041\ : LocalMux
    port map (
            O => \N__44742\,
            I => \N__44737\
        );

    \I__10040\ : InMux
    port map (
            O => \N__44741\,
            I => \N__44734\
        );

    \I__10039\ : InMux
    port map (
            O => \N__44740\,
            I => \N__44729\
        );

    \I__10038\ : Span4Mux_v
    port map (
            O => \N__44737\,
            I => \N__44726\
        );

    \I__10037\ : LocalMux
    port map (
            O => \N__44734\,
            I => \N__44723\
        );

    \I__10036\ : InMux
    port map (
            O => \N__44733\,
            I => \N__44718\
        );

    \I__10035\ : InMux
    port map (
            O => \N__44732\,
            I => \N__44718\
        );

    \I__10034\ : LocalMux
    port map (
            O => \N__44729\,
            I => \N__44715\
        );

    \I__10033\ : Span4Mux_h
    port map (
            O => \N__44726\,
            I => \N__44712\
        );

    \I__10032\ : Span4Mux_h
    port map (
            O => \N__44723\,
            I => \N__44709\
        );

    \I__10031\ : LocalMux
    port map (
            O => \N__44718\,
            I => \N__44706\
        );

    \I__10030\ : Span4Mux_v
    port map (
            O => \N__44715\,
            I => \N__44701\
        );

    \I__10029\ : Span4Mux_h
    port map (
            O => \N__44712\,
            I => \N__44701\
        );

    \I__10028\ : Odrv4
    port map (
            O => \N__44709\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__10027\ : Odrv4
    port map (
            O => \N__44706\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__10026\ : Odrv4
    port map (
            O => \N__44701\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__10025\ : InMux
    port map (
            O => \N__44694\,
            I => \N__44691\
        );

    \I__10024\ : LocalMux
    port map (
            O => \N__44691\,
            I => \N__44688\
        );

    \I__10023\ : Span4Mux_h
    port map (
            O => \N__44688\,
            I => \N__44685\
        );

    \I__10022\ : Span4Mux_h
    port map (
            O => \N__44685\,
            I => \N__44682\
        );

    \I__10021\ : Span4Mux_h
    port map (
            O => \N__44682\,
            I => \N__44679\
        );

    \I__10020\ : Odrv4
    port map (
            O => \N__44679\,
            I => \current_shift_inst.PI_CTRL.integrator_i_25\
        );

    \I__10019\ : CascadeMux
    port map (
            O => \N__44676\,
            I => \N__44672\
        );

    \I__10018\ : CascadeMux
    port map (
            O => \N__44675\,
            I => \N__44668\
        );

    \I__10017\ : InMux
    port map (
            O => \N__44672\,
            I => \N__44665\
        );

    \I__10016\ : InMux
    port map (
            O => \N__44671\,
            I => \N__44662\
        );

    \I__10015\ : InMux
    port map (
            O => \N__44668\,
            I => \N__44659\
        );

    \I__10014\ : LocalMux
    port map (
            O => \N__44665\,
            I => \N__44656\
        );

    \I__10013\ : LocalMux
    port map (
            O => \N__44662\,
            I => \N__44653\
        );

    \I__10012\ : LocalMux
    port map (
            O => \N__44659\,
            I => \N__44649\
        );

    \I__10011\ : Span4Mux_v
    port map (
            O => \N__44656\,
            I => \N__44644\
        );

    \I__10010\ : Span4Mux_h
    port map (
            O => \N__44653\,
            I => \N__44644\
        );

    \I__10009\ : InMux
    port map (
            O => \N__44652\,
            I => \N__44641\
        );

    \I__10008\ : Odrv12
    port map (
            O => \N__44649\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__10007\ : Odrv4
    port map (
            O => \N__44644\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__10006\ : LocalMux
    port map (
            O => \N__44641\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__10005\ : InMux
    port map (
            O => \N__44634\,
            I => \N__44631\
        );

    \I__10004\ : LocalMux
    port map (
            O => \N__44631\,
            I => \N__44628\
        );

    \I__10003\ : Span4Mux_h
    port map (
            O => \N__44628\,
            I => \N__44623\
        );

    \I__10002\ : InMux
    port map (
            O => \N__44627\,
            I => \N__44620\
        );

    \I__10001\ : InMux
    port map (
            O => \N__44626\,
            I => \N__44617\
        );

    \I__10000\ : Odrv4
    port map (
            O => \N__44623\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__9999\ : LocalMux
    port map (
            O => \N__44620\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__9998\ : LocalMux
    port map (
            O => \N__44617\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__9997\ : InMux
    port map (
            O => \N__44610\,
            I => \N__44607\
        );

    \I__9996\ : LocalMux
    port map (
            O => \N__44607\,
            I => \N__44604\
        );

    \I__9995\ : Span4Mux_v
    port map (
            O => \N__44604\,
            I => \N__44601\
        );

    \I__9994\ : Odrv4
    port map (
            O => \N__44601\,
            I => \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\
        );

    \I__9993\ : CascadeMux
    port map (
            O => \N__44598\,
            I => \N__44577\
        );

    \I__9992\ : CascadeMux
    port map (
            O => \N__44597\,
            I => \N__44571\
        );

    \I__9991\ : CascadeMux
    port map (
            O => \N__44596\,
            I => \N__44566\
        );

    \I__9990\ : InMux
    port map (
            O => \N__44595\,
            I => \N__44560\
        );

    \I__9989\ : InMux
    port map (
            O => \N__44594\,
            I => \N__44560\
        );

    \I__9988\ : CascadeMux
    port map (
            O => \N__44593\,
            I => \N__44556\
        );

    \I__9987\ : CascadeMux
    port map (
            O => \N__44592\,
            I => \N__44551\
        );

    \I__9986\ : CascadeMux
    port map (
            O => \N__44591\,
            I => \N__44548\
        );

    \I__9985\ : CascadeMux
    port map (
            O => \N__44590\,
            I => \N__44545\
        );

    \I__9984\ : InMux
    port map (
            O => \N__44589\,
            I => \N__44542\
        );

    \I__9983\ : InMux
    port map (
            O => \N__44588\,
            I => \N__44539\
        );

    \I__9982\ : InMux
    port map (
            O => \N__44587\,
            I => \N__44536\
        );

    \I__9981\ : InMux
    port map (
            O => \N__44586\,
            I => \N__44532\
        );

    \I__9980\ : CascadeMux
    port map (
            O => \N__44585\,
            I => \N__44528\
        );

    \I__9979\ : CascadeMux
    port map (
            O => \N__44584\,
            I => \N__44525\
        );

    \I__9978\ : CascadeMux
    port map (
            O => \N__44583\,
            I => \N__44519\
        );

    \I__9977\ : InMux
    port map (
            O => \N__44582\,
            I => \N__44505\
        );

    \I__9976\ : InMux
    port map (
            O => \N__44581\,
            I => \N__44505\
        );

    \I__9975\ : InMux
    port map (
            O => \N__44580\,
            I => \N__44502\
        );

    \I__9974\ : InMux
    port map (
            O => \N__44577\,
            I => \N__44499\
        );

    \I__9973\ : InMux
    port map (
            O => \N__44576\,
            I => \N__44496\
        );

    \I__9972\ : InMux
    port map (
            O => \N__44575\,
            I => \N__44492\
        );

    \I__9971\ : InMux
    port map (
            O => \N__44574\,
            I => \N__44481\
        );

    \I__9970\ : InMux
    port map (
            O => \N__44571\,
            I => \N__44481\
        );

    \I__9969\ : InMux
    port map (
            O => \N__44570\,
            I => \N__44481\
        );

    \I__9968\ : InMux
    port map (
            O => \N__44569\,
            I => \N__44481\
        );

    \I__9967\ : InMux
    port map (
            O => \N__44566\,
            I => \N__44481\
        );

    \I__9966\ : InMux
    port map (
            O => \N__44565\,
            I => \N__44478\
        );

    \I__9965\ : LocalMux
    port map (
            O => \N__44560\,
            I => \N__44475\
        );

    \I__9964\ : InMux
    port map (
            O => \N__44559\,
            I => \N__44461\
        );

    \I__9963\ : InMux
    port map (
            O => \N__44556\,
            I => \N__44461\
        );

    \I__9962\ : InMux
    port map (
            O => \N__44555\,
            I => \N__44461\
        );

    \I__9961\ : InMux
    port map (
            O => \N__44554\,
            I => \N__44461\
        );

    \I__9960\ : InMux
    port map (
            O => \N__44551\,
            I => \N__44461\
        );

    \I__9959\ : InMux
    port map (
            O => \N__44548\,
            I => \N__44461\
        );

    \I__9958\ : InMux
    port map (
            O => \N__44545\,
            I => \N__44458\
        );

    \I__9957\ : LocalMux
    port map (
            O => \N__44542\,
            I => \N__44453\
        );

    \I__9956\ : LocalMux
    port map (
            O => \N__44539\,
            I => \N__44453\
        );

    \I__9955\ : LocalMux
    port map (
            O => \N__44536\,
            I => \N__44450\
        );

    \I__9954\ : InMux
    port map (
            O => \N__44535\,
            I => \N__44447\
        );

    \I__9953\ : LocalMux
    port map (
            O => \N__44532\,
            I => \N__44444\
        );

    \I__9952\ : InMux
    port map (
            O => \N__44531\,
            I => \N__44427\
        );

    \I__9951\ : InMux
    port map (
            O => \N__44528\,
            I => \N__44427\
        );

    \I__9950\ : InMux
    port map (
            O => \N__44525\,
            I => \N__44427\
        );

    \I__9949\ : InMux
    port map (
            O => \N__44524\,
            I => \N__44427\
        );

    \I__9948\ : InMux
    port map (
            O => \N__44523\,
            I => \N__44427\
        );

    \I__9947\ : InMux
    port map (
            O => \N__44522\,
            I => \N__44427\
        );

    \I__9946\ : InMux
    port map (
            O => \N__44519\,
            I => \N__44427\
        );

    \I__9945\ : InMux
    port map (
            O => \N__44518\,
            I => \N__44427\
        );

    \I__9944\ : InMux
    port map (
            O => \N__44517\,
            I => \N__44420\
        );

    \I__9943\ : InMux
    port map (
            O => \N__44516\,
            I => \N__44420\
        );

    \I__9942\ : InMux
    port map (
            O => \N__44515\,
            I => \N__44420\
        );

    \I__9941\ : InMux
    port map (
            O => \N__44514\,
            I => \N__44417\
        );

    \I__9940\ : InMux
    port map (
            O => \N__44513\,
            I => \N__44414\
        );

    \I__9939\ : InMux
    port map (
            O => \N__44512\,
            I => \N__44407\
        );

    \I__9938\ : InMux
    port map (
            O => \N__44511\,
            I => \N__44407\
        );

    \I__9937\ : InMux
    port map (
            O => \N__44510\,
            I => \N__44407\
        );

    \I__9936\ : LocalMux
    port map (
            O => \N__44505\,
            I => \N__44404\
        );

    \I__9935\ : LocalMux
    port map (
            O => \N__44502\,
            I => \N__44401\
        );

    \I__9934\ : LocalMux
    port map (
            O => \N__44499\,
            I => \N__44397\
        );

    \I__9933\ : LocalMux
    port map (
            O => \N__44496\,
            I => \N__44394\
        );

    \I__9932\ : InMux
    port map (
            O => \N__44495\,
            I => \N__44391\
        );

    \I__9931\ : LocalMux
    port map (
            O => \N__44492\,
            I => \N__44386\
        );

    \I__9930\ : LocalMux
    port map (
            O => \N__44481\,
            I => \N__44386\
        );

    \I__9929\ : LocalMux
    port map (
            O => \N__44478\,
            I => \N__44381\
        );

    \I__9928\ : Span4Mux_h
    port map (
            O => \N__44475\,
            I => \N__44381\
        );

    \I__9927\ : CascadeMux
    port map (
            O => \N__44474\,
            I => \N__44377\
        );

    \I__9926\ : LocalMux
    port map (
            O => \N__44461\,
            I => \N__44371\
        );

    \I__9925\ : LocalMux
    port map (
            O => \N__44458\,
            I => \N__44368\
        );

    \I__9924\ : Span4Mux_v
    port map (
            O => \N__44453\,
            I => \N__44365\
        );

    \I__9923\ : Span4Mux_v
    port map (
            O => \N__44450\,
            I => \N__44358\
        );

    \I__9922\ : LocalMux
    port map (
            O => \N__44447\,
            I => \N__44358\
        );

    \I__9921\ : Span4Mux_h
    port map (
            O => \N__44444\,
            I => \N__44358\
        );

    \I__9920\ : LocalMux
    port map (
            O => \N__44427\,
            I => \N__44353\
        );

    \I__9919\ : LocalMux
    port map (
            O => \N__44420\,
            I => \N__44353\
        );

    \I__9918\ : LocalMux
    port map (
            O => \N__44417\,
            I => \N__44342\
        );

    \I__9917\ : LocalMux
    port map (
            O => \N__44414\,
            I => \N__44342\
        );

    \I__9916\ : LocalMux
    port map (
            O => \N__44407\,
            I => \N__44342\
        );

    \I__9915\ : Span4Mux_h
    port map (
            O => \N__44404\,
            I => \N__44342\
        );

    \I__9914\ : Span4Mux_h
    port map (
            O => \N__44401\,
            I => \N__44342\
        );

    \I__9913\ : InMux
    port map (
            O => \N__44400\,
            I => \N__44339\
        );

    \I__9912\ : Span4Mux_h
    port map (
            O => \N__44397\,
            I => \N__44336\
        );

    \I__9911\ : Span4Mux_h
    port map (
            O => \N__44394\,
            I => \N__44333\
        );

    \I__9910\ : LocalMux
    port map (
            O => \N__44391\,
            I => \N__44330\
        );

    \I__9909\ : Span4Mux_h
    port map (
            O => \N__44386\,
            I => \N__44325\
        );

    \I__9908\ : Span4Mux_h
    port map (
            O => \N__44381\,
            I => \N__44325\
        );

    \I__9907\ : InMux
    port map (
            O => \N__44380\,
            I => \N__44314\
        );

    \I__9906\ : InMux
    port map (
            O => \N__44377\,
            I => \N__44314\
        );

    \I__9905\ : InMux
    port map (
            O => \N__44376\,
            I => \N__44314\
        );

    \I__9904\ : InMux
    port map (
            O => \N__44375\,
            I => \N__44314\
        );

    \I__9903\ : InMux
    port map (
            O => \N__44374\,
            I => \N__44314\
        );

    \I__9902\ : Span4Mux_h
    port map (
            O => \N__44371\,
            I => \N__44305\
        );

    \I__9901\ : Span4Mux_h
    port map (
            O => \N__44368\,
            I => \N__44305\
        );

    \I__9900\ : Span4Mux_h
    port map (
            O => \N__44365\,
            I => \N__44305\
        );

    \I__9899\ : Span4Mux_v
    port map (
            O => \N__44358\,
            I => \N__44305\
        );

    \I__9898\ : Span4Mux_h
    port map (
            O => \N__44353\,
            I => \N__44300\
        );

    \I__9897\ : Span4Mux_v
    port map (
            O => \N__44342\,
            I => \N__44300\
        );

    \I__9896\ : LocalMux
    port map (
            O => \N__44339\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__9895\ : Odrv4
    port map (
            O => \N__44336\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__9894\ : Odrv4
    port map (
            O => \N__44333\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__9893\ : Odrv12
    port map (
            O => \N__44330\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__9892\ : Odrv4
    port map (
            O => \N__44325\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__9891\ : LocalMux
    port map (
            O => \N__44314\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__9890\ : Odrv4
    port map (
            O => \N__44305\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__9889\ : Odrv4
    port map (
            O => \N__44300\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__9888\ : InMux
    port map (
            O => \N__44283\,
            I => \N__44279\
        );

    \I__9887\ : InMux
    port map (
            O => \N__44282\,
            I => \N__44276\
        );

    \I__9886\ : LocalMux
    port map (
            O => \N__44279\,
            I => \N__44273\
        );

    \I__9885\ : LocalMux
    port map (
            O => \N__44276\,
            I => \N__44270\
        );

    \I__9884\ : Span4Mux_h
    port map (
            O => \N__44273\,
            I => \N__44266\
        );

    \I__9883\ : Span4Mux_h
    port map (
            O => \N__44270\,
            I => \N__44263\
        );

    \I__9882\ : InMux
    port map (
            O => \N__44269\,
            I => \N__44260\
        );

    \I__9881\ : Span4Mux_h
    port map (
            O => \N__44266\,
            I => \N__44257\
        );

    \I__9880\ : Span4Mux_h
    port map (
            O => \N__44263\,
            I => \N__44254\
        );

    \I__9879\ : LocalMux
    port map (
            O => \N__44260\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\
        );

    \I__9878\ : Odrv4
    port map (
            O => \N__44257\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\
        );

    \I__9877\ : Odrv4
    port map (
            O => \N__44254\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\
        );

    \I__9876\ : InMux
    port map (
            O => \N__44247\,
            I => \N__44244\
        );

    \I__9875\ : LocalMux
    port map (
            O => \N__44244\,
            I => \N__44240\
        );

    \I__9874\ : CascadeMux
    port map (
            O => \N__44243\,
            I => \N__44237\
        );

    \I__9873\ : Span4Mux_v
    port map (
            O => \N__44240\,
            I => \N__44233\
        );

    \I__9872\ : InMux
    port map (
            O => \N__44237\,
            I => \N__44230\
        );

    \I__9871\ : InMux
    port map (
            O => \N__44236\,
            I => \N__44227\
        );

    \I__9870\ : Odrv4
    port map (
            O => \N__44233\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__9869\ : LocalMux
    port map (
            O => \N__44230\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__9868\ : LocalMux
    port map (
            O => \N__44227\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__9867\ : CascadeMux
    port map (
            O => \N__44220\,
            I => \N__44217\
        );

    \I__9866\ : InMux
    port map (
            O => \N__44217\,
            I => \N__44213\
        );

    \I__9865\ : InMux
    port map (
            O => \N__44216\,
            I => \N__44209\
        );

    \I__9864\ : LocalMux
    port map (
            O => \N__44213\,
            I => \N__44206\
        );

    \I__9863\ : InMux
    port map (
            O => \N__44212\,
            I => \N__44203\
        );

    \I__9862\ : LocalMux
    port map (
            O => \N__44209\,
            I => \N__44200\
        );

    \I__9861\ : Span4Mux_v
    port map (
            O => \N__44206\,
            I => \N__44194\
        );

    \I__9860\ : LocalMux
    port map (
            O => \N__44203\,
            I => \N__44194\
        );

    \I__9859\ : Span4Mux_v
    port map (
            O => \N__44200\,
            I => \N__44191\
        );

    \I__9858\ : InMux
    port map (
            O => \N__44199\,
            I => \N__44188\
        );

    \I__9857\ : Sp12to4
    port map (
            O => \N__44194\,
            I => \N__44181\
        );

    \I__9856\ : Sp12to4
    port map (
            O => \N__44191\,
            I => \N__44181\
        );

    \I__9855\ : LocalMux
    port map (
            O => \N__44188\,
            I => \N__44181\
        );

    \I__9854\ : Odrv12
    port map (
            O => \N__44181\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__9853\ : CascadeMux
    port map (
            O => \N__44178\,
            I => \N__44175\
        );

    \I__9852\ : InMux
    port map (
            O => \N__44175\,
            I => \N__44172\
        );

    \I__9851\ : LocalMux
    port map (
            O => \N__44172\,
            I => \N__44169\
        );

    \I__9850\ : Span4Mux_v
    port map (
            O => \N__44169\,
            I => \N__44166\
        );

    \I__9849\ : Odrv4
    port map (
            O => \N__44166\,
            I => \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\
        );

    \I__9848\ : InMux
    port map (
            O => \N__44163\,
            I => \N__44160\
        );

    \I__9847\ : LocalMux
    port map (
            O => \N__44160\,
            I => \N__44156\
        );

    \I__9846\ : InMux
    port map (
            O => \N__44159\,
            I => \N__44152\
        );

    \I__9845\ : Span4Mux_v
    port map (
            O => \N__44156\,
            I => \N__44149\
        );

    \I__9844\ : InMux
    port map (
            O => \N__44155\,
            I => \N__44146\
        );

    \I__9843\ : LocalMux
    port map (
            O => \N__44152\,
            I => \N__44143\
        );

    \I__9842\ : Odrv4
    port map (
            O => \N__44149\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__9841\ : LocalMux
    port map (
            O => \N__44146\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__9840\ : Odrv4
    port map (
            O => \N__44143\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__9839\ : CEMux
    port map (
            O => \N__44136\,
            I => \N__44109\
        );

    \I__9838\ : CEMux
    port map (
            O => \N__44135\,
            I => \N__44109\
        );

    \I__9837\ : CEMux
    port map (
            O => \N__44134\,
            I => \N__44109\
        );

    \I__9836\ : CEMux
    port map (
            O => \N__44133\,
            I => \N__44109\
        );

    \I__9835\ : CEMux
    port map (
            O => \N__44132\,
            I => \N__44109\
        );

    \I__9834\ : CEMux
    port map (
            O => \N__44131\,
            I => \N__44109\
        );

    \I__9833\ : CEMux
    port map (
            O => \N__44130\,
            I => \N__44109\
        );

    \I__9832\ : CEMux
    port map (
            O => \N__44129\,
            I => \N__44109\
        );

    \I__9831\ : CEMux
    port map (
            O => \N__44128\,
            I => \N__44109\
        );

    \I__9830\ : GlobalMux
    port map (
            O => \N__44109\,
            I => \N__44106\
        );

    \I__9829\ : gio2CtrlBuf
    port map (
            O => \N__44106\,
            I => \current_shift_inst.timer_s1.N_166_i_g\
        );

    \I__9828\ : CascadeMux
    port map (
            O => \N__44103\,
            I => \N__44099\
        );

    \I__9827\ : InMux
    port map (
            O => \N__44102\,
            I => \N__44094\
        );

    \I__9826\ : InMux
    port map (
            O => \N__44099\,
            I => \N__44094\
        );

    \I__9825\ : LocalMux
    port map (
            O => \N__44094\,
            I => \N__44090\
        );

    \I__9824\ : InMux
    port map (
            O => \N__44093\,
            I => \N__44087\
        );

    \I__9823\ : Span4Mux_h
    port map (
            O => \N__44090\,
            I => \N__44081\
        );

    \I__9822\ : LocalMux
    port map (
            O => \N__44087\,
            I => \N__44081\
        );

    \I__9821\ : InMux
    port map (
            O => \N__44086\,
            I => \N__44078\
        );

    \I__9820\ : Span4Mux_v
    port map (
            O => \N__44081\,
            I => \N__44075\
        );

    \I__9819\ : LocalMux
    port map (
            O => \N__44078\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__9818\ : Odrv4
    port map (
            O => \N__44075\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__9817\ : CascadeMux
    port map (
            O => \N__44070\,
            I => \N__44067\
        );

    \I__9816\ : InMux
    port map (
            O => \N__44067\,
            I => \N__44064\
        );

    \I__9815\ : LocalMux
    port map (
            O => \N__44064\,
            I => \N__44061\
        );

    \I__9814\ : Span4Mux_h
    port map (
            O => \N__44061\,
            I => \N__44058\
        );

    \I__9813\ : Odrv4
    port map (
            O => \N__44058\,
            I => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\
        );

    \I__9812\ : InMux
    port map (
            O => \N__44055\,
            I => \N__44042\
        );

    \I__9811\ : InMux
    port map (
            O => \N__44054\,
            I => \N__44033\
        );

    \I__9810\ : InMux
    port map (
            O => \N__44053\,
            I => \N__44028\
        );

    \I__9809\ : InMux
    port map (
            O => \N__44052\,
            I => \N__44028\
        );

    \I__9808\ : InMux
    port map (
            O => \N__44051\,
            I => \N__44025\
        );

    \I__9807\ : InMux
    port map (
            O => \N__44050\,
            I => \N__44004\
        );

    \I__9806\ : InMux
    port map (
            O => \N__44049\,
            I => \N__44004\
        );

    \I__9805\ : InMux
    port map (
            O => \N__44048\,
            I => \N__44004\
        );

    \I__9804\ : InMux
    port map (
            O => \N__44047\,
            I => \N__44004\
        );

    \I__9803\ : InMux
    port map (
            O => \N__44046\,
            I => \N__44004\
        );

    \I__9802\ : InMux
    port map (
            O => \N__44045\,
            I => \N__44004\
        );

    \I__9801\ : LocalMux
    port map (
            O => \N__44042\,
            I => \N__44001\
        );

    \I__9800\ : InMux
    port map (
            O => \N__44041\,
            I => \N__43992\
        );

    \I__9799\ : InMux
    port map (
            O => \N__44040\,
            I => \N__43992\
        );

    \I__9798\ : InMux
    port map (
            O => \N__44039\,
            I => \N__43992\
        );

    \I__9797\ : InMux
    port map (
            O => \N__44038\,
            I => \N__43992\
        );

    \I__9796\ : InMux
    port map (
            O => \N__44037\,
            I => \N__43987\
        );

    \I__9795\ : InMux
    port map (
            O => \N__44036\,
            I => \N__43987\
        );

    \I__9794\ : LocalMux
    port map (
            O => \N__44033\,
            I => \N__43984\
        );

    \I__9793\ : LocalMux
    port map (
            O => \N__44028\,
            I => \N__43981\
        );

    \I__9792\ : LocalMux
    port map (
            O => \N__44025\,
            I => \N__43978\
        );

    \I__9791\ : InMux
    port map (
            O => \N__44024\,
            I => \N__43975\
        );

    \I__9790\ : InMux
    port map (
            O => \N__44023\,
            I => \N__43960\
        );

    \I__9789\ : InMux
    port map (
            O => \N__44022\,
            I => \N__43960\
        );

    \I__9788\ : InMux
    port map (
            O => \N__44021\,
            I => \N__43960\
        );

    \I__9787\ : InMux
    port map (
            O => \N__44020\,
            I => \N__43960\
        );

    \I__9786\ : InMux
    port map (
            O => \N__44019\,
            I => \N__43960\
        );

    \I__9785\ : InMux
    port map (
            O => \N__44018\,
            I => \N__43960\
        );

    \I__9784\ : InMux
    port map (
            O => \N__44017\,
            I => \N__43960\
        );

    \I__9783\ : LocalMux
    port map (
            O => \N__44004\,
            I => \N__43955\
        );

    \I__9782\ : Span4Mux_h
    port map (
            O => \N__44001\,
            I => \N__43955\
        );

    \I__9781\ : LocalMux
    port map (
            O => \N__43992\,
            I => \N__43952\
        );

    \I__9780\ : LocalMux
    port map (
            O => \N__43987\,
            I => \N__43945\
        );

    \I__9779\ : Span4Mux_v
    port map (
            O => \N__43984\,
            I => \N__43945\
        );

    \I__9778\ : Span4Mux_v
    port map (
            O => \N__43981\,
            I => \N__43945\
        );

    \I__9777\ : Odrv4
    port map (
            O => \N__43978\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__9776\ : LocalMux
    port map (
            O => \N__43975\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__9775\ : LocalMux
    port map (
            O => \N__43960\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__9774\ : Odrv4
    port map (
            O => \N__43955\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__9773\ : Odrv12
    port map (
            O => \N__43952\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__9772\ : Odrv4
    port map (
            O => \N__43945\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__9771\ : CascadeMux
    port map (
            O => \N__43932\,
            I => \N__43928\
        );

    \I__9770\ : InMux
    port map (
            O => \N__43931\,
            I => \N__43920\
        );

    \I__9769\ : InMux
    port map (
            O => \N__43928\,
            I => \N__43920\
        );

    \I__9768\ : InMux
    port map (
            O => \N__43927\,
            I => \N__43920\
        );

    \I__9767\ : LocalMux
    port map (
            O => \N__43920\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__9766\ : InMux
    port map (
            O => \N__43917\,
            I => \N__43907\
        );

    \I__9765\ : InMux
    port map (
            O => \N__43916\,
            I => \N__43907\
        );

    \I__9764\ : InMux
    port map (
            O => \N__43915\,
            I => \N__43907\
        );

    \I__9763\ : InMux
    port map (
            O => \N__43914\,
            I => \N__43904\
        );

    \I__9762\ : LocalMux
    port map (
            O => \N__43907\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__9761\ : LocalMux
    port map (
            O => \N__43904\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__9760\ : CascadeMux
    port map (
            O => \N__43899\,
            I => \N__43896\
        );

    \I__9759\ : InMux
    port map (
            O => \N__43896\,
            I => \N__43893\
        );

    \I__9758\ : LocalMux
    port map (
            O => \N__43893\,
            I => \N__43890\
        );

    \I__9757\ : Span4Mux_h
    port map (
            O => \N__43890\,
            I => \N__43887\
        );

    \I__9756\ : Odrv4
    port map (
            O => \N__43887\,
            I => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\
        );

    \I__9755\ : CascadeMux
    port map (
            O => \N__43884\,
            I => \N__43881\
        );

    \I__9754\ : InMux
    port map (
            O => \N__43881\,
            I => \N__43878\
        );

    \I__9753\ : LocalMux
    port map (
            O => \N__43878\,
            I => \N__43875\
        );

    \I__9752\ : Span4Mux_h
    port map (
            O => \N__43875\,
            I => \N__43872\
        );

    \I__9751\ : Odrv4
    port map (
            O => \N__43872\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\
        );

    \I__9750\ : CascadeMux
    port map (
            O => \N__43869\,
            I => \N__43866\
        );

    \I__9749\ : InMux
    port map (
            O => \N__43866\,
            I => \N__43863\
        );

    \I__9748\ : LocalMux
    port map (
            O => \N__43863\,
            I => \N__43860\
        );

    \I__9747\ : Span12Mux_h
    port map (
            O => \N__43860\,
            I => \N__43857\
        );

    \I__9746\ : Odrv12
    port map (
            O => \N__43857\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\
        );

    \I__9745\ : CascadeMux
    port map (
            O => \N__43854\,
            I => \N__43851\
        );

    \I__9744\ : InMux
    port map (
            O => \N__43851\,
            I => \N__43847\
        );

    \I__9743\ : InMux
    port map (
            O => \N__43850\,
            I => \N__43844\
        );

    \I__9742\ : LocalMux
    port map (
            O => \N__43847\,
            I => \N__43836\
        );

    \I__9741\ : LocalMux
    port map (
            O => \N__43844\,
            I => \N__43836\
        );

    \I__9740\ : InMux
    port map (
            O => \N__43843\,
            I => \N__43831\
        );

    \I__9739\ : InMux
    port map (
            O => \N__43842\,
            I => \N__43831\
        );

    \I__9738\ : InMux
    port map (
            O => \N__43841\,
            I => \N__43828\
        );

    \I__9737\ : Span4Mux_h
    port map (
            O => \N__43836\,
            I => \N__43823\
        );

    \I__9736\ : LocalMux
    port map (
            O => \N__43831\,
            I => \N__43823\
        );

    \I__9735\ : LocalMux
    port map (
            O => \N__43828\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__9734\ : Odrv4
    port map (
            O => \N__43823\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__9733\ : InMux
    port map (
            O => \N__43818\,
            I => \N__43813\
        );

    \I__9732\ : InMux
    port map (
            O => \N__43817\,
            I => \N__43808\
        );

    \I__9731\ : InMux
    port map (
            O => \N__43816\,
            I => \N__43808\
        );

    \I__9730\ : LocalMux
    port map (
            O => \N__43813\,
            I => \N__43803\
        );

    \I__9729\ : LocalMux
    port map (
            O => \N__43808\,
            I => \N__43803\
        );

    \I__9728\ : Odrv4
    port map (
            O => \N__43803\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__9727\ : CascadeMux
    port map (
            O => \N__43800\,
            I => \N__43797\
        );

    \I__9726\ : InMux
    port map (
            O => \N__43797\,
            I => \N__43794\
        );

    \I__9725\ : LocalMux
    port map (
            O => \N__43794\,
            I => \N__43791\
        );

    \I__9724\ : Span4Mux_h
    port map (
            O => \N__43791\,
            I => \N__43788\
        );

    \I__9723\ : Span4Mux_v
    port map (
            O => \N__43788\,
            I => \N__43785\
        );

    \I__9722\ : Odrv4
    port map (
            O => \N__43785\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\
        );

    \I__9721\ : CascadeMux
    port map (
            O => \N__43782\,
            I => \N__43779\
        );

    \I__9720\ : InMux
    port map (
            O => \N__43779\,
            I => \N__43776\
        );

    \I__9719\ : LocalMux
    port map (
            O => \N__43776\,
            I => \N__43770\
        );

    \I__9718\ : InMux
    port map (
            O => \N__43775\,
            I => \N__43765\
        );

    \I__9717\ : InMux
    port map (
            O => \N__43774\,
            I => \N__43765\
        );

    \I__9716\ : InMux
    port map (
            O => \N__43773\,
            I => \N__43762\
        );

    \I__9715\ : Span4Mux_v
    port map (
            O => \N__43770\,
            I => \N__43759\
        );

    \I__9714\ : LocalMux
    port map (
            O => \N__43765\,
            I => \N__43756\
        );

    \I__9713\ : LocalMux
    port map (
            O => \N__43762\,
            I => \N__43753\
        );

    \I__9712\ : Span4Mux_h
    port map (
            O => \N__43759\,
            I => \N__43750\
        );

    \I__9711\ : Span4Mux_h
    port map (
            O => \N__43756\,
            I => \N__43747\
        );

    \I__9710\ : Odrv4
    port map (
            O => \N__43753\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__9709\ : Odrv4
    port map (
            O => \N__43750\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__9708\ : Odrv4
    port map (
            O => \N__43747\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__9707\ : CascadeMux
    port map (
            O => \N__43740\,
            I => \N__43737\
        );

    \I__9706\ : InMux
    port map (
            O => \N__43737\,
            I => \N__43733\
        );

    \I__9705\ : InMux
    port map (
            O => \N__43736\,
            I => \N__43729\
        );

    \I__9704\ : LocalMux
    port map (
            O => \N__43733\,
            I => \N__43726\
        );

    \I__9703\ : InMux
    port map (
            O => \N__43732\,
            I => \N__43723\
        );

    \I__9702\ : LocalMux
    port map (
            O => \N__43729\,
            I => \N__43718\
        );

    \I__9701\ : Span4Mux_v
    port map (
            O => \N__43726\,
            I => \N__43718\
        );

    \I__9700\ : LocalMux
    port map (
            O => \N__43723\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__9699\ : Odrv4
    port map (
            O => \N__43718\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__9698\ : InMux
    port map (
            O => \N__43713\,
            I => \N__43710\
        );

    \I__9697\ : LocalMux
    port map (
            O => \N__43710\,
            I => \N__43707\
        );

    \I__9696\ : Span4Mux_v
    port map (
            O => \N__43707\,
            I => \N__43704\
        );

    \I__9695\ : Odrv4
    port map (
            O => \N__43704\,
            I => \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\
        );

    \I__9694\ : CascadeMux
    port map (
            O => \N__43701\,
            I => \N__43697\
        );

    \I__9693\ : CascadeMux
    port map (
            O => \N__43700\,
            I => \N__43694\
        );

    \I__9692\ : InMux
    port map (
            O => \N__43697\,
            I => \N__43690\
        );

    \I__9691\ : InMux
    port map (
            O => \N__43694\,
            I => \N__43687\
        );

    \I__9690\ : InMux
    port map (
            O => \N__43693\,
            I => \N__43684\
        );

    \I__9689\ : LocalMux
    port map (
            O => \N__43690\,
            I => \N__43680\
        );

    \I__9688\ : LocalMux
    port map (
            O => \N__43687\,
            I => \N__43677\
        );

    \I__9687\ : LocalMux
    port map (
            O => \N__43684\,
            I => \N__43674\
        );

    \I__9686\ : InMux
    port map (
            O => \N__43683\,
            I => \N__43671\
        );

    \I__9685\ : Span4Mux_h
    port map (
            O => \N__43680\,
            I => \N__43668\
        );

    \I__9684\ : Span4Mux_v
    port map (
            O => \N__43677\,
            I => \N__43663\
        );

    \I__9683\ : Span4Mux_h
    port map (
            O => \N__43674\,
            I => \N__43663\
        );

    \I__9682\ : LocalMux
    port map (
            O => \N__43671\,
            I => \N__43660\
        );

    \I__9681\ : Span4Mux_h
    port map (
            O => \N__43668\,
            I => \N__43657\
        );

    \I__9680\ : Span4Mux_h
    port map (
            O => \N__43663\,
            I => \N__43654\
        );

    \I__9679\ : Odrv12
    port map (
            O => \N__43660\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__9678\ : Odrv4
    port map (
            O => \N__43657\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__9677\ : Odrv4
    port map (
            O => \N__43654\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__9676\ : InMux
    port map (
            O => \N__43647\,
            I => \N__43643\
        );

    \I__9675\ : InMux
    port map (
            O => \N__43646\,
            I => \N__43639\
        );

    \I__9674\ : LocalMux
    port map (
            O => \N__43643\,
            I => \N__43636\
        );

    \I__9673\ : InMux
    port map (
            O => \N__43642\,
            I => \N__43633\
        );

    \I__9672\ : LocalMux
    port map (
            O => \N__43639\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__9671\ : Odrv4
    port map (
            O => \N__43636\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__9670\ : LocalMux
    port map (
            O => \N__43633\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__9669\ : CascadeMux
    port map (
            O => \N__43626\,
            I => \N__43623\
        );

    \I__9668\ : InMux
    port map (
            O => \N__43623\,
            I => \N__43620\
        );

    \I__9667\ : LocalMux
    port map (
            O => \N__43620\,
            I => \N__43617\
        );

    \I__9666\ : Span4Mux_v
    port map (
            O => \N__43617\,
            I => \N__43614\
        );

    \I__9665\ : Odrv4
    port map (
            O => \N__43614\,
            I => \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\
        );

    \I__9664\ : InMux
    port map (
            O => \N__43611\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__9663\ : CascadeMux
    port map (
            O => \N__43608\,
            I => \N__43604\
        );

    \I__9662\ : InMux
    port map (
            O => \N__43607\,
            I => \N__43600\
        );

    \I__9661\ : InMux
    port map (
            O => \N__43604\,
            I => \N__43597\
        );

    \I__9660\ : InMux
    port map (
            O => \N__43603\,
            I => \N__43594\
        );

    \I__9659\ : LocalMux
    port map (
            O => \N__43600\,
            I => \N__43591\
        );

    \I__9658\ : LocalMux
    port map (
            O => \N__43597\,
            I => \N__43588\
        );

    \I__9657\ : LocalMux
    port map (
            O => \N__43594\,
            I => \N__43585\
        );

    \I__9656\ : Span4Mux_v
    port map (
            O => \N__43591\,
            I => \N__43580\
        );

    \I__9655\ : Span4Mux_h
    port map (
            O => \N__43588\,
            I => \N__43580\
        );

    \I__9654\ : Span12Mux_h
    port map (
            O => \N__43585\,
            I => \N__43576\
        );

    \I__9653\ : Span4Mux_h
    port map (
            O => \N__43580\,
            I => \N__43573\
        );

    \I__9652\ : InMux
    port map (
            O => \N__43579\,
            I => \N__43570\
        );

    \I__9651\ : Odrv12
    port map (
            O => \N__43576\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__9650\ : Odrv4
    port map (
            O => \N__43573\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__9649\ : LocalMux
    port map (
            O => \N__43570\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__9648\ : CascadeMux
    port map (
            O => \N__43563\,
            I => \N__43560\
        );

    \I__9647\ : InMux
    port map (
            O => \N__43560\,
            I => \N__43557\
        );

    \I__9646\ : LocalMux
    port map (
            O => \N__43557\,
            I => \N__43554\
        );

    \I__9645\ : Span4Mux_v
    port map (
            O => \N__43554\,
            I => \N__43549\
        );

    \I__9644\ : InMux
    port map (
            O => \N__43553\,
            I => \N__43546\
        );

    \I__9643\ : InMux
    port map (
            O => \N__43552\,
            I => \N__43543\
        );

    \I__9642\ : Odrv4
    port map (
            O => \N__43549\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__9641\ : LocalMux
    port map (
            O => \N__43546\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__9640\ : LocalMux
    port map (
            O => \N__43543\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__9639\ : CascadeMux
    port map (
            O => \N__43536\,
            I => \N__43533\
        );

    \I__9638\ : InMux
    port map (
            O => \N__43533\,
            I => \N__43530\
        );

    \I__9637\ : LocalMux
    port map (
            O => \N__43530\,
            I => \N__43527\
        );

    \I__9636\ : Sp12to4
    port map (
            O => \N__43527\,
            I => \N__43524\
        );

    \I__9635\ : Odrv12
    port map (
            O => \N__43524\,
            I => \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\
        );

    \I__9634\ : CascadeMux
    port map (
            O => \N__43521\,
            I => \N__43518\
        );

    \I__9633\ : InMux
    port map (
            O => \N__43518\,
            I => \N__43515\
        );

    \I__9632\ : LocalMux
    port map (
            O => \N__43515\,
            I => \current_shift_inst.un4_control_input_1_axb_12\
        );

    \I__9631\ : InMux
    port map (
            O => \N__43512\,
            I => \N__43509\
        );

    \I__9630\ : LocalMux
    port map (
            O => \N__43509\,
            I => \N__43506\
        );

    \I__9629\ : Odrv4
    port map (
            O => \N__43506\,
            I => \current_shift_inst.un4_control_input_1_axb_1\
        );

    \I__9628\ : CascadeMux
    port map (
            O => \N__43503\,
            I => \N__43499\
        );

    \I__9627\ : CascadeMux
    port map (
            O => \N__43502\,
            I => \N__43496\
        );

    \I__9626\ : InMux
    port map (
            O => \N__43499\,
            I => \N__43493\
        );

    \I__9625\ : InMux
    port map (
            O => \N__43496\,
            I => \N__43490\
        );

    \I__9624\ : LocalMux
    port map (
            O => \N__43493\,
            I => \N__43485\
        );

    \I__9623\ : LocalMux
    port map (
            O => \N__43490\,
            I => \N__43482\
        );

    \I__9622\ : InMux
    port map (
            O => \N__43489\,
            I => \N__43477\
        );

    \I__9621\ : InMux
    port map (
            O => \N__43488\,
            I => \N__43477\
        );

    \I__9620\ : Span4Mux_v
    port map (
            O => \N__43485\,
            I => \N__43474\
        );

    \I__9619\ : Span12Mux_s7_v
    port map (
            O => \N__43482\,
            I => \N__43469\
        );

    \I__9618\ : LocalMux
    port map (
            O => \N__43477\,
            I => \N__43469\
        );

    \I__9617\ : Odrv4
    port map (
            O => \N__43474\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__9616\ : Odrv12
    port map (
            O => \N__43469\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__9615\ : InMux
    port map (
            O => \N__43464\,
            I => \N__43461\
        );

    \I__9614\ : LocalMux
    port map (
            O => \N__43461\,
            I => \N__43458\
        );

    \I__9613\ : Span4Mux_v
    port map (
            O => \N__43458\,
            I => \N__43453\
        );

    \I__9612\ : InMux
    port map (
            O => \N__43457\,
            I => \N__43450\
        );

    \I__9611\ : InMux
    port map (
            O => \N__43456\,
            I => \N__43447\
        );

    \I__9610\ : Odrv4
    port map (
            O => \N__43453\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__9609\ : LocalMux
    port map (
            O => \N__43450\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__9608\ : LocalMux
    port map (
            O => \N__43447\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__9607\ : InMux
    port map (
            O => \N__43440\,
            I => \N__43437\
        );

    \I__9606\ : LocalMux
    port map (
            O => \N__43437\,
            I => \N__43434\
        );

    \I__9605\ : Span4Mux_v
    port map (
            O => \N__43434\,
            I => \N__43431\
        );

    \I__9604\ : Odrv4
    port map (
            O => \N__43431\,
            I => \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\
        );

    \I__9603\ : CascadeMux
    port map (
            O => \N__43428\,
            I => \N__43425\
        );

    \I__9602\ : InMux
    port map (
            O => \N__43425\,
            I => \N__43422\
        );

    \I__9601\ : LocalMux
    port map (
            O => \N__43422\,
            I => \N__43418\
        );

    \I__9600\ : CascadeMux
    port map (
            O => \N__43421\,
            I => \N__43415\
        );

    \I__9599\ : Span4Mux_v
    port map (
            O => \N__43418\,
            I => \N__43410\
        );

    \I__9598\ : InMux
    port map (
            O => \N__43415\,
            I => \N__43407\
        );

    \I__9597\ : InMux
    port map (
            O => \N__43414\,
            I => \N__43402\
        );

    \I__9596\ : InMux
    port map (
            O => \N__43413\,
            I => \N__43402\
        );

    \I__9595\ : Span4Mux_h
    port map (
            O => \N__43410\,
            I => \N__43399\
        );

    \I__9594\ : LocalMux
    port map (
            O => \N__43407\,
            I => \N__43396\
        );

    \I__9593\ : LocalMux
    port map (
            O => \N__43402\,
            I => \N__43393\
        );

    \I__9592\ : Odrv4
    port map (
            O => \N__43399\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__9591\ : Odrv12
    port map (
            O => \N__43396\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__9590\ : Odrv4
    port map (
            O => \N__43393\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__9589\ : InMux
    port map (
            O => \N__43386\,
            I => \N__43382\
        );

    \I__9588\ : InMux
    port map (
            O => \N__43385\,
            I => \N__43379\
        );

    \I__9587\ : LocalMux
    port map (
            O => \N__43382\,
            I => \N__43375\
        );

    \I__9586\ : LocalMux
    port map (
            O => \N__43379\,
            I => \N__43372\
        );

    \I__9585\ : InMux
    port map (
            O => \N__43378\,
            I => \N__43369\
        );

    \I__9584\ : Span4Mux_v
    port map (
            O => \N__43375\,
            I => \N__43364\
        );

    \I__9583\ : Span4Mux_h
    port map (
            O => \N__43372\,
            I => \N__43364\
        );

    \I__9582\ : LocalMux
    port map (
            O => \N__43369\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__9581\ : Odrv4
    port map (
            O => \N__43364\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__9580\ : CascadeMux
    port map (
            O => \N__43359\,
            I => \N__43356\
        );

    \I__9579\ : InMux
    port map (
            O => \N__43356\,
            I => \N__43353\
        );

    \I__9578\ : LocalMux
    port map (
            O => \N__43353\,
            I => \N__43350\
        );

    \I__9577\ : Span4Mux_v
    port map (
            O => \N__43350\,
            I => \N__43347\
        );

    \I__9576\ : Odrv4
    port map (
            O => \N__43347\,
            I => \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\
        );

    \I__9575\ : InMux
    port map (
            O => \N__43344\,
            I => \N__43341\
        );

    \I__9574\ : LocalMux
    port map (
            O => \N__43341\,
            I => \current_shift_inst.un4_control_input_1_axb_14\
        );

    \I__9573\ : CascadeMux
    port map (
            O => \N__43338\,
            I => \N__43335\
        );

    \I__9572\ : InMux
    port map (
            O => \N__43335\,
            I => \N__43331\
        );

    \I__9571\ : InMux
    port map (
            O => \N__43334\,
            I => \N__43328\
        );

    \I__9570\ : LocalMux
    port map (
            O => \N__43331\,
            I => \N__43322\
        );

    \I__9569\ : LocalMux
    port map (
            O => \N__43328\,
            I => \N__43322\
        );

    \I__9568\ : InMux
    port map (
            O => \N__43327\,
            I => \N__43319\
        );

    \I__9567\ : Odrv4
    port map (
            O => \N__43322\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__9566\ : LocalMux
    port map (
            O => \N__43319\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__9565\ : InMux
    port map (
            O => \N__43314\,
            I => \N__43309\
        );

    \I__9564\ : InMux
    port map (
            O => \N__43313\,
            I => \N__43306\
        );

    \I__9563\ : CascadeMux
    port map (
            O => \N__43312\,
            I => \N__43303\
        );

    \I__9562\ : LocalMux
    port map (
            O => \N__43309\,
            I => \N__43299\
        );

    \I__9561\ : LocalMux
    port map (
            O => \N__43306\,
            I => \N__43296\
        );

    \I__9560\ : InMux
    port map (
            O => \N__43303\,
            I => \N__43291\
        );

    \I__9559\ : InMux
    port map (
            O => \N__43302\,
            I => \N__43291\
        );

    \I__9558\ : Span4Mux_h
    port map (
            O => \N__43299\,
            I => \N__43284\
        );

    \I__9557\ : Span4Mux_v
    port map (
            O => \N__43296\,
            I => \N__43284\
        );

    \I__9556\ : LocalMux
    port map (
            O => \N__43291\,
            I => \N__43284\
        );

    \I__9555\ : Odrv4
    port map (
            O => \N__43284\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__9554\ : CascadeMux
    port map (
            O => \N__43281\,
            I => \N__43278\
        );

    \I__9553\ : InMux
    port map (
            O => \N__43278\,
            I => \N__43275\
        );

    \I__9552\ : LocalMux
    port map (
            O => \N__43275\,
            I => \N__43272\
        );

    \I__9551\ : Sp12to4
    port map (
            O => \N__43272\,
            I => \N__43269\
        );

    \I__9550\ : Odrv12
    port map (
            O => \N__43269\,
            I => \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\
        );

    \I__9549\ : CascadeMux
    port map (
            O => \N__43266\,
            I => \N__43263\
        );

    \I__9548\ : InMux
    port map (
            O => \N__43263\,
            I => \N__43260\
        );

    \I__9547\ : LocalMux
    port map (
            O => \N__43260\,
            I => \N__43257\
        );

    \I__9546\ : Span4Mux_h
    port map (
            O => \N__43257\,
            I => \N__43254\
        );

    \I__9545\ : Span4Mux_v
    port map (
            O => \N__43254\,
            I => \N__43251\
        );

    \I__9544\ : Odrv4
    port map (
            O => \N__43251\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2\
        );

    \I__9543\ : CascadeMux
    port map (
            O => \N__43248\,
            I => \N__43245\
        );

    \I__9542\ : InMux
    port map (
            O => \N__43245\,
            I => \N__43242\
        );

    \I__9541\ : LocalMux
    port map (
            O => \N__43242\,
            I => \N__43238\
        );

    \I__9540\ : InMux
    port map (
            O => \N__43241\,
            I => \N__43235\
        );

    \I__9539\ : Odrv12
    port map (
            O => \N__43238\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__9538\ : LocalMux
    port map (
            O => \N__43235\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__9537\ : InMux
    port map (
            O => \N__43230\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__9536\ : CascadeMux
    port map (
            O => \N__43227\,
            I => \N__43224\
        );

    \I__9535\ : InMux
    port map (
            O => \N__43224\,
            I => \N__43221\
        );

    \I__9534\ : LocalMux
    port map (
            O => \N__43221\,
            I => \N__43217\
        );

    \I__9533\ : InMux
    port map (
            O => \N__43220\,
            I => \N__43214\
        );

    \I__9532\ : Span4Mux_v
    port map (
            O => \N__43217\,
            I => \N__43209\
        );

    \I__9531\ : LocalMux
    port map (
            O => \N__43214\,
            I => \N__43209\
        );

    \I__9530\ : Odrv4
    port map (
            O => \N__43209\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__9529\ : InMux
    port map (
            O => \N__43206\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__9528\ : CascadeMux
    port map (
            O => \N__43203\,
            I => \N__43200\
        );

    \I__9527\ : InMux
    port map (
            O => \N__43200\,
            I => \N__43196\
        );

    \I__9526\ : CascadeMux
    port map (
            O => \N__43199\,
            I => \N__43193\
        );

    \I__9525\ : LocalMux
    port map (
            O => \N__43196\,
            I => \N__43190\
        );

    \I__9524\ : InMux
    port map (
            O => \N__43193\,
            I => \N__43187\
        );

    \I__9523\ : Span4Mux_v
    port map (
            O => \N__43190\,
            I => \N__43182\
        );

    \I__9522\ : LocalMux
    port map (
            O => \N__43187\,
            I => \N__43182\
        );

    \I__9521\ : Odrv4
    port map (
            O => \N__43182\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__9520\ : InMux
    port map (
            O => \N__43179\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__9519\ : InMux
    port map (
            O => \N__43176\,
            I => \N__43173\
        );

    \I__9518\ : LocalMux
    port map (
            O => \N__43173\,
            I => \N__43170\
        );

    \I__9517\ : Span4Mux_v
    port map (
            O => \N__43170\,
            I => \N__43166\
        );

    \I__9516\ : InMux
    port map (
            O => \N__43169\,
            I => \N__43163\
        );

    \I__9515\ : Odrv4
    port map (
            O => \N__43166\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__9514\ : LocalMux
    port map (
            O => \N__43163\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__9513\ : InMux
    port map (
            O => \N__43158\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__9512\ : InMux
    port map (
            O => \N__43155\,
            I => \N__43152\
        );

    \I__9511\ : LocalMux
    port map (
            O => \N__43152\,
            I => \N__43148\
        );

    \I__9510\ : CascadeMux
    port map (
            O => \N__43151\,
            I => \N__43145\
        );

    \I__9509\ : Span4Mux_v
    port map (
            O => \N__43148\,
            I => \N__43142\
        );

    \I__9508\ : InMux
    port map (
            O => \N__43145\,
            I => \N__43139\
        );

    \I__9507\ : Odrv4
    port map (
            O => \N__43142\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__9506\ : LocalMux
    port map (
            O => \N__43139\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__9505\ : InMux
    port map (
            O => \N__43134\,
            I => \bfn_17_22_0_\
        );

    \I__9504\ : InMux
    port map (
            O => \N__43131\,
            I => \N__43128\
        );

    \I__9503\ : LocalMux
    port map (
            O => \N__43128\,
            I => \N__43125\
        );

    \I__9502\ : Span4Mux_v
    port map (
            O => \N__43125\,
            I => \N__43121\
        );

    \I__9501\ : InMux
    port map (
            O => \N__43124\,
            I => \N__43118\
        );

    \I__9500\ : Odrv4
    port map (
            O => \N__43121\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__9499\ : LocalMux
    port map (
            O => \N__43118\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__9498\ : InMux
    port map (
            O => \N__43113\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__9497\ : InMux
    port map (
            O => \N__43110\,
            I => \N__43106\
        );

    \I__9496\ : InMux
    port map (
            O => \N__43109\,
            I => \N__43103\
        );

    \I__9495\ : LocalMux
    port map (
            O => \N__43106\,
            I => \N__43100\
        );

    \I__9494\ : LocalMux
    port map (
            O => \N__43103\,
            I => \N__43097\
        );

    \I__9493\ : Odrv12
    port map (
            O => \N__43100\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__9492\ : Odrv4
    port map (
            O => \N__43097\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__9491\ : InMux
    port map (
            O => \N__43092\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__9490\ : InMux
    port map (
            O => \N__43089\,
            I => \N__43085\
        );

    \I__9489\ : InMux
    port map (
            O => \N__43088\,
            I => \N__43082\
        );

    \I__9488\ : LocalMux
    port map (
            O => \N__43085\,
            I => \N__43079\
        );

    \I__9487\ : LocalMux
    port map (
            O => \N__43082\,
            I => \N__43076\
        );

    \I__9486\ : Odrv12
    port map (
            O => \N__43079\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__9485\ : Odrv4
    port map (
            O => \N__43076\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__9484\ : InMux
    port map (
            O => \N__43071\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__9483\ : InMux
    port map (
            O => \N__43068\,
            I => \N__43063\
        );

    \I__9482\ : InMux
    port map (
            O => \N__43067\,
            I => \N__43057\
        );

    \I__9481\ : InMux
    port map (
            O => \N__43066\,
            I => \N__43057\
        );

    \I__9480\ : LocalMux
    port map (
            O => \N__43063\,
            I => \N__43054\
        );

    \I__9479\ : InMux
    port map (
            O => \N__43062\,
            I => \N__43051\
        );

    \I__9478\ : LocalMux
    port map (
            O => \N__43057\,
            I => \N__43048\
        );

    \I__9477\ : Odrv4
    port map (
            O => \N__43054\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\
        );

    \I__9476\ : LocalMux
    port map (
            O => \N__43051\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\
        );

    \I__9475\ : Odrv4
    port map (
            O => \N__43048\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\
        );

    \I__9474\ : InMux
    port map (
            O => \N__43041\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__9473\ : InMux
    port map (
            O => \N__43038\,
            I => \N__43034\
        );

    \I__9472\ : InMux
    port map (
            O => \N__43037\,
            I => \N__43031\
        );

    \I__9471\ : LocalMux
    port map (
            O => \N__43034\,
            I => \N__43028\
        );

    \I__9470\ : LocalMux
    port map (
            O => \N__43031\,
            I => \N__43025\
        );

    \I__9469\ : Span4Mux_v
    port map (
            O => \N__43028\,
            I => \N__43019\
        );

    \I__9468\ : Span4Mux_h
    port map (
            O => \N__43025\,
            I => \N__43019\
        );

    \I__9467\ : InMux
    port map (
            O => \N__43024\,
            I => \N__43016\
        );

    \I__9466\ : Odrv4
    port map (
            O => \N__43019\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto15\
        );

    \I__9465\ : LocalMux
    port map (
            O => \N__43016\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto15\
        );

    \I__9464\ : InMux
    port map (
            O => \N__43011\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__9463\ : InMux
    port map (
            O => \N__43008\,
            I => \N__43003\
        );

    \I__9462\ : CascadeMux
    port map (
            O => \N__43007\,
            I => \N__43000\
        );

    \I__9461\ : CascadeMux
    port map (
            O => \N__43006\,
            I => \N__42997\
        );

    \I__9460\ : LocalMux
    port map (
            O => \N__43003\,
            I => \N__42994\
        );

    \I__9459\ : InMux
    port map (
            O => \N__43000\,
            I => \N__42991\
        );

    \I__9458\ : InMux
    port map (
            O => \N__42997\,
            I => \N__42988\
        );

    \I__9457\ : Odrv4
    port map (
            O => \N__42994\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__42991\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__9455\ : LocalMux
    port map (
            O => \N__42988\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__9454\ : InMux
    port map (
            O => \N__42981\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__9453\ : InMux
    port map (
            O => \N__42978\,
            I => \N__42975\
        );

    \I__9452\ : LocalMux
    port map (
            O => \N__42975\,
            I => \N__42971\
        );

    \I__9451\ : InMux
    port map (
            O => \N__42974\,
            I => \N__42968\
        );

    \I__9450\ : Span4Mux_v
    port map (
            O => \N__42971\,
            I => \N__42964\
        );

    \I__9449\ : LocalMux
    port map (
            O => \N__42968\,
            I => \N__42961\
        );

    \I__9448\ : InMux
    port map (
            O => \N__42967\,
            I => \N__42958\
        );

    \I__9447\ : Odrv4
    port map (
            O => \N__42964\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__9446\ : Odrv4
    port map (
            O => \N__42961\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__9445\ : LocalMux
    port map (
            O => \N__42958\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__9444\ : InMux
    port map (
            O => \N__42951\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__9443\ : InMux
    port map (
            O => \N__42948\,
            I => \N__42945\
        );

    \I__9442\ : LocalMux
    port map (
            O => \N__42945\,
            I => \N__42942\
        );

    \I__9441\ : Span4Mux_v
    port map (
            O => \N__42942\,
            I => \N__42937\
        );

    \I__9440\ : InMux
    port map (
            O => \N__42941\,
            I => \N__42934\
        );

    \I__9439\ : InMux
    port map (
            O => \N__42940\,
            I => \N__42931\
        );

    \I__9438\ : Odrv4
    port map (
            O => \N__42937\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__9437\ : LocalMux
    port map (
            O => \N__42934\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__9436\ : LocalMux
    port map (
            O => \N__42931\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__9435\ : InMux
    port map (
            O => \N__42924\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__9434\ : InMux
    port map (
            O => \N__42921\,
            I => \bfn_17_21_0_\
        );

    \I__9433\ : CascadeMux
    port map (
            O => \N__42918\,
            I => \N__42915\
        );

    \I__9432\ : InMux
    port map (
            O => \N__42915\,
            I => \N__42912\
        );

    \I__9431\ : LocalMux
    port map (
            O => \N__42912\,
            I => \N__42909\
        );

    \I__9430\ : Span4Mux_v
    port map (
            O => \N__42909\,
            I => \N__42905\
        );

    \I__9429\ : InMux
    port map (
            O => \N__42908\,
            I => \N__42902\
        );

    \I__9428\ : Odrv4
    port map (
            O => \N__42905\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__9427\ : LocalMux
    port map (
            O => \N__42902\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__9426\ : InMux
    port map (
            O => \N__42897\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__9425\ : InMux
    port map (
            O => \N__42894\,
            I => \N__42891\
        );

    \I__9424\ : LocalMux
    port map (
            O => \N__42891\,
            I => \N__42886\
        );

    \I__9423\ : InMux
    port map (
            O => \N__42890\,
            I => \N__42881\
        );

    \I__9422\ : InMux
    port map (
            O => \N__42889\,
            I => \N__42881\
        );

    \I__9421\ : Span4Mux_v
    port map (
            O => \N__42886\,
            I => \N__42876\
        );

    \I__9420\ : LocalMux
    port map (
            O => \N__42881\,
            I => \N__42876\
        );

    \I__9419\ : Odrv4
    port map (
            O => \N__42876\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__9418\ : InMux
    port map (
            O => \N__42873\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__9417\ : InMux
    port map (
            O => \N__42870\,
            I => \N__42865\
        );

    \I__9416\ : InMux
    port map (
            O => \N__42869\,
            I => \N__42860\
        );

    \I__9415\ : InMux
    port map (
            O => \N__42868\,
            I => \N__42860\
        );

    \I__9414\ : LocalMux
    port map (
            O => \N__42865\,
            I => \N__42857\
        );

    \I__9413\ : LocalMux
    port map (
            O => \N__42860\,
            I => \N__42854\
        );

    \I__9412\ : Span4Mux_v
    port map (
            O => \N__42857\,
            I => \N__42849\
        );

    \I__9411\ : Span4Mux_h
    port map (
            O => \N__42854\,
            I => \N__42849\
        );

    \I__9410\ : Odrv4
    port map (
            O => \N__42849\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__9409\ : InMux
    port map (
            O => \N__42846\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__9408\ : InMux
    port map (
            O => \N__42843\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__9407\ : InMux
    port map (
            O => \N__42840\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__9406\ : InMux
    port map (
            O => \N__42837\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__9405\ : InMux
    port map (
            O => \N__42834\,
            I => \N__42831\
        );

    \I__9404\ : LocalMux
    port map (
            O => \N__42831\,
            I => \N__42826\
        );

    \I__9403\ : CascadeMux
    port map (
            O => \N__42830\,
            I => \N__42822\
        );

    \I__9402\ : CascadeMux
    port map (
            O => \N__42829\,
            I => \N__42819\
        );

    \I__9401\ : Span4Mux_h
    port map (
            O => \N__42826\,
            I => \N__42816\
        );

    \I__9400\ : InMux
    port map (
            O => \N__42825\,
            I => \N__42813\
        );

    \I__9399\ : InMux
    port map (
            O => \N__42822\,
            I => \N__42810\
        );

    \I__9398\ : InMux
    port map (
            O => \N__42819\,
            I => \N__42807\
        );

    \I__9397\ : Odrv4
    port map (
            O => \N__42816\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\
        );

    \I__9396\ : LocalMux
    port map (
            O => \N__42813\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\
        );

    \I__9395\ : LocalMux
    port map (
            O => \N__42810\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\
        );

    \I__9394\ : LocalMux
    port map (
            O => \N__42807\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\
        );

    \I__9393\ : InMux
    port map (
            O => \N__42798\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__9392\ : InMux
    port map (
            O => \N__42795\,
            I => \N__42792\
        );

    \I__9391\ : LocalMux
    port map (
            O => \N__42792\,
            I => \N__42788\
        );

    \I__9390\ : InMux
    port map (
            O => \N__42791\,
            I => \N__42785\
        );

    \I__9389\ : Odrv12
    port map (
            O => \N__42788\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__9388\ : LocalMux
    port map (
            O => \N__42785\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__9387\ : InMux
    port map (
            O => \N__42780\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__9386\ : InMux
    port map (
            O => \N__42777\,
            I => \N__42774\
        );

    \I__9385\ : LocalMux
    port map (
            O => \N__42774\,
            I => \N__42770\
        );

    \I__9384\ : InMux
    port map (
            O => \N__42773\,
            I => \N__42767\
        );

    \I__9383\ : Odrv12
    port map (
            O => \N__42770\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__9382\ : LocalMux
    port map (
            O => \N__42767\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__9381\ : InMux
    port map (
            O => \N__42762\,
            I => \bfn_17_20_0_\
        );

    \I__9380\ : InMux
    port map (
            O => \N__42759\,
            I => \N__42756\
        );

    \I__9379\ : LocalMux
    port map (
            O => \N__42756\,
            I => \N__42752\
        );

    \I__9378\ : CascadeMux
    port map (
            O => \N__42755\,
            I => \N__42749\
        );

    \I__9377\ : Span4Mux_h
    port map (
            O => \N__42752\,
            I => \N__42746\
        );

    \I__9376\ : InMux
    port map (
            O => \N__42749\,
            I => \N__42743\
        );

    \I__9375\ : Odrv4
    port map (
            O => \N__42746\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__9374\ : LocalMux
    port map (
            O => \N__42743\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__9373\ : InMux
    port map (
            O => \N__42738\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__9372\ : InMux
    port map (
            O => \N__42735\,
            I => \N__42732\
        );

    \I__9371\ : LocalMux
    port map (
            O => \N__42732\,
            I => \N__42729\
        );

    \I__9370\ : Span4Mux_v
    port map (
            O => \N__42729\,
            I => \N__42725\
        );

    \I__9369\ : InMux
    port map (
            O => \N__42728\,
            I => \N__42722\
        );

    \I__9368\ : Odrv4
    port map (
            O => \N__42725\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__42722\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__9366\ : InMux
    port map (
            O => \N__42717\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__9365\ : InMux
    port map (
            O => \N__42714\,
            I => \N__42711\
        );

    \I__9364\ : LocalMux
    port map (
            O => \N__42711\,
            I => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4\
        );

    \I__9363\ : CascadeMux
    port map (
            O => \N__42708\,
            I => \N__42705\
        );

    \I__9362\ : InMux
    port map (
            O => \N__42705\,
            I => \N__42702\
        );

    \I__9361\ : LocalMux
    port map (
            O => \N__42702\,
            I => \delay_measurement_inst.delay_tr_timer.N_344\
        );

    \I__9360\ : CascadeMux
    port map (
            O => \N__42699\,
            I => \delay_measurement_inst.delay_tr_timer.N_344_cascade_\
        );

    \I__9359\ : InMux
    port map (
            O => \N__42696\,
            I => \N__42693\
        );

    \I__9358\ : LocalMux
    port map (
            O => \N__42693\,
            I => \delay_measurement_inst.delay_tr_timer.N_347\
        );

    \I__9357\ : CascadeMux
    port map (
            O => \N__42690\,
            I => \delay_measurement_inst.delay_tr_timer.N_347_cascade_\
        );

    \I__9356\ : CascadeMux
    port map (
            O => \N__42687\,
            I => \delay_measurement_inst.delay_tr_timer.N_373_cascade_\
        );

    \I__9355\ : InMux
    port map (
            O => \N__42684\,
            I => \N__42681\
        );

    \I__9354\ : LocalMux
    port map (
            O => \N__42681\,
            I => \delay_measurement_inst.delay_tr_timer.N_351\
        );

    \I__9353\ : InMux
    port map (
            O => \N__42678\,
            I => \N__42675\
        );

    \I__9352\ : LocalMux
    port map (
            O => \N__42675\,
            I => \delay_measurement_inst.delay_tr_timer.N_353\
        );

    \I__9351\ : InMux
    port map (
            O => \N__42672\,
            I => \N__42668\
        );

    \I__9350\ : InMux
    port map (
            O => \N__42671\,
            I => \N__42665\
        );

    \I__9349\ : LocalMux
    port map (
            O => \N__42668\,
            I => \delay_measurement_inst.delay_tr_timer.N_348\
        );

    \I__9348\ : LocalMux
    port map (
            O => \N__42665\,
            I => \delay_measurement_inst.delay_tr_timer.N_348\
        );

    \I__9347\ : CascadeMux
    port map (
            O => \N__42660\,
            I => \N__42657\
        );

    \I__9346\ : InMux
    port map (
            O => \N__42657\,
            I => \N__42654\
        );

    \I__9345\ : LocalMux
    port map (
            O => \N__42654\,
            I => \N__42649\
        );

    \I__9344\ : InMux
    port map (
            O => \N__42653\,
            I => \N__42644\
        );

    \I__9343\ : InMux
    port map (
            O => \N__42652\,
            I => \N__42644\
        );

    \I__9342\ : Odrv12
    port map (
            O => \N__42649\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__9341\ : LocalMux
    port map (
            O => \N__42644\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__9340\ : InMux
    port map (
            O => \N__42639\,
            I => \N__42636\
        );

    \I__9339\ : LocalMux
    port map (
            O => \N__42636\,
            I => \N__42632\
        );

    \I__9338\ : InMux
    port map (
            O => \N__42635\,
            I => \N__42629\
        );

    \I__9337\ : Odrv4
    port map (
            O => \N__42632\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__9336\ : LocalMux
    port map (
            O => \N__42629\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__9335\ : InMux
    port map (
            O => \N__42624\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__9334\ : InMux
    port map (
            O => \N__42621\,
            I => \N__42618\
        );

    \I__9333\ : LocalMux
    port map (
            O => \N__42618\,
            I => \N__42614\
        );

    \I__9332\ : InMux
    port map (
            O => \N__42617\,
            I => \N__42611\
        );

    \I__9331\ : Odrv4
    port map (
            O => \N__42614\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__9330\ : LocalMux
    port map (
            O => \N__42611\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__9329\ : InMux
    port map (
            O => \N__42606\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__9328\ : CascadeMux
    port map (
            O => \N__42603\,
            I => \N__42600\
        );

    \I__9327\ : InMux
    port map (
            O => \N__42600\,
            I => \N__42596\
        );

    \I__9326\ : InMux
    port map (
            O => \N__42599\,
            I => \N__42593\
        );

    \I__9325\ : LocalMux
    port map (
            O => \N__42596\,
            I => \elapsed_time_ns_1_RNI3JIF91_0_29\
        );

    \I__9324\ : LocalMux
    port map (
            O => \N__42593\,
            I => \elapsed_time_ns_1_RNI3JIF91_0_29\
        );

    \I__9323\ : InMux
    port map (
            O => \N__42588\,
            I => \N__42585\
        );

    \I__9322\ : LocalMux
    port map (
            O => \N__42585\,
            I => \elapsed_time_ns_1_RNITCIF91_0_23\
        );

    \I__9321\ : CascadeMux
    port map (
            O => \N__42582\,
            I => \elapsed_time_ns_1_RNITCIF91_0_23_cascade_\
        );

    \I__9320\ : InMux
    port map (
            O => \N__42579\,
            I => \N__42575\
        );

    \I__9319\ : InMux
    port map (
            O => \N__42578\,
            I => \N__42572\
        );

    \I__9318\ : LocalMux
    port map (
            O => \N__42575\,
            I => \elapsed_time_ns_1_RNIUDIF91_0_24\
        );

    \I__9317\ : LocalMux
    port map (
            O => \N__42572\,
            I => \elapsed_time_ns_1_RNIUDIF91_0_24\
        );

    \I__9316\ : InMux
    port map (
            O => \N__42567\,
            I => \N__42564\
        );

    \I__9315\ : LocalMux
    port map (
            O => \N__42564\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15\
        );

    \I__9314\ : InMux
    port map (
            O => \N__42561\,
            I => \N__42557\
        );

    \I__9313\ : InMux
    port map (
            O => \N__42560\,
            I => \N__42551\
        );

    \I__9312\ : LocalMux
    port map (
            O => \N__42557\,
            I => \N__42548\
        );

    \I__9311\ : InMux
    port map (
            O => \N__42556\,
            I => \N__42545\
        );

    \I__9310\ : InMux
    port map (
            O => \N__42555\,
            I => \N__42542\
        );

    \I__9309\ : InMux
    port map (
            O => \N__42554\,
            I => \N__42539\
        );

    \I__9308\ : LocalMux
    port map (
            O => \N__42551\,
            I => \elapsed_time_ns_1_RNIA965M1_0_18\
        );

    \I__9307\ : Odrv12
    port map (
            O => \N__42548\,
            I => \elapsed_time_ns_1_RNIA965M1_0_18\
        );

    \I__9306\ : LocalMux
    port map (
            O => \N__42545\,
            I => \elapsed_time_ns_1_RNIA965M1_0_18\
        );

    \I__9305\ : LocalMux
    port map (
            O => \N__42542\,
            I => \elapsed_time_ns_1_RNIA965M1_0_18\
        );

    \I__9304\ : LocalMux
    port map (
            O => \N__42539\,
            I => \elapsed_time_ns_1_RNIA965M1_0_18\
        );

    \I__9303\ : CascadeMux
    port map (
            O => \N__42528\,
            I => \elapsed_time_ns_1_RNICG2591_0_4_cascade_\
        );

    \I__9302\ : InMux
    port map (
            O => \N__42525\,
            I => \N__42522\
        );

    \I__9301\ : LocalMux
    port map (
            O => \N__42522\,
            I => \N__42518\
        );

    \I__9300\ : InMux
    port map (
            O => \N__42521\,
            I => \N__42512\
        );

    \I__9299\ : Span4Mux_v
    port map (
            O => \N__42518\,
            I => \N__42509\
        );

    \I__9298\ : InMux
    port map (
            O => \N__42517\,
            I => \N__42506\
        );

    \I__9297\ : InMux
    port map (
            O => \N__42516\,
            I => \N__42503\
        );

    \I__9296\ : InMux
    port map (
            O => \N__42515\,
            I => \N__42500\
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__42512\,
            I => \elapsed_time_ns_1_RNI9865M1_0_17\
        );

    \I__9294\ : Odrv4
    port map (
            O => \N__42509\,
            I => \elapsed_time_ns_1_RNI9865M1_0_17\
        );

    \I__9293\ : LocalMux
    port map (
            O => \N__42506\,
            I => \elapsed_time_ns_1_RNI9865M1_0_17\
        );

    \I__9292\ : LocalMux
    port map (
            O => \N__42503\,
            I => \elapsed_time_ns_1_RNI9865M1_0_17\
        );

    \I__9291\ : LocalMux
    port map (
            O => \N__42500\,
            I => \elapsed_time_ns_1_RNI9865M1_0_17\
        );

    \I__9290\ : CascadeMux
    port map (
            O => \N__42489\,
            I => \N__42486\
        );

    \I__9289\ : InMux
    port map (
            O => \N__42486\,
            I => \N__42482\
        );

    \I__9288\ : InMux
    port map (
            O => \N__42485\,
            I => \N__42479\
        );

    \I__9287\ : LocalMux
    port map (
            O => \N__42482\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_9\
        );

    \I__9286\ : LocalMux
    port map (
            O => \N__42479\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_9\
        );

    \I__9285\ : CascadeMux
    port map (
            O => \N__42474\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2_cascade_\
        );

    \I__9284\ : CascadeMux
    port map (
            O => \N__42471\,
            I => \N__42468\
        );

    \I__9283\ : InMux
    port map (
            O => \N__42468\,
            I => \N__42464\
        );

    \I__9282\ : InMux
    port map (
            O => \N__42467\,
            I => \N__42461\
        );

    \I__9281\ : LocalMux
    port map (
            O => \N__42464\,
            I => \elapsed_time_ns_1_RNIRBJF91_0_30\
        );

    \I__9280\ : LocalMux
    port map (
            O => \N__42461\,
            I => \elapsed_time_ns_1_RNIRBJF91_0_30\
        );

    \I__9279\ : InMux
    port map (
            O => \N__42456\,
            I => \N__42453\
        );

    \I__9278\ : LocalMux
    port map (
            O => \N__42453\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16\
        );

    \I__9277\ : InMux
    port map (
            O => \N__42450\,
            I => \N__42446\
        );

    \I__9276\ : InMux
    port map (
            O => \N__42449\,
            I => \N__42443\
        );

    \I__9275\ : LocalMux
    port map (
            O => \N__42446\,
            I => \N__42439\
        );

    \I__9274\ : LocalMux
    port map (
            O => \N__42443\,
            I => \N__42436\
        );

    \I__9273\ : InMux
    port map (
            O => \N__42442\,
            I => \N__42433\
        );

    \I__9272\ : Span12Mux_v
    port map (
            O => \N__42439\,
            I => \N__42430\
        );

    \I__9271\ : Odrv4
    port map (
            O => \N__42436\,
            I => \delay_measurement_inst.N_363\
        );

    \I__9270\ : LocalMux
    port map (
            O => \N__42433\,
            I => \delay_measurement_inst.N_363\
        );

    \I__9269\ : Odrv12
    port map (
            O => \N__42430\,
            I => \delay_measurement_inst.N_363\
        );

    \I__9268\ : CascadeMux
    port map (
            O => \N__42423\,
            I => \N__42420\
        );

    \I__9267\ : InMux
    port map (
            O => \N__42420\,
            I => \N__42417\
        );

    \I__9266\ : LocalMux
    port map (
            O => \N__42417\,
            I => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0\
        );

    \I__9265\ : CascadeMux
    port map (
            O => \N__42414\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_\
        );

    \I__9264\ : CascadeMux
    port map (
            O => \N__42411\,
            I => \elapsed_time_ns_1_RNIBA65M1_0_19_cascade_\
        );

    \I__9263\ : CascadeMux
    port map (
            O => \N__42408\,
            I => \N__42405\
        );

    \I__9262\ : InMux
    port map (
            O => \N__42405\,
            I => \N__42401\
        );

    \I__9261\ : InMux
    port map (
            O => \N__42404\,
            I => \N__42398\
        );

    \I__9260\ : LocalMux
    port map (
            O => \N__42401\,
            I => \N__42392\
        );

    \I__9259\ : LocalMux
    port map (
            O => \N__42398\,
            I => \N__42392\
        );

    \I__9258\ : InMux
    port map (
            O => \N__42397\,
            I => \N__42389\
        );

    \I__9257\ : Span4Mux_h
    port map (
            O => \N__42392\,
            I => \N__42385\
        );

    \I__9256\ : LocalMux
    port map (
            O => \N__42389\,
            I => \N__42382\
        );

    \I__9255\ : InMux
    port map (
            O => \N__42388\,
            I => \N__42379\
        );

    \I__9254\ : Odrv4
    port map (
            O => \N__42385\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_9\
        );

    \I__9253\ : Odrv4
    port map (
            O => \N__42382\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_9\
        );

    \I__9252\ : LocalMux
    port map (
            O => \N__42379\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_9\
        );

    \I__9251\ : InMux
    port map (
            O => \N__42372\,
            I => \N__42369\
        );

    \I__9250\ : LocalMux
    port map (
            O => \N__42369\,
            I => \elapsed_time_ns_1_RNIQ9IF91_0_20\
        );

    \I__9249\ : CascadeMux
    port map (
            O => \N__42366\,
            I => \elapsed_time_ns_1_RNIQ9IF91_0_20_cascade_\
        );

    \I__9248\ : CascadeMux
    port map (
            O => \N__42363\,
            I => \N__42360\
        );

    \I__9247\ : InMux
    port map (
            O => \N__42360\,
            I => \N__42357\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__42357\,
            I => \N__42353\
        );

    \I__9245\ : InMux
    port map (
            O => \N__42356\,
            I => \N__42350\
        );

    \I__9244\ : Odrv4
    port map (
            O => \N__42353\,
            I => \elapsed_time_ns_1_RNIRAIF91_0_21\
        );

    \I__9243\ : LocalMux
    port map (
            O => \N__42350\,
            I => \elapsed_time_ns_1_RNIRAIF91_0_21\
        );

    \I__9242\ : InMux
    port map (
            O => \N__42345\,
            I => \N__42342\
        );

    \I__9241\ : LocalMux
    port map (
            O => \N__42342\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15\
        );

    \I__9240\ : CascadeMux
    port map (
            O => \N__42339\,
            I => \N__42336\
        );

    \I__9239\ : InMux
    port map (
            O => \N__42336\,
            I => \N__42331\
        );

    \I__9238\ : CascadeMux
    port map (
            O => \N__42335\,
            I => \N__42328\
        );

    \I__9237\ : InMux
    port map (
            O => \N__42334\,
            I => \N__42325\
        );

    \I__9236\ : LocalMux
    port map (
            O => \N__42331\,
            I => \N__42322\
        );

    \I__9235\ : InMux
    port map (
            O => \N__42328\,
            I => \N__42318\
        );

    \I__9234\ : LocalMux
    port map (
            O => \N__42325\,
            I => \N__42315\
        );

    \I__9233\ : Span4Mux_h
    port map (
            O => \N__42322\,
            I => \N__42312\
        );

    \I__9232\ : InMux
    port map (
            O => \N__42321\,
            I => \N__42309\
        );

    \I__9231\ : LocalMux
    port map (
            O => \N__42318\,
            I => \elapsed_time_ns_1_RNIQ8HF91_0_11\
        );

    \I__9230\ : Odrv4
    port map (
            O => \N__42315\,
            I => \elapsed_time_ns_1_RNIQ8HF91_0_11\
        );

    \I__9229\ : Odrv4
    port map (
            O => \N__42312\,
            I => \elapsed_time_ns_1_RNIQ8HF91_0_11\
        );

    \I__9228\ : LocalMux
    port map (
            O => \N__42309\,
            I => \elapsed_time_ns_1_RNIQ8HF91_0_11\
        );

    \I__9227\ : InMux
    port map (
            O => \N__42300\,
            I => \N__42297\
        );

    \I__9226\ : LocalMux
    port map (
            O => \N__42297\,
            I => \N__42294\
        );

    \I__9225\ : Span4Mux_h
    port map (
            O => \N__42294\,
            I => \N__42291\
        );

    \I__9224\ : Odrv4
    port map (
            O => \N__42291\,
            I => \current_shift_inst.un38_control_input_0_s1_30\
        );

    \I__9223\ : InMux
    port map (
            O => \N__42288\,
            I => \current_shift_inst.un38_control_input_cry_29_s1\
        );

    \I__9222\ : InMux
    port map (
            O => \N__42285\,
            I => \current_shift_inst.un38_control_input_cry_30_s1\
        );

    \I__9221\ : CascadeMux
    port map (
            O => \N__42282\,
            I => \N__42279\
        );

    \I__9220\ : InMux
    port map (
            O => \N__42279\,
            I => \N__42276\
        );

    \I__9219\ : LocalMux
    port map (
            O => \N__42276\,
            I => \N__42273\
        );

    \I__9218\ : Span4Mux_h
    port map (
            O => \N__42273\,
            I => \N__42270\
        );

    \I__9217\ : Odrv4
    port map (
            O => \N__42270\,
            I => \current_shift_inst.un38_control_input_0_s1_31\
        );

    \I__9216\ : CascadeMux
    port map (
            O => \N__42267\,
            I => \N__42263\
        );

    \I__9215\ : CascadeMux
    port map (
            O => \N__42266\,
            I => \N__42260\
        );

    \I__9214\ : InMux
    port map (
            O => \N__42263\,
            I => \N__42257\
        );

    \I__9213\ : InMux
    port map (
            O => \N__42260\,
            I => \N__42254\
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__42257\,
            I => \N__42248\
        );

    \I__9211\ : LocalMux
    port map (
            O => \N__42254\,
            I => \N__42248\
        );

    \I__9210\ : CascadeMux
    port map (
            O => \N__42253\,
            I => \N__42245\
        );

    \I__9209\ : Span4Mux_v
    port map (
            O => \N__42248\,
            I => \N__42242\
        );

    \I__9208\ : InMux
    port map (
            O => \N__42245\,
            I => \N__42239\
        );

    \I__9207\ : Odrv4
    port map (
            O => \N__42242\,
            I => \elapsed_time_ns_1_RNIP7HF91_0_10\
        );

    \I__9206\ : LocalMux
    port map (
            O => \N__42239\,
            I => \elapsed_time_ns_1_RNIP7HF91_0_10\
        );

    \I__9205\ : InMux
    port map (
            O => \N__42234\,
            I => \N__42231\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__42231\,
            I => \N__42226\
        );

    \I__9203\ : InMux
    port map (
            O => \N__42230\,
            I => \N__42222\
        );

    \I__9202\ : InMux
    port map (
            O => \N__42229\,
            I => \N__42219\
        );

    \I__9201\ : Span12Mux_s11_v
    port map (
            O => \N__42226\,
            I => \N__42216\
        );

    \I__9200\ : InMux
    port map (
            O => \N__42225\,
            I => \N__42213\
        );

    \I__9199\ : LocalMux
    port map (
            O => \N__42222\,
            I => \elapsed_time_ns_1_RNIR9HF91_0_12\
        );

    \I__9198\ : LocalMux
    port map (
            O => \N__42219\,
            I => \elapsed_time_ns_1_RNIR9HF91_0_12\
        );

    \I__9197\ : Odrv12
    port map (
            O => \N__42216\,
            I => \elapsed_time_ns_1_RNIR9HF91_0_12\
        );

    \I__9196\ : LocalMux
    port map (
            O => \N__42213\,
            I => \elapsed_time_ns_1_RNIR9HF91_0_12\
        );

    \I__9195\ : CascadeMux
    port map (
            O => \N__42204\,
            I => \N__42200\
        );

    \I__9194\ : InMux
    port map (
            O => \N__42203\,
            I => \N__42196\
        );

    \I__9193\ : InMux
    port map (
            O => \N__42200\,
            I => \N__42193\
        );

    \I__9192\ : InMux
    port map (
            O => \N__42199\,
            I => \N__42190\
        );

    \I__9191\ : LocalMux
    port map (
            O => \N__42196\,
            I => \elapsed_time_ns_1_RNISAHF91_0_13\
        );

    \I__9190\ : LocalMux
    port map (
            O => \N__42193\,
            I => \elapsed_time_ns_1_RNISAHF91_0_13\
        );

    \I__9189\ : LocalMux
    port map (
            O => \N__42190\,
            I => \elapsed_time_ns_1_RNISAHF91_0_13\
        );

    \I__9188\ : CascadeMux
    port map (
            O => \N__42183\,
            I => \elapsed_time_ns_1_RNIP7HF91_0_10_cascade_\
        );

    \I__9187\ : CascadeMux
    port map (
            O => \N__42180\,
            I => \N__42177\
        );

    \I__9186\ : InMux
    port map (
            O => \N__42177\,
            I => \N__42174\
        );

    \I__9185\ : LocalMux
    port map (
            O => \N__42174\,
            I => \N__42171\
        );

    \I__9184\ : Span4Mux_v
    port map (
            O => \N__42171\,
            I => \N__42165\
        );

    \I__9183\ : InMux
    port map (
            O => \N__42170\,
            I => \N__42162\
        );

    \I__9182\ : InMux
    port map (
            O => \N__42169\,
            I => \N__42159\
        );

    \I__9181\ : InMux
    port map (
            O => \N__42168\,
            I => \N__42155\
        );

    \I__9180\ : Sp12to4
    port map (
            O => \N__42165\,
            I => \N__42152\
        );

    \I__9179\ : LocalMux
    port map (
            O => \N__42162\,
            I => \N__42149\
        );

    \I__9178\ : LocalMux
    port map (
            O => \N__42159\,
            I => \N__42146\
        );

    \I__9177\ : InMux
    port map (
            O => \N__42158\,
            I => \N__42143\
        );

    \I__9176\ : LocalMux
    port map (
            O => \N__42155\,
            I => \elapsed_time_ns_1_RNI6565M1_0_14\
        );

    \I__9175\ : Odrv12
    port map (
            O => \N__42152\,
            I => \elapsed_time_ns_1_RNI6565M1_0_14\
        );

    \I__9174\ : Odrv4
    port map (
            O => \N__42149\,
            I => \elapsed_time_ns_1_RNI6565M1_0_14\
        );

    \I__9173\ : Odrv4
    port map (
            O => \N__42146\,
            I => \elapsed_time_ns_1_RNI6565M1_0_14\
        );

    \I__9172\ : LocalMux
    port map (
            O => \N__42143\,
            I => \elapsed_time_ns_1_RNI6565M1_0_14\
        );

    \I__9171\ : CascadeMux
    port map (
            O => \N__42132\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2_cascade_\
        );

    \I__9170\ : InMux
    port map (
            O => \N__42129\,
            I => \N__42124\
        );

    \I__9169\ : InMux
    port map (
            O => \N__42128\,
            I => \N__42120\
        );

    \I__9168\ : InMux
    port map (
            O => \N__42127\,
            I => \N__42117\
        );

    \I__9167\ : LocalMux
    port map (
            O => \N__42124\,
            I => \N__42114\
        );

    \I__9166\ : InMux
    port map (
            O => \N__42123\,
            I => \N__42111\
        );

    \I__9165\ : LocalMux
    port map (
            O => \N__42120\,
            I => \N__42106\
        );

    \I__9164\ : LocalMux
    port map (
            O => \N__42117\,
            I => \N__42106\
        );

    \I__9163\ : Span4Mux_v
    port map (
            O => \N__42114\,
            I => \N__42102\
        );

    \I__9162\ : LocalMux
    port map (
            O => \N__42111\,
            I => \N__42097\
        );

    \I__9161\ : Span4Mux_h
    port map (
            O => \N__42106\,
            I => \N__42097\
        );

    \I__9160\ : InMux
    port map (
            O => \N__42105\,
            I => \N__42094\
        );

    \I__9159\ : Odrv4
    port map (
            O => \N__42102\,
            I => \elapsed_time_ns_1_RNIQENQL1_0_9\
        );

    \I__9158\ : Odrv4
    port map (
            O => \N__42097\,
            I => \elapsed_time_ns_1_RNIQENQL1_0_9\
        );

    \I__9157\ : LocalMux
    port map (
            O => \N__42094\,
            I => \elapsed_time_ns_1_RNIQENQL1_0_9\
        );

    \I__9156\ : CascadeMux
    port map (
            O => \N__42087\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_0_6_cascade_\
        );

    \I__9155\ : CascadeMux
    port map (
            O => \N__42084\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_\
        );

    \I__9154\ : CascadeMux
    port map (
            O => \N__42081\,
            I => \elapsed_time_ns_1_RNIK8NQL1_0_3_cascade_\
        );

    \I__9153\ : CascadeMux
    port map (
            O => \N__42078\,
            I => \N__42075\
        );

    \I__9152\ : InMux
    port map (
            O => \N__42075\,
            I => \N__42072\
        );

    \I__9151\ : LocalMux
    port map (
            O => \N__42072\,
            I => \N__42069\
        );

    \I__9150\ : Span4Mux_v
    port map (
            O => \N__42069\,
            I => \N__42066\
        );

    \I__9149\ : Odrv4
    port map (
            O => \N__42066\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\
        );

    \I__9148\ : InMux
    port map (
            O => \N__42063\,
            I => \N__42060\
        );

    \I__9147\ : LocalMux
    port map (
            O => \N__42060\,
            I => \N__42057\
        );

    \I__9146\ : Span4Mux_h
    port map (
            O => \N__42057\,
            I => \N__42054\
        );

    \I__9145\ : Odrv4
    port map (
            O => \N__42054\,
            I => \current_shift_inst.un38_control_input_0_s1_22\
        );

    \I__9144\ : InMux
    port map (
            O => \N__42051\,
            I => \current_shift_inst.un38_control_input_cry_21_s1\
        );

    \I__9143\ : InMux
    port map (
            O => \N__42048\,
            I => \N__42045\
        );

    \I__9142\ : LocalMux
    port map (
            O => \N__42045\,
            I => \N__42042\
        );

    \I__9141\ : Span4Mux_h
    port map (
            O => \N__42042\,
            I => \N__42039\
        );

    \I__9140\ : Odrv4
    port map (
            O => \N__42039\,
            I => \current_shift_inst.un38_control_input_0_s1_23\
        );

    \I__9139\ : InMux
    port map (
            O => \N__42036\,
            I => \current_shift_inst.un38_control_input_cry_22_s1\
        );

    \I__9138\ : CascadeMux
    port map (
            O => \N__42033\,
            I => \N__42030\
        );

    \I__9137\ : InMux
    port map (
            O => \N__42030\,
            I => \N__42027\
        );

    \I__9136\ : LocalMux
    port map (
            O => \N__42027\,
            I => \N__42024\
        );

    \I__9135\ : Odrv12
    port map (
            O => \N__42024\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\
        );

    \I__9134\ : InMux
    port map (
            O => \N__42021\,
            I => \N__42018\
        );

    \I__9133\ : LocalMux
    port map (
            O => \N__42018\,
            I => \N__42015\
        );

    \I__9132\ : Span4Mux_h
    port map (
            O => \N__42015\,
            I => \N__42012\
        );

    \I__9131\ : Odrv4
    port map (
            O => \N__42012\,
            I => \current_shift_inst.un38_control_input_0_s1_24\
        );

    \I__9130\ : InMux
    port map (
            O => \N__42009\,
            I => \bfn_17_14_0_\
        );

    \I__9129\ : InMux
    port map (
            O => \N__42006\,
            I => \N__42003\
        );

    \I__9128\ : LocalMux
    port map (
            O => \N__42003\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\
        );

    \I__9127\ : InMux
    port map (
            O => \N__42000\,
            I => \N__41997\
        );

    \I__9126\ : LocalMux
    port map (
            O => \N__41997\,
            I => \N__41994\
        );

    \I__9125\ : Span4Mux_h
    port map (
            O => \N__41994\,
            I => \N__41991\
        );

    \I__9124\ : Odrv4
    port map (
            O => \N__41991\,
            I => \current_shift_inst.un38_control_input_0_s1_25\
        );

    \I__9123\ : InMux
    port map (
            O => \N__41988\,
            I => \current_shift_inst.un38_control_input_cry_24_s1\
        );

    \I__9122\ : CascadeMux
    port map (
            O => \N__41985\,
            I => \N__41982\
        );

    \I__9121\ : InMux
    port map (
            O => \N__41982\,
            I => \N__41979\
        );

    \I__9120\ : LocalMux
    port map (
            O => \N__41979\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\
        );

    \I__9119\ : CascadeMux
    port map (
            O => \N__41976\,
            I => \N__41973\
        );

    \I__9118\ : InMux
    port map (
            O => \N__41973\,
            I => \N__41970\
        );

    \I__9117\ : LocalMux
    port map (
            O => \N__41970\,
            I => \N__41967\
        );

    \I__9116\ : Span4Mux_v
    port map (
            O => \N__41967\,
            I => \N__41964\
        );

    \I__9115\ : Odrv4
    port map (
            O => \N__41964\,
            I => \current_shift_inst.un38_control_input_0_s1_26\
        );

    \I__9114\ : InMux
    port map (
            O => \N__41961\,
            I => \current_shift_inst.un38_control_input_cry_25_s1\
        );

    \I__9113\ : InMux
    port map (
            O => \N__41958\,
            I => \N__41955\
        );

    \I__9112\ : LocalMux
    port map (
            O => \N__41955\,
            I => \N__41952\
        );

    \I__9111\ : Span4Mux_v
    port map (
            O => \N__41952\,
            I => \N__41949\
        );

    \I__9110\ : Odrv4
    port map (
            O => \N__41949\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\
        );

    \I__9109\ : InMux
    port map (
            O => \N__41946\,
            I => \N__41943\
        );

    \I__9108\ : LocalMux
    port map (
            O => \N__41943\,
            I => \N__41940\
        );

    \I__9107\ : Span4Mux_v
    port map (
            O => \N__41940\,
            I => \N__41937\
        );

    \I__9106\ : Odrv4
    port map (
            O => \N__41937\,
            I => \current_shift_inst.un38_control_input_0_s1_27\
        );

    \I__9105\ : InMux
    port map (
            O => \N__41934\,
            I => \current_shift_inst.un38_control_input_cry_26_s1\
        );

    \I__9104\ : CascadeMux
    port map (
            O => \N__41931\,
            I => \N__41928\
        );

    \I__9103\ : InMux
    port map (
            O => \N__41928\,
            I => \N__41925\
        );

    \I__9102\ : LocalMux
    port map (
            O => \N__41925\,
            I => \N__41922\
        );

    \I__9101\ : Span4Mux_v
    port map (
            O => \N__41922\,
            I => \N__41919\
        );

    \I__9100\ : Odrv4
    port map (
            O => \N__41919\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\
        );

    \I__9099\ : InMux
    port map (
            O => \N__41916\,
            I => \N__41913\
        );

    \I__9098\ : LocalMux
    port map (
            O => \N__41913\,
            I => \N__41910\
        );

    \I__9097\ : Span4Mux_h
    port map (
            O => \N__41910\,
            I => \N__41907\
        );

    \I__9096\ : Odrv4
    port map (
            O => \N__41907\,
            I => \current_shift_inst.un38_control_input_0_s1_28\
        );

    \I__9095\ : InMux
    port map (
            O => \N__41904\,
            I => \current_shift_inst.un38_control_input_cry_27_s1\
        );

    \I__9094\ : InMux
    port map (
            O => \N__41901\,
            I => \N__41898\
        );

    \I__9093\ : LocalMux
    port map (
            O => \N__41898\,
            I => \N__41895\
        );

    \I__9092\ : Span4Mux_h
    port map (
            O => \N__41895\,
            I => \N__41892\
        );

    \I__9091\ : Odrv4
    port map (
            O => \N__41892\,
            I => \current_shift_inst.un38_control_input_0_s1_29\
        );

    \I__9090\ : InMux
    port map (
            O => \N__41889\,
            I => \current_shift_inst.un38_control_input_cry_28_s1\
        );

    \I__9089\ : InMux
    port map (
            O => \N__41886\,
            I => \N__41883\
        );

    \I__9088\ : LocalMux
    port map (
            O => \N__41883\,
            I => \N__41880\
        );

    \I__9087\ : Span4Mux_v
    port map (
            O => \N__41880\,
            I => \N__41877\
        );

    \I__9086\ : Odrv4
    port map (
            O => \N__41877\,
            I => \current_shift_inst.un38_control_input_0_s1_20\
        );

    \I__9085\ : InMux
    port map (
            O => \N__41874\,
            I => \current_shift_inst.un38_control_input_cry_19_s1\
        );

    \I__9084\ : InMux
    port map (
            O => \N__41871\,
            I => \N__41868\
        );

    \I__9083\ : LocalMux
    port map (
            O => \N__41868\,
            I => \N__41865\
        );

    \I__9082\ : Odrv4
    port map (
            O => \N__41865\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\
        );

    \I__9081\ : InMux
    port map (
            O => \N__41862\,
            I => \N__41859\
        );

    \I__9080\ : LocalMux
    port map (
            O => \N__41859\,
            I => \N__41856\
        );

    \I__9079\ : Span4Mux_h
    port map (
            O => \N__41856\,
            I => \N__41853\
        );

    \I__9078\ : Odrv4
    port map (
            O => \N__41853\,
            I => \current_shift_inst.un38_control_input_0_s1_21\
        );

    \I__9077\ : InMux
    port map (
            O => \N__41850\,
            I => \current_shift_inst.un38_control_input_cry_20_s1\
        );

    \I__9076\ : InMux
    port map (
            O => \N__41847\,
            I => \N__41844\
        );

    \I__9075\ : LocalMux
    port map (
            O => \N__41844\,
            I => \N__41841\
        );

    \I__9074\ : Odrv12
    port map (
            O => \N__41841\,
            I => \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\
        );

    \I__9073\ : InMux
    port map (
            O => \N__41838\,
            I => \N__41835\
        );

    \I__9072\ : LocalMux
    port map (
            O => \N__41835\,
            I => \N__41832\
        );

    \I__9071\ : Odrv12
    port map (
            O => \N__41832\,
            I => \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\
        );

    \I__9070\ : InMux
    port map (
            O => \N__41829\,
            I => \N__41826\
        );

    \I__9069\ : LocalMux
    port map (
            O => \N__41826\,
            I => \N__41823\
        );

    \I__9068\ : Span4Mux_v
    port map (
            O => \N__41823\,
            I => \N__41820\
        );

    \I__9067\ : Odrv4
    port map (
            O => \N__41820\,
            I => \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\
        );

    \I__9066\ : InMux
    port map (
            O => \N__41817\,
            I => \N__41814\
        );

    \I__9065\ : LocalMux
    port map (
            O => \N__41814\,
            I => \N__41811\
        );

    \I__9064\ : Odrv4
    port map (
            O => \N__41811\,
            I => \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\
        );

    \I__9063\ : CascadeMux
    port map (
            O => \N__41808\,
            I => \N__41805\
        );

    \I__9062\ : InMux
    port map (
            O => \N__41805\,
            I => \N__41802\
        );

    \I__9061\ : LocalMux
    port map (
            O => \N__41802\,
            I => \N__41799\
        );

    \I__9060\ : Odrv12
    port map (
            O => \N__41799\,
            I => \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\
        );

    \I__9059\ : InMux
    port map (
            O => \N__41796\,
            I => \N__41793\
        );

    \I__9058\ : LocalMux
    port map (
            O => \N__41793\,
            I => \N__41790\
        );

    \I__9057\ : Odrv12
    port map (
            O => \N__41790\,
            I => \current_shift_inst.un4_control_input_1_axb_29\
        );

    \I__9056\ : InMux
    port map (
            O => \N__41787\,
            I => \current_shift_inst.un4_control_input_1_cry_28\
        );

    \I__9055\ : InMux
    port map (
            O => \N__41784\,
            I => \current_shift_inst.un4_control_input1_31\
        );

    \I__9054\ : CascadeMux
    port map (
            O => \N__41781\,
            I => \N__41777\
        );

    \I__9053\ : CascadeMux
    port map (
            O => \N__41780\,
            I => \N__41774\
        );

    \I__9052\ : InMux
    port map (
            O => \N__41777\,
            I => \N__41771\
        );

    \I__9051\ : InMux
    port map (
            O => \N__41774\,
            I => \N__41768\
        );

    \I__9050\ : LocalMux
    port map (
            O => \N__41771\,
            I => \N__41765\
        );

    \I__9049\ : LocalMux
    port map (
            O => \N__41768\,
            I => \N__41762\
        );

    \I__9048\ : Span4Mux_v
    port map (
            O => \N__41765\,
            I => \N__41756\
        );

    \I__9047\ : Span4Mux_h
    port map (
            O => \N__41762\,
            I => \N__41756\
        );

    \I__9046\ : CascadeMux
    port map (
            O => \N__41761\,
            I => \N__41753\
        );

    \I__9045\ : Span4Mux_h
    port map (
            O => \N__41756\,
            I => \N__41749\
        );

    \I__9044\ : InMux
    port map (
            O => \N__41753\,
            I => \N__41744\
        );

    \I__9043\ : InMux
    port map (
            O => \N__41752\,
            I => \N__41744\
        );

    \I__9042\ : Odrv4
    port map (
            O => \N__41749\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__9041\ : LocalMux
    port map (
            O => \N__41744\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__9040\ : InMux
    port map (
            O => \N__41739\,
            I => \N__41736\
        );

    \I__9039\ : LocalMux
    port map (
            O => \N__41736\,
            I => \N__41731\
        );

    \I__9038\ : InMux
    port map (
            O => \N__41735\,
            I => \N__41728\
        );

    \I__9037\ : InMux
    port map (
            O => \N__41734\,
            I => \N__41725\
        );

    \I__9036\ : Span4Mux_v
    port map (
            O => \N__41731\,
            I => \N__41720\
        );

    \I__9035\ : LocalMux
    port map (
            O => \N__41728\,
            I => \N__41720\
        );

    \I__9034\ : LocalMux
    port map (
            O => \N__41725\,
            I => \N__41717\
        );

    \I__9033\ : Span4Mux_h
    port map (
            O => \N__41720\,
            I => \N__41714\
        );

    \I__9032\ : Odrv4
    port map (
            O => \N__41717\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__9031\ : Odrv4
    port map (
            O => \N__41714\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__9030\ : CascadeMux
    port map (
            O => \N__41709\,
            I => \N__41705\
        );

    \I__9029\ : InMux
    port map (
            O => \N__41708\,
            I => \N__41702\
        );

    \I__9028\ : InMux
    port map (
            O => \N__41705\,
            I => \N__41698\
        );

    \I__9027\ : LocalMux
    port map (
            O => \N__41702\,
            I => \N__41694\
        );

    \I__9026\ : InMux
    port map (
            O => \N__41701\,
            I => \N__41691\
        );

    \I__9025\ : LocalMux
    port map (
            O => \N__41698\,
            I => \N__41688\
        );

    \I__9024\ : InMux
    port map (
            O => \N__41697\,
            I => \N__41685\
        );

    \I__9023\ : Span4Mux_v
    port map (
            O => \N__41694\,
            I => \N__41680\
        );

    \I__9022\ : LocalMux
    port map (
            O => \N__41691\,
            I => \N__41680\
        );

    \I__9021\ : Span4Mux_v
    port map (
            O => \N__41688\,
            I => \N__41677\
        );

    \I__9020\ : LocalMux
    port map (
            O => \N__41685\,
            I => \N__41674\
        );

    \I__9019\ : Span4Mux_h
    port map (
            O => \N__41680\,
            I => \N__41671\
        );

    \I__9018\ : Span4Mux_h
    port map (
            O => \N__41677\,
            I => \N__41666\
        );

    \I__9017\ : Span4Mux_h
    port map (
            O => \N__41674\,
            I => \N__41666\
        );

    \I__9016\ : Odrv4
    port map (
            O => \N__41671\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__9015\ : Odrv4
    port map (
            O => \N__41666\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__9014\ : InMux
    port map (
            O => \N__41661\,
            I => \N__41658\
        );

    \I__9013\ : LocalMux
    port map (
            O => \N__41658\,
            I => \N__41653\
        );

    \I__9012\ : InMux
    port map (
            O => \N__41657\,
            I => \N__41650\
        );

    \I__9011\ : InMux
    port map (
            O => \N__41656\,
            I => \N__41647\
        );

    \I__9010\ : Span4Mux_v
    port map (
            O => \N__41653\,
            I => \N__41642\
        );

    \I__9009\ : LocalMux
    port map (
            O => \N__41650\,
            I => \N__41642\
        );

    \I__9008\ : LocalMux
    port map (
            O => \N__41647\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__9007\ : Odrv4
    port map (
            O => \N__41642\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__9006\ : InMux
    port map (
            O => \N__41637\,
            I => \N__41634\
        );

    \I__9005\ : LocalMux
    port map (
            O => \N__41634\,
            I => \N__41630\
        );

    \I__9004\ : InMux
    port map (
            O => \N__41633\,
            I => \N__41627\
        );

    \I__9003\ : Span4Mux_h
    port map (
            O => \N__41630\,
            I => \N__41624\
        );

    \I__9002\ : LocalMux
    port map (
            O => \N__41627\,
            I => \N__41621\
        );

    \I__9001\ : Odrv4
    port map (
            O => \N__41624\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__9000\ : Odrv4
    port map (
            O => \N__41621\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__8999\ : InMux
    port map (
            O => \N__41616\,
            I => \N__41613\
        );

    \I__8998\ : LocalMux
    port map (
            O => \N__41613\,
            I => \N__41609\
        );

    \I__8997\ : CascadeMux
    port map (
            O => \N__41612\,
            I => \N__41606\
        );

    \I__8996\ : Span4Mux_v
    port map (
            O => \N__41609\,
            I => \N__41603\
        );

    \I__8995\ : InMux
    port map (
            O => \N__41606\,
            I => \N__41600\
        );

    \I__8994\ : Odrv4
    port map (
            O => \N__41603\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__8993\ : LocalMux
    port map (
            O => \N__41600\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__8992\ : CascadeMux
    port map (
            O => \N__41595\,
            I => \N__41592\
        );

    \I__8991\ : InMux
    port map (
            O => \N__41592\,
            I => \N__41589\
        );

    \I__8990\ : LocalMux
    port map (
            O => \N__41589\,
            I => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\
        );

    \I__8989\ : InMux
    port map (
            O => \N__41586\,
            I => \N__41583\
        );

    \I__8988\ : LocalMux
    port map (
            O => \N__41583\,
            I => \N__41580\
        );

    \I__8987\ : Span4Mux_v
    port map (
            O => \N__41580\,
            I => \N__41577\
        );

    \I__8986\ : Odrv4
    port map (
            O => \N__41577\,
            I => \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\
        );

    \I__8985\ : CascadeMux
    port map (
            O => \N__41574\,
            I => \N__41571\
        );

    \I__8984\ : InMux
    port map (
            O => \N__41571\,
            I => \N__41568\
        );

    \I__8983\ : LocalMux
    port map (
            O => \N__41568\,
            I => \N__41565\
        );

    \I__8982\ : Span4Mux_v
    port map (
            O => \N__41565\,
            I => \N__41562\
        );

    \I__8981\ : Odrv4
    port map (
            O => \N__41562\,
            I => \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\
        );

    \I__8980\ : InMux
    port map (
            O => \N__41559\,
            I => \N__41556\
        );

    \I__8979\ : LocalMux
    port map (
            O => \N__41556\,
            I => \N__41553\
        );

    \I__8978\ : Odrv4
    port map (
            O => \N__41553\,
            I => \current_shift_inst.un4_control_input_1_axb_21\
        );

    \I__8977\ : InMux
    port map (
            O => \N__41550\,
            I => \N__41541\
        );

    \I__8976\ : InMux
    port map (
            O => \N__41549\,
            I => \N__41541\
        );

    \I__8975\ : InMux
    port map (
            O => \N__41548\,
            I => \N__41541\
        );

    \I__8974\ : LocalMux
    port map (
            O => \N__41541\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__8973\ : InMux
    port map (
            O => \N__41538\,
            I => \current_shift_inst.un4_control_input_1_cry_20\
        );

    \I__8972\ : InMux
    port map (
            O => \N__41535\,
            I => \N__41532\
        );

    \I__8971\ : LocalMux
    port map (
            O => \N__41532\,
            I => \N__41529\
        );

    \I__8970\ : Odrv4
    port map (
            O => \N__41529\,
            I => \current_shift_inst.un4_control_input_1_axb_22\
        );

    \I__8969\ : InMux
    port map (
            O => \N__41526\,
            I => \current_shift_inst.un4_control_input_1_cry_21\
        );

    \I__8968\ : InMux
    port map (
            O => \N__41523\,
            I => \N__41520\
        );

    \I__8967\ : LocalMux
    port map (
            O => \N__41520\,
            I => \N__41517\
        );

    \I__8966\ : Odrv4
    port map (
            O => \N__41517\,
            I => \current_shift_inst.un4_control_input_1_axb_23\
        );

    \I__8965\ : InMux
    port map (
            O => \N__41514\,
            I => \current_shift_inst.un4_control_input_1_cry_22\
        );

    \I__8964\ : InMux
    port map (
            O => \N__41511\,
            I => \N__41508\
        );

    \I__8963\ : LocalMux
    port map (
            O => \N__41508\,
            I => \N__41505\
        );

    \I__8962\ : Span4Mux_h
    port map (
            O => \N__41505\,
            I => \N__41502\
        );

    \I__8961\ : Span4Mux_h
    port map (
            O => \N__41502\,
            I => \N__41499\
        );

    \I__8960\ : Odrv4
    port map (
            O => \N__41499\,
            I => \current_shift_inst.un4_control_input_1_axb_24\
        );

    \I__8959\ : InMux
    port map (
            O => \N__41496\,
            I => \current_shift_inst.un4_control_input_1_cry_23\
        );

    \I__8958\ : InMux
    port map (
            O => \N__41493\,
            I => \N__41490\
        );

    \I__8957\ : LocalMux
    port map (
            O => \N__41490\,
            I => \N__41487\
        );

    \I__8956\ : Odrv4
    port map (
            O => \N__41487\,
            I => \current_shift_inst.un4_control_input_1_axb_25\
        );

    \I__8955\ : CascadeMux
    port map (
            O => \N__41484\,
            I => \N__41481\
        );

    \I__8954\ : InMux
    port map (
            O => \N__41481\,
            I => \N__41477\
        );

    \I__8953\ : InMux
    port map (
            O => \N__41480\,
            I => \N__41474\
        );

    \I__8952\ : LocalMux
    port map (
            O => \N__41477\,
            I => \N__41468\
        );

    \I__8951\ : LocalMux
    port map (
            O => \N__41474\,
            I => \N__41468\
        );

    \I__8950\ : InMux
    port map (
            O => \N__41473\,
            I => \N__41465\
        );

    \I__8949\ : Span4Mux_v
    port map (
            O => \N__41468\,
            I => \N__41462\
        );

    \I__8948\ : LocalMux
    port map (
            O => \N__41465\,
            I => \N__41459\
        );

    \I__8947\ : Odrv4
    port map (
            O => \N__41462\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__8946\ : Odrv12
    port map (
            O => \N__41459\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__8945\ : InMux
    port map (
            O => \N__41454\,
            I => \bfn_17_10_0_\
        );

    \I__8944\ : InMux
    port map (
            O => \N__41451\,
            I => \N__41448\
        );

    \I__8943\ : LocalMux
    port map (
            O => \N__41448\,
            I => \N__41445\
        );

    \I__8942\ : Odrv12
    port map (
            O => \N__41445\,
            I => \current_shift_inst.un4_control_input_1_axb_26\
        );

    \I__8941\ : CascadeMux
    port map (
            O => \N__41442\,
            I => \N__41439\
        );

    \I__8940\ : InMux
    port map (
            O => \N__41439\,
            I => \N__41435\
        );

    \I__8939\ : InMux
    port map (
            O => \N__41438\,
            I => \N__41432\
        );

    \I__8938\ : LocalMux
    port map (
            O => \N__41435\,
            I => \N__41428\
        );

    \I__8937\ : LocalMux
    port map (
            O => \N__41432\,
            I => \N__41425\
        );

    \I__8936\ : InMux
    port map (
            O => \N__41431\,
            I => \N__41422\
        );

    \I__8935\ : Sp12to4
    port map (
            O => \N__41428\,
            I => \N__41419\
        );

    \I__8934\ : Span4Mux_v
    port map (
            O => \N__41425\,
            I => \N__41414\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__41422\,
            I => \N__41414\
        );

    \I__8932\ : Odrv12
    port map (
            O => \N__41419\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__8931\ : Odrv4
    port map (
            O => \N__41414\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__8930\ : InMux
    port map (
            O => \N__41409\,
            I => \current_shift_inst.un4_control_input_1_cry_25\
        );

    \I__8929\ : InMux
    port map (
            O => \N__41406\,
            I => \N__41403\
        );

    \I__8928\ : LocalMux
    port map (
            O => \N__41403\,
            I => \N__41400\
        );

    \I__8927\ : Odrv12
    port map (
            O => \N__41400\,
            I => \current_shift_inst.un4_control_input_1_axb_27\
        );

    \I__8926\ : CascadeMux
    port map (
            O => \N__41397\,
            I => \N__41394\
        );

    \I__8925\ : InMux
    port map (
            O => \N__41394\,
            I => \N__41391\
        );

    \I__8924\ : LocalMux
    port map (
            O => \N__41391\,
            I => \N__41387\
        );

    \I__8923\ : CascadeMux
    port map (
            O => \N__41390\,
            I => \N__41384\
        );

    \I__8922\ : Span4Mux_v
    port map (
            O => \N__41387\,
            I => \N__41380\
        );

    \I__8921\ : InMux
    port map (
            O => \N__41384\,
            I => \N__41375\
        );

    \I__8920\ : InMux
    port map (
            O => \N__41383\,
            I => \N__41375\
        );

    \I__8919\ : Odrv4
    port map (
            O => \N__41380\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__8918\ : LocalMux
    port map (
            O => \N__41375\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__8917\ : InMux
    port map (
            O => \N__41370\,
            I => \current_shift_inst.un4_control_input_1_cry_26\
        );

    \I__8916\ : InMux
    port map (
            O => \N__41367\,
            I => \N__41364\
        );

    \I__8915\ : LocalMux
    port map (
            O => \N__41364\,
            I => \N__41361\
        );

    \I__8914\ : Odrv12
    port map (
            O => \N__41361\,
            I => \current_shift_inst.un4_control_input_1_axb_28\
        );

    \I__8913\ : InMux
    port map (
            O => \N__41358\,
            I => \N__41349\
        );

    \I__8912\ : InMux
    port map (
            O => \N__41357\,
            I => \N__41349\
        );

    \I__8911\ : InMux
    port map (
            O => \N__41356\,
            I => \N__41349\
        );

    \I__8910\ : LocalMux
    port map (
            O => \N__41349\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__8909\ : InMux
    port map (
            O => \N__41346\,
            I => \current_shift_inst.un4_control_input_1_cry_27\
        );

    \I__8908\ : InMux
    port map (
            O => \N__41343\,
            I => \N__41340\
        );

    \I__8907\ : LocalMux
    port map (
            O => \N__41340\,
            I => \current_shift_inst.un4_control_input_1_axb_13\
        );

    \I__8906\ : InMux
    port map (
            O => \N__41337\,
            I => \current_shift_inst.un4_control_input_1_cry_12\
        );

    \I__8905\ : InMux
    port map (
            O => \N__41334\,
            I => \current_shift_inst.un4_control_input_1_cry_13\
        );

    \I__8904\ : InMux
    port map (
            O => \N__41331\,
            I => \N__41328\
        );

    \I__8903\ : LocalMux
    port map (
            O => \N__41328\,
            I => \N__41325\
        );

    \I__8902\ : Span4Mux_h
    port map (
            O => \N__41325\,
            I => \N__41322\
        );

    \I__8901\ : Odrv4
    port map (
            O => \N__41322\,
            I => \current_shift_inst.un4_control_input_1_axb_15\
        );

    \I__8900\ : InMux
    port map (
            O => \N__41319\,
            I => \current_shift_inst.un4_control_input_1_cry_14\
        );

    \I__8899\ : InMux
    port map (
            O => \N__41316\,
            I => \N__41313\
        );

    \I__8898\ : LocalMux
    port map (
            O => \N__41313\,
            I => \N__41310\
        );

    \I__8897\ : Odrv12
    port map (
            O => \N__41310\,
            I => \current_shift_inst.un4_control_input_1_axb_16\
        );

    \I__8896\ : InMux
    port map (
            O => \N__41307\,
            I => \current_shift_inst.un4_control_input_1_cry_15\
        );

    \I__8895\ : InMux
    port map (
            O => \N__41304\,
            I => \N__41301\
        );

    \I__8894\ : LocalMux
    port map (
            O => \N__41301\,
            I => \N__41298\
        );

    \I__8893\ : Odrv4
    port map (
            O => \N__41298\,
            I => \current_shift_inst.un4_control_input_1_axb_17\
        );

    \I__8892\ : InMux
    port map (
            O => \N__41295\,
            I => \bfn_17_9_0_\
        );

    \I__8891\ : InMux
    port map (
            O => \N__41292\,
            I => \N__41289\
        );

    \I__8890\ : LocalMux
    port map (
            O => \N__41289\,
            I => \N__41286\
        );

    \I__8889\ : Odrv12
    port map (
            O => \N__41286\,
            I => \current_shift_inst.un4_control_input_1_axb_18\
        );

    \I__8888\ : InMux
    port map (
            O => \N__41283\,
            I => \current_shift_inst.un4_control_input_1_cry_17\
        );

    \I__8887\ : InMux
    port map (
            O => \N__41280\,
            I => \N__41277\
        );

    \I__8886\ : LocalMux
    port map (
            O => \N__41277\,
            I => \N__41274\
        );

    \I__8885\ : Odrv12
    port map (
            O => \N__41274\,
            I => \current_shift_inst.un4_control_input_1_axb_19\
        );

    \I__8884\ : InMux
    port map (
            O => \N__41271\,
            I => \current_shift_inst.un4_control_input_1_cry_18\
        );

    \I__8883\ : InMux
    port map (
            O => \N__41268\,
            I => \current_shift_inst.un4_control_input_1_cry_19\
        );

    \I__8882\ : InMux
    port map (
            O => \N__41265\,
            I => \N__41262\
        );

    \I__8881\ : LocalMux
    port map (
            O => \N__41262\,
            I => \N__41259\
        );

    \I__8880\ : Odrv4
    port map (
            O => \N__41259\,
            I => \current_shift_inst.un4_control_input_1_axb_5\
        );

    \I__8879\ : InMux
    port map (
            O => \N__41256\,
            I => \N__41253\
        );

    \I__8878\ : LocalMux
    port map (
            O => \N__41253\,
            I => \N__41248\
        );

    \I__8877\ : InMux
    port map (
            O => \N__41252\,
            I => \N__41245\
        );

    \I__8876\ : InMux
    port map (
            O => \N__41251\,
            I => \N__41242\
        );

    \I__8875\ : Odrv4
    port map (
            O => \N__41248\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__8874\ : LocalMux
    port map (
            O => \N__41245\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__8873\ : LocalMux
    port map (
            O => \N__41242\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__8872\ : InMux
    port map (
            O => \N__41235\,
            I => \current_shift_inst.un4_control_input_1_cry_4\
        );

    \I__8871\ : InMux
    port map (
            O => \N__41232\,
            I => \N__41229\
        );

    \I__8870\ : LocalMux
    port map (
            O => \N__41229\,
            I => \N__41226\
        );

    \I__8869\ : Span4Mux_h
    port map (
            O => \N__41226\,
            I => \N__41223\
        );

    \I__8868\ : Odrv4
    port map (
            O => \N__41223\,
            I => \current_shift_inst.un4_control_input_1_axb_6\
        );

    \I__8867\ : InMux
    port map (
            O => \N__41220\,
            I => \current_shift_inst.un4_control_input_1_cry_5\
        );

    \I__8866\ : InMux
    port map (
            O => \N__41217\,
            I => \N__41214\
        );

    \I__8865\ : LocalMux
    port map (
            O => \N__41214\,
            I => \N__41211\
        );

    \I__8864\ : Odrv4
    port map (
            O => \N__41211\,
            I => \current_shift_inst.un4_control_input_1_axb_7\
        );

    \I__8863\ : InMux
    port map (
            O => \N__41208\,
            I => \N__41205\
        );

    \I__8862\ : LocalMux
    port map (
            O => \N__41205\,
            I => \N__41200\
        );

    \I__8861\ : InMux
    port map (
            O => \N__41204\,
            I => \N__41197\
        );

    \I__8860\ : InMux
    port map (
            O => \N__41203\,
            I => \N__41194\
        );

    \I__8859\ : Span4Mux_v
    port map (
            O => \N__41200\,
            I => \N__41189\
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__41197\,
            I => \N__41189\
        );

    \I__8857\ : LocalMux
    port map (
            O => \N__41194\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__8856\ : Odrv4
    port map (
            O => \N__41189\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__8855\ : InMux
    port map (
            O => \N__41184\,
            I => \current_shift_inst.un4_control_input_1_cry_6\
        );

    \I__8854\ : InMux
    port map (
            O => \N__41181\,
            I => \N__41178\
        );

    \I__8853\ : LocalMux
    port map (
            O => \N__41178\,
            I => \N__41175\
        );

    \I__8852\ : Odrv4
    port map (
            O => \N__41175\,
            I => \current_shift_inst.un4_control_input_1_axb_8\
        );

    \I__8851\ : InMux
    port map (
            O => \N__41172\,
            I => \current_shift_inst.un4_control_input_1_cry_7\
        );

    \I__8850\ : InMux
    port map (
            O => \N__41169\,
            I => \N__41166\
        );

    \I__8849\ : LocalMux
    port map (
            O => \N__41166\,
            I => \N__41163\
        );

    \I__8848\ : Span4Mux_h
    port map (
            O => \N__41163\,
            I => \N__41160\
        );

    \I__8847\ : Odrv4
    port map (
            O => \N__41160\,
            I => \current_shift_inst.un4_control_input_1_axb_9\
        );

    \I__8846\ : InMux
    port map (
            O => \N__41157\,
            I => \N__41153\
        );

    \I__8845\ : CascadeMux
    port map (
            O => \N__41156\,
            I => \N__41150\
        );

    \I__8844\ : LocalMux
    port map (
            O => \N__41153\,
            I => \N__41146\
        );

    \I__8843\ : InMux
    port map (
            O => \N__41150\,
            I => \N__41141\
        );

    \I__8842\ : InMux
    port map (
            O => \N__41149\,
            I => \N__41141\
        );

    \I__8841\ : Span4Mux_h
    port map (
            O => \N__41146\,
            I => \N__41138\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__41141\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__8839\ : Odrv4
    port map (
            O => \N__41138\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__8838\ : InMux
    port map (
            O => \N__41133\,
            I => \bfn_17_8_0_\
        );

    \I__8837\ : InMux
    port map (
            O => \N__41130\,
            I => \N__41127\
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__41127\,
            I => \current_shift_inst.un4_control_input_1_axb_10\
        );

    \I__8835\ : InMux
    port map (
            O => \N__41124\,
            I => \current_shift_inst.un4_control_input_1_cry_9\
        );

    \I__8834\ : InMux
    port map (
            O => \N__41121\,
            I => \N__41118\
        );

    \I__8833\ : LocalMux
    port map (
            O => \N__41118\,
            I => \N__41115\
        );

    \I__8832\ : Span4Mux_h
    port map (
            O => \N__41115\,
            I => \N__41112\
        );

    \I__8831\ : Odrv4
    port map (
            O => \N__41112\,
            I => \current_shift_inst.un4_control_input_1_axb_11\
        );

    \I__8830\ : InMux
    port map (
            O => \N__41109\,
            I => \current_shift_inst.un4_control_input_1_cry_10\
        );

    \I__8829\ : InMux
    port map (
            O => \N__41106\,
            I => \current_shift_inst.un4_control_input_1_cry_11\
        );

    \I__8828\ : CascadeMux
    port map (
            O => \N__41103\,
            I => \N__41099\
        );

    \I__8827\ : CascadeMux
    port map (
            O => \N__41102\,
            I => \N__41096\
        );

    \I__8826\ : InMux
    port map (
            O => \N__41099\,
            I => \N__41093\
        );

    \I__8825\ : InMux
    port map (
            O => \N__41096\,
            I => \N__41090\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__41093\,
            I => \N__41085\
        );

    \I__8823\ : LocalMux
    port map (
            O => \N__41090\,
            I => \N__41082\
        );

    \I__8822\ : InMux
    port map (
            O => \N__41089\,
            I => \N__41077\
        );

    \I__8821\ : InMux
    port map (
            O => \N__41088\,
            I => \N__41077\
        );

    \I__8820\ : Span4Mux_h
    port map (
            O => \N__41085\,
            I => \N__41074\
        );

    \I__8819\ : Span4Mux_v
    port map (
            O => \N__41082\,
            I => \N__41069\
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__41077\,
            I => \N__41069\
        );

    \I__8817\ : Odrv4
    port map (
            O => \N__41074\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__8816\ : Odrv4
    port map (
            O => \N__41069\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__8815\ : InMux
    port map (
            O => \N__41064\,
            I => \N__41060\
        );

    \I__8814\ : InMux
    port map (
            O => \N__41063\,
            I => \N__41057\
        );

    \I__8813\ : LocalMux
    port map (
            O => \N__41060\,
            I => \N__41053\
        );

    \I__8812\ : LocalMux
    port map (
            O => \N__41057\,
            I => \N__41050\
        );

    \I__8811\ : CascadeMux
    port map (
            O => \N__41056\,
            I => \N__41046\
        );

    \I__8810\ : Span4Mux_h
    port map (
            O => \N__41053\,
            I => \N__41041\
        );

    \I__8809\ : Span4Mux_v
    port map (
            O => \N__41050\,
            I => \N__41041\
        );

    \I__8808\ : InMux
    port map (
            O => \N__41049\,
            I => \N__41038\
        );

    \I__8807\ : InMux
    port map (
            O => \N__41046\,
            I => \N__41035\
        );

    \I__8806\ : Odrv4
    port map (
            O => \N__41041\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__8805\ : LocalMux
    port map (
            O => \N__41038\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__41035\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__8803\ : InMux
    port map (
            O => \N__41028\,
            I => \N__41025\
        );

    \I__8802\ : LocalMux
    port map (
            O => \N__41025\,
            I => \N__41022\
        );

    \I__8801\ : Odrv4
    port map (
            O => \N__41022\,
            I => \current_shift_inst.un4_control_input_1_axb_2\
        );

    \I__8800\ : InMux
    port map (
            O => \N__41019\,
            I => \N__41013\
        );

    \I__8799\ : InMux
    port map (
            O => \N__41018\,
            I => \N__41013\
        );

    \I__8798\ : LocalMux
    port map (
            O => \N__41013\,
            I => \N__41010\
        );

    \I__8797\ : Span4Mux_v
    port map (
            O => \N__41010\,
            I => \N__41006\
        );

    \I__8796\ : InMux
    port map (
            O => \N__41009\,
            I => \N__41003\
        );

    \I__8795\ : Odrv4
    port map (
            O => \N__41006\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__8794\ : LocalMux
    port map (
            O => \N__41003\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__8793\ : InMux
    port map (
            O => \N__40998\,
            I => \current_shift_inst.un4_control_input_1_cry_1\
        );

    \I__8792\ : InMux
    port map (
            O => \N__40995\,
            I => \N__40992\
        );

    \I__8791\ : LocalMux
    port map (
            O => \N__40992\,
            I => \N__40989\
        );

    \I__8790\ : Odrv12
    port map (
            O => \N__40989\,
            I => \current_shift_inst.un4_control_input_1_axb_3\
        );

    \I__8789\ : InMux
    port map (
            O => \N__40986\,
            I => \N__40983\
        );

    \I__8788\ : LocalMux
    port map (
            O => \N__40983\,
            I => \N__40980\
        );

    \I__8787\ : Span4Mux_v
    port map (
            O => \N__40980\,
            I => \N__40975\
        );

    \I__8786\ : InMux
    port map (
            O => \N__40979\,
            I => \N__40972\
        );

    \I__8785\ : InMux
    port map (
            O => \N__40978\,
            I => \N__40969\
        );

    \I__8784\ : Odrv4
    port map (
            O => \N__40975\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__8783\ : LocalMux
    port map (
            O => \N__40972\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__8782\ : LocalMux
    port map (
            O => \N__40969\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__8781\ : InMux
    port map (
            O => \N__40962\,
            I => \current_shift_inst.un4_control_input_1_cry_2\
        );

    \I__8780\ : InMux
    port map (
            O => \N__40959\,
            I => \N__40956\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__40956\,
            I => \N__40953\
        );

    \I__8778\ : Odrv4
    port map (
            O => \N__40953\,
            I => \current_shift_inst.un4_control_input_1_axb_4\
        );

    \I__8777\ : CascadeMux
    port map (
            O => \N__40950\,
            I => \N__40947\
        );

    \I__8776\ : InMux
    port map (
            O => \N__40947\,
            I => \N__40944\
        );

    \I__8775\ : LocalMux
    port map (
            O => \N__40944\,
            I => \N__40939\
        );

    \I__8774\ : InMux
    port map (
            O => \N__40943\,
            I => \N__40934\
        );

    \I__8773\ : InMux
    port map (
            O => \N__40942\,
            I => \N__40934\
        );

    \I__8772\ : Span4Mux_h
    port map (
            O => \N__40939\,
            I => \N__40931\
        );

    \I__8771\ : LocalMux
    port map (
            O => \N__40934\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__8770\ : Odrv4
    port map (
            O => \N__40931\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__8769\ : InMux
    port map (
            O => \N__40926\,
            I => \current_shift_inst.un4_control_input_1_cry_3\
        );

    \I__8768\ : InMux
    port map (
            O => \N__40923\,
            I => \N__40918\
        );

    \I__8767\ : InMux
    port map (
            O => \N__40922\,
            I => \N__40915\
        );

    \I__8766\ : InMux
    port map (
            O => \N__40921\,
            I => \N__40911\
        );

    \I__8765\ : LocalMux
    port map (
            O => \N__40918\,
            I => \N__40908\
        );

    \I__8764\ : LocalMux
    port map (
            O => \N__40915\,
            I => \N__40905\
        );

    \I__8763\ : InMux
    port map (
            O => \N__40914\,
            I => \N__40902\
        );

    \I__8762\ : LocalMux
    port map (
            O => \N__40911\,
            I => \N__40899\
        );

    \I__8761\ : Span12Mux_v
    port map (
            O => \N__40908\,
            I => \N__40896\
        );

    \I__8760\ : Span12Mux_v
    port map (
            O => \N__40905\,
            I => \N__40893\
        );

    \I__8759\ : LocalMux
    port map (
            O => \N__40902\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__8758\ : Odrv4
    port map (
            O => \N__40899\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__8757\ : Odrv12
    port map (
            O => \N__40896\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__8756\ : Odrv12
    port map (
            O => \N__40893\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__8755\ : InMux
    port map (
            O => \N__40884\,
            I => \N__40881\
        );

    \I__8754\ : LocalMux
    port map (
            O => \N__40881\,
            I => \N__40878\
        );

    \I__8753\ : Span4Mux_h
    port map (
            O => \N__40878\,
            I => \N__40875\
        );

    \I__8752\ : Odrv4
    port map (
            O => \N__40875\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_5\
        );

    \I__8751\ : CascadeMux
    port map (
            O => \N__40872\,
            I => \N__40869\
        );

    \I__8750\ : InMux
    port map (
            O => \N__40869\,
            I => \N__40861\
        );

    \I__8749\ : InMux
    port map (
            O => \N__40868\,
            I => \N__40855\
        );

    \I__8748\ : InMux
    port map (
            O => \N__40867\,
            I => \N__40850\
        );

    \I__8747\ : InMux
    port map (
            O => \N__40866\,
            I => \N__40850\
        );

    \I__8746\ : InMux
    port map (
            O => \N__40865\,
            I => \N__40845\
        );

    \I__8745\ : InMux
    port map (
            O => \N__40864\,
            I => \N__40845\
        );

    \I__8744\ : LocalMux
    port map (
            O => \N__40861\,
            I => \N__40842\
        );

    \I__8743\ : CascadeMux
    port map (
            O => \N__40860\,
            I => \N__40839\
        );

    \I__8742\ : CascadeMux
    port map (
            O => \N__40859\,
            I => \N__40835\
        );

    \I__8741\ : CascadeMux
    port map (
            O => \N__40858\,
            I => \N__40832\
        );

    \I__8740\ : LocalMux
    port map (
            O => \N__40855\,
            I => \N__40828\
        );

    \I__8739\ : LocalMux
    port map (
            O => \N__40850\,
            I => \N__40825\
        );

    \I__8738\ : LocalMux
    port map (
            O => \N__40845\,
            I => \N__40820\
        );

    \I__8737\ : Span4Mux_v
    port map (
            O => \N__40842\,
            I => \N__40820\
        );

    \I__8736\ : InMux
    port map (
            O => \N__40839\,
            I => \N__40815\
        );

    \I__8735\ : InMux
    port map (
            O => \N__40838\,
            I => \N__40815\
        );

    \I__8734\ : InMux
    port map (
            O => \N__40835\,
            I => \N__40812\
        );

    \I__8733\ : InMux
    port map (
            O => \N__40832\,
            I => \N__40807\
        );

    \I__8732\ : InMux
    port map (
            O => \N__40831\,
            I => \N__40807\
        );

    \I__8731\ : Span4Mux_h
    port map (
            O => \N__40828\,
            I => \N__40804\
        );

    \I__8730\ : Span4Mux_v
    port map (
            O => \N__40825\,
            I => \N__40801\
        );

    \I__8729\ : Span4Mux_v
    port map (
            O => \N__40820\,
            I => \N__40798\
        );

    \I__8728\ : LocalMux
    port map (
            O => \N__40815\,
            I => \phase_controller_inst1.stoper_tr.N_242\
        );

    \I__8727\ : LocalMux
    port map (
            O => \N__40812\,
            I => \phase_controller_inst1.stoper_tr.N_242\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__40807\,
            I => \phase_controller_inst1.stoper_tr.N_242\
        );

    \I__8725\ : Odrv4
    port map (
            O => \N__40804\,
            I => \phase_controller_inst1.stoper_tr.N_242\
        );

    \I__8724\ : Odrv4
    port map (
            O => \N__40801\,
            I => \phase_controller_inst1.stoper_tr.N_242\
        );

    \I__8723\ : Odrv4
    port map (
            O => \N__40798\,
            I => \phase_controller_inst1.stoper_tr.N_242\
        );

    \I__8722\ : InMux
    port map (
            O => \N__40785\,
            I => \N__40782\
        );

    \I__8721\ : LocalMux
    port map (
            O => \N__40782\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\
        );

    \I__8720\ : CascadeMux
    port map (
            O => \N__40779\,
            I => \N__40776\
        );

    \I__8719\ : InMux
    port map (
            O => \N__40776\,
            I => \N__40770\
        );

    \I__8718\ : InMux
    port map (
            O => \N__40775\,
            I => \N__40770\
        );

    \I__8717\ : LocalMux
    port map (
            O => \N__40770\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\
        );

    \I__8716\ : CascadeMux
    port map (
            O => \N__40767\,
            I => \N__40763\
        );

    \I__8715\ : CascadeMux
    port map (
            O => \N__40766\,
            I => \N__40760\
        );

    \I__8714\ : InMux
    port map (
            O => \N__40763\,
            I => \N__40757\
        );

    \I__8713\ : InMux
    port map (
            O => \N__40760\,
            I => \N__40754\
        );

    \I__8712\ : LocalMux
    port map (
            O => \N__40757\,
            I => \N__40751\
        );

    \I__8711\ : LocalMux
    port map (
            O => \N__40754\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\
        );

    \I__8710\ : Odrv4
    port map (
            O => \N__40751\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\
        );

    \I__8709\ : InMux
    port map (
            O => \N__40746\,
            I => \N__40742\
        );

    \I__8708\ : InMux
    port map (
            O => \N__40745\,
            I => \N__40739\
        );

    \I__8707\ : LocalMux
    port map (
            O => \N__40742\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__8706\ : LocalMux
    port map (
            O => \N__40739\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__8705\ : InMux
    port map (
            O => \N__40734\,
            I => \N__40730\
        );

    \I__8704\ : InMux
    port map (
            O => \N__40733\,
            I => \N__40727\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__40730\,
            I => \N__40723\
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__40727\,
            I => \N__40720\
        );

    \I__8701\ : InMux
    port map (
            O => \N__40726\,
            I => \N__40717\
        );

    \I__8700\ : Span4Mux_h
    port map (
            O => \N__40723\,
            I => \N__40714\
        );

    \I__8699\ : Odrv4
    port map (
            O => \N__40720\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__8698\ : LocalMux
    port map (
            O => \N__40717\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__8697\ : Odrv4
    port map (
            O => \N__40714\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__8696\ : CascadeMux
    port map (
            O => \N__40707\,
            I => \N__40704\
        );

    \I__8695\ : InMux
    port map (
            O => \N__40704\,
            I => \N__40699\
        );

    \I__8694\ : InMux
    port map (
            O => \N__40703\,
            I => \N__40696\
        );

    \I__8693\ : CascadeMux
    port map (
            O => \N__40702\,
            I => \N__40693\
        );

    \I__8692\ : LocalMux
    port map (
            O => \N__40699\,
            I => \N__40689\
        );

    \I__8691\ : LocalMux
    port map (
            O => \N__40696\,
            I => \N__40686\
        );

    \I__8690\ : InMux
    port map (
            O => \N__40693\,
            I => \N__40681\
        );

    \I__8689\ : InMux
    port map (
            O => \N__40692\,
            I => \N__40681\
        );

    \I__8688\ : Span4Mux_v
    port map (
            O => \N__40689\,
            I => \N__40678\
        );

    \I__8687\ : Span4Mux_h
    port map (
            O => \N__40686\,
            I => \N__40673\
        );

    \I__8686\ : LocalMux
    port map (
            O => \N__40681\,
            I => \N__40673\
        );

    \I__8685\ : Odrv4
    port map (
            O => \N__40678\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__8684\ : Odrv4
    port map (
            O => \N__40673\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__8683\ : InMux
    port map (
            O => \N__40668\,
            I => \N__40661\
        );

    \I__8682\ : InMux
    port map (
            O => \N__40667\,
            I => \N__40661\
        );

    \I__8681\ : InMux
    port map (
            O => \N__40666\,
            I => \N__40658\
        );

    \I__8680\ : LocalMux
    port map (
            O => \N__40661\,
            I => \N__40655\
        );

    \I__8679\ : LocalMux
    port map (
            O => \N__40658\,
            I => \N__40652\
        );

    \I__8678\ : Span4Mux_v
    port map (
            O => \N__40655\,
            I => \N__40648\
        );

    \I__8677\ : Span4Mux_v
    port map (
            O => \N__40652\,
            I => \N__40645\
        );

    \I__8676\ : InMux
    port map (
            O => \N__40651\,
            I => \N__40642\
        );

    \I__8675\ : Odrv4
    port map (
            O => \N__40648\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__8674\ : Odrv4
    port map (
            O => \N__40645\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__8673\ : LocalMux
    port map (
            O => \N__40642\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__8672\ : CascadeMux
    port map (
            O => \N__40635\,
            I => \N__40632\
        );

    \I__8671\ : InMux
    port map (
            O => \N__40632\,
            I => \N__40628\
        );

    \I__8670\ : InMux
    port map (
            O => \N__40631\,
            I => \N__40625\
        );

    \I__8669\ : LocalMux
    port map (
            O => \N__40628\,
            I => \delay_measurement_inst.delay_tr_timer.N_382\
        );

    \I__8668\ : LocalMux
    port map (
            O => \N__40625\,
            I => \delay_measurement_inst.delay_tr_timer.N_382\
        );

    \I__8667\ : CascadeMux
    port map (
            O => \N__40620\,
            I => \delay_measurement_inst.delay_tr_timer.N_382_cascade_\
        );

    \I__8666\ : InMux
    port map (
            O => \N__40617\,
            I => \N__40613\
        );

    \I__8665\ : InMux
    port map (
            O => \N__40616\,
            I => \N__40610\
        );

    \I__8664\ : LocalMux
    port map (
            O => \N__40613\,
            I => \delay_measurement_inst.delay_tr_timer.N_371\
        );

    \I__8663\ : LocalMux
    port map (
            O => \N__40610\,
            I => \delay_measurement_inst.delay_tr_timer.N_371\
        );

    \I__8662\ : InMux
    port map (
            O => \N__40605\,
            I => \N__40599\
        );

    \I__8661\ : InMux
    port map (
            O => \N__40604\,
            I => \N__40599\
        );

    \I__8660\ : LocalMux
    port map (
            O => \N__40599\,
            I => \delay_measurement_inst.delay_tr_timer.N_356\
        );

    \I__8659\ : InMux
    port map (
            O => \N__40596\,
            I => \N__40593\
        );

    \I__8658\ : LocalMux
    port map (
            O => \N__40593\,
            I => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5\
        );

    \I__8657\ : CascadeMux
    port map (
            O => \N__40590\,
            I => \delay_measurement_inst.delay_tr_timer.N_351_cascade_\
        );

    \I__8656\ : InMux
    port map (
            O => \N__40587\,
            I => \N__40583\
        );

    \I__8655\ : CascadeMux
    port map (
            O => \N__40586\,
            I => \N__40580\
        );

    \I__8654\ : LocalMux
    port map (
            O => \N__40583\,
            I => \N__40577\
        );

    \I__8653\ : InMux
    port map (
            O => \N__40580\,
            I => \N__40574\
        );

    \I__8652\ : Odrv4
    port map (
            O => \N__40577\,
            I => \delay_measurement_inst.delay_tr_timer.N_378\
        );

    \I__8651\ : LocalMux
    port map (
            O => \N__40574\,
            I => \delay_measurement_inst.delay_tr_timer.N_378\
        );

    \I__8650\ : InMux
    port map (
            O => \N__40569\,
            I => \N__40566\
        );

    \I__8649\ : LocalMux
    port map (
            O => \N__40566\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_4\
        );

    \I__8648\ : InMux
    port map (
            O => \N__40563\,
            I => \N__40560\
        );

    \I__8647\ : LocalMux
    port map (
            O => \N__40560\,
            I => \N__40556\
        );

    \I__8646\ : InMux
    port map (
            O => \N__40559\,
            I => \N__40553\
        );

    \I__8645\ : Odrv4
    port map (
            O => \N__40556\,
            I => \delay_measurement_inst.delay_tr_timer.N_360\
        );

    \I__8644\ : LocalMux
    port map (
            O => \N__40553\,
            I => \delay_measurement_inst.delay_tr_timer.N_360\
        );

    \I__8643\ : CascadeMux
    port map (
            O => \N__40548\,
            I => \delay_measurement_inst.delay_tr9_cascade_\
        );

    \I__8642\ : InMux
    port map (
            O => \N__40545\,
            I => \N__40542\
        );

    \I__8641\ : LocalMux
    port map (
            O => \N__40542\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0\
        );

    \I__8640\ : InMux
    port map (
            O => \N__40539\,
            I => \N__40533\
        );

    \I__8639\ : InMux
    port map (
            O => \N__40538\,
            I => \N__40533\
        );

    \I__8638\ : LocalMux
    port map (
            O => \N__40533\,
            I => \delay_measurement_inst.delay_tr_timer.N_390\
        );

    \I__8637\ : CascadeMux
    port map (
            O => \N__40530\,
            I => \delay_measurement_inst.delay_tr_timer.N_390_cascade_\
        );

    \I__8636\ : CascadeMux
    port map (
            O => \N__40527\,
            I => \delay_measurement_inst.delay_tr_timer.N_391_cascade_\
        );

    \I__8635\ : CascadeMux
    port map (
            O => \N__40524\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_\
        );

    \I__8634\ : CascadeMux
    port map (
            O => \N__40521\,
            I => \elapsed_time_ns_1_RNI6565M1_0_14_cascade_\
        );

    \I__8633\ : InMux
    port map (
            O => \N__40518\,
            I => \N__40515\
        );

    \I__8632\ : LocalMux
    port map (
            O => \N__40515\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14\
        );

    \I__8631\ : InMux
    port map (
            O => \N__40512\,
            I => \N__40509\
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__40509\,
            I => \elapsed_time_ns_1_RNIVEIF91_0_25\
        );

    \I__8629\ : InMux
    port map (
            O => \N__40506\,
            I => \N__40500\
        );

    \I__8628\ : InMux
    port map (
            O => \N__40505\,
            I => \N__40500\
        );

    \I__8627\ : LocalMux
    port map (
            O => \N__40500\,
            I => \elapsed_time_ns_1_RNI1HIF91_0_27\
        );

    \I__8626\ : CascadeMux
    port map (
            O => \N__40497\,
            I => \elapsed_time_ns_1_RNIVEIF91_0_25_cascade_\
        );

    \I__8625\ : InMux
    port map (
            O => \N__40494\,
            I => \N__40488\
        );

    \I__8624\ : InMux
    port map (
            O => \N__40493\,
            I => \N__40488\
        );

    \I__8623\ : LocalMux
    port map (
            O => \N__40488\,
            I => \elapsed_time_ns_1_RNISBIF91_0_22\
        );

    \I__8622\ : CascadeMux
    port map (
            O => \N__40485\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15_cascade_\
        );

    \I__8621\ : InMux
    port map (
            O => \N__40482\,
            I => \N__40476\
        );

    \I__8620\ : InMux
    port map (
            O => \N__40481\,
            I => \N__40476\
        );

    \I__8619\ : LocalMux
    port map (
            O => \N__40476\,
            I => \elapsed_time_ns_1_RNI2IIF91_0_28\
        );

    \I__8618\ : CascadeMux
    port map (
            O => \N__40473\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_\
        );

    \I__8617\ : InMux
    port map (
            O => \N__40470\,
            I => \N__40466\
        );

    \I__8616\ : InMux
    port map (
            O => \N__40469\,
            I => \N__40463\
        );

    \I__8615\ : LocalMux
    port map (
            O => \N__40466\,
            I => \elapsed_time_ns_1_RNI0GIF91_0_26\
        );

    \I__8614\ : LocalMux
    port map (
            O => \N__40463\,
            I => \elapsed_time_ns_1_RNI0GIF91_0_26\
        );

    \I__8613\ : InMux
    port map (
            O => \N__40458\,
            I => \N__40455\
        );

    \I__8612\ : LocalMux
    port map (
            O => \N__40455\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18\
        );

    \I__8611\ : InMux
    port map (
            O => \N__40452\,
            I => \N__40449\
        );

    \I__8610\ : LocalMux
    port map (
            O => \N__40449\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17\
        );

    \I__8609\ : InMux
    port map (
            O => \N__40446\,
            I => \N__40442\
        );

    \I__8608\ : InMux
    port map (
            O => \N__40445\,
            I => \N__40439\
        );

    \I__8607\ : LocalMux
    port map (
            O => \N__40442\,
            I => \N__40434\
        );

    \I__8606\ : LocalMux
    port map (
            O => \N__40439\,
            I => \N__40434\
        );

    \I__8605\ : Span4Mux_h
    port map (
            O => \N__40434\,
            I => \N__40430\
        );

    \I__8604\ : InMux
    port map (
            O => \N__40433\,
            I => \N__40427\
        );

    \I__8603\ : Span4Mux_h
    port map (
            O => \N__40430\,
            I => \N__40424\
        );

    \I__8602\ : LocalMux
    port map (
            O => \N__40427\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\
        );

    \I__8601\ : Odrv4
    port map (
            O => \N__40424\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\
        );

    \I__8600\ : InMux
    port map (
            O => \N__40419\,
            I => \N__40416\
        );

    \I__8599\ : LocalMux
    port map (
            O => \N__40416\,
            I => \N__40411\
        );

    \I__8598\ : InMux
    port map (
            O => \N__40415\,
            I => \N__40408\
        );

    \I__8597\ : InMux
    port map (
            O => \N__40414\,
            I => \N__40405\
        );

    \I__8596\ : Span4Mux_v
    port map (
            O => \N__40411\,
            I => \N__40398\
        );

    \I__8595\ : LocalMux
    port map (
            O => \N__40408\,
            I => \N__40398\
        );

    \I__8594\ : LocalMux
    port map (
            O => \N__40405\,
            I => \N__40398\
        );

    \I__8593\ : Span4Mux_h
    port map (
            O => \N__40398\,
            I => \N__40394\
        );

    \I__8592\ : InMux
    port map (
            O => \N__40397\,
            I => \N__40391\
        );

    \I__8591\ : Odrv4
    port map (
            O => \N__40394\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__8590\ : LocalMux
    port map (
            O => \N__40391\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__8589\ : InMux
    port map (
            O => \N__40386\,
            I => \N__40383\
        );

    \I__8588\ : LocalMux
    port map (
            O => \N__40383\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\
        );

    \I__8587\ : CascadeMux
    port map (
            O => \N__40380\,
            I => \elapsed_time_ns_1_RNISAHF91_0_13_cascade_\
        );

    \I__8586\ : InMux
    port map (
            O => \N__40377\,
            I => \N__40374\
        );

    \I__8585\ : LocalMux
    port map (
            O => \N__40374\,
            I => \N__40371\
        );

    \I__8584\ : Span4Mux_v
    port map (
            O => \N__40371\,
            I => \N__40368\
        );

    \I__8583\ : Odrv4
    port map (
            O => \N__40368\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\
        );

    \I__8582\ : InMux
    port map (
            O => \N__40365\,
            I => \N__40362\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__40362\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9\
        );

    \I__8580\ : InMux
    port map (
            O => \N__40359\,
            I => \N__40356\
        );

    \I__8579\ : LocalMux
    port map (
            O => \N__40356\,
            I => \N__40353\
        );

    \I__8578\ : Span4Mux_v
    port map (
            O => \N__40353\,
            I => \N__40350\
        );

    \I__8577\ : Odrv4
    port map (
            O => \N__40350\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\
        );

    \I__8576\ : InMux
    port map (
            O => \N__40347\,
            I => \N__40344\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__40344\,
            I => \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\
        );

    \I__8574\ : InMux
    port map (
            O => \N__40341\,
            I => \N__40338\
        );

    \I__8573\ : LocalMux
    port map (
            O => \N__40338\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\
        );

    \I__8572\ : InMux
    port map (
            O => \N__40335\,
            I => \N__40332\
        );

    \I__8571\ : LocalMux
    port map (
            O => \N__40332\,
            I => \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\
        );

    \I__8570\ : CascadeMux
    port map (
            O => \N__40329\,
            I => \N__40326\
        );

    \I__8569\ : InMux
    port map (
            O => \N__40326\,
            I => \N__40323\
        );

    \I__8568\ : LocalMux
    port map (
            O => \N__40323\,
            I => \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\
        );

    \I__8567\ : InMux
    port map (
            O => \N__40320\,
            I => \N__40315\
        );

    \I__8566\ : InMux
    port map (
            O => \N__40319\,
            I => \N__40311\
        );

    \I__8565\ : InMux
    port map (
            O => \N__40318\,
            I => \N__40308\
        );

    \I__8564\ : LocalMux
    port map (
            O => \N__40315\,
            I => \N__40305\
        );

    \I__8563\ : InMux
    port map (
            O => \N__40314\,
            I => \N__40302\
        );

    \I__8562\ : LocalMux
    port map (
            O => \N__40311\,
            I => \N__40297\
        );

    \I__8561\ : LocalMux
    port map (
            O => \N__40308\,
            I => \N__40297\
        );

    \I__8560\ : Span4Mux_h
    port map (
            O => \N__40305\,
            I => \N__40294\
        );

    \I__8559\ : LocalMux
    port map (
            O => \N__40302\,
            I => \N__40291\
        );

    \I__8558\ : Span4Mux_h
    port map (
            O => \N__40297\,
            I => \N__40288\
        );

    \I__8557\ : Span4Mux_h
    port map (
            O => \N__40294\,
            I => \N__40285\
        );

    \I__8556\ : Odrv12
    port map (
            O => \N__40291\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__8555\ : Odrv4
    port map (
            O => \N__40288\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__8554\ : Odrv4
    port map (
            O => \N__40285\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__8553\ : CascadeMux
    port map (
            O => \N__40278\,
            I => \N__40275\
        );

    \I__8552\ : InMux
    port map (
            O => \N__40275\,
            I => \N__40272\
        );

    \I__8551\ : LocalMux
    port map (
            O => \N__40272\,
            I => \N__40269\
        );

    \I__8550\ : Span4Mux_h
    port map (
            O => \N__40269\,
            I => \N__40266\
        );

    \I__8549\ : Span4Mux_h
    port map (
            O => \N__40266\,
            I => \N__40263\
        );

    \I__8548\ : Odrv4
    port map (
            O => \N__40263\,
            I => \current_shift_inst.PI_CTRL.integrator_i_29\
        );

    \I__8547\ : InMux
    port map (
            O => \N__40260\,
            I => \N__40257\
        );

    \I__8546\ : LocalMux
    port map (
            O => \N__40257\,
            I => \N__40253\
        );

    \I__8545\ : InMux
    port map (
            O => \N__40256\,
            I => \N__40250\
        );

    \I__8544\ : Span4Mux_v
    port map (
            O => \N__40253\,
            I => \N__40245\
        );

    \I__8543\ : LocalMux
    port map (
            O => \N__40250\,
            I => \N__40245\
        );

    \I__8542\ : Span4Mux_v
    port map (
            O => \N__40245\,
            I => \N__40240\
        );

    \I__8541\ : InMux
    port map (
            O => \N__40244\,
            I => \N__40235\
        );

    \I__8540\ : InMux
    port map (
            O => \N__40243\,
            I => \N__40235\
        );

    \I__8539\ : Odrv4
    port map (
            O => \N__40240\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__40235\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__8537\ : InMux
    port map (
            O => \N__40230\,
            I => \N__40227\
        );

    \I__8536\ : LocalMux
    port map (
            O => \N__40227\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\
        );

    \I__8535\ : InMux
    port map (
            O => \N__40224\,
            I => \N__40219\
        );

    \I__8534\ : InMux
    port map (
            O => \N__40223\,
            I => \N__40216\
        );

    \I__8533\ : InMux
    port map (
            O => \N__40222\,
            I => \N__40213\
        );

    \I__8532\ : LocalMux
    port map (
            O => \N__40219\,
            I => \N__40208\
        );

    \I__8531\ : LocalMux
    port map (
            O => \N__40216\,
            I => \N__40208\
        );

    \I__8530\ : LocalMux
    port map (
            O => \N__40213\,
            I => \N__40205\
        );

    \I__8529\ : Span4Mux_v
    port map (
            O => \N__40208\,
            I => \N__40201\
        );

    \I__8528\ : Span4Mux_h
    port map (
            O => \N__40205\,
            I => \N__40198\
        );

    \I__8527\ : InMux
    port map (
            O => \N__40204\,
            I => \N__40195\
        );

    \I__8526\ : Odrv4
    port map (
            O => \N__40201\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__8525\ : Odrv4
    port map (
            O => \N__40198\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__8524\ : LocalMux
    port map (
            O => \N__40195\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__8523\ : CascadeMux
    port map (
            O => \N__40188\,
            I => \N__40185\
        );

    \I__8522\ : InMux
    port map (
            O => \N__40185\,
            I => \N__40182\
        );

    \I__8521\ : LocalMux
    port map (
            O => \N__40182\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\
        );

    \I__8520\ : CascadeMux
    port map (
            O => \N__40179\,
            I => \N__40176\
        );

    \I__8519\ : InMux
    port map (
            O => \N__40176\,
            I => \N__40173\
        );

    \I__8518\ : LocalMux
    port map (
            O => \N__40173\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\
        );

    \I__8517\ : CascadeMux
    port map (
            O => \N__40170\,
            I => \N__40167\
        );

    \I__8516\ : InMux
    port map (
            O => \N__40167\,
            I => \N__40164\
        );

    \I__8515\ : LocalMux
    port map (
            O => \N__40164\,
            I => \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\
        );

    \I__8514\ : InMux
    port map (
            O => \N__40161\,
            I => \N__40158\
        );

    \I__8513\ : LocalMux
    port map (
            O => \N__40158\,
            I => \N__40155\
        );

    \I__8512\ : Span4Mux_h
    port map (
            O => \N__40155\,
            I => \N__40152\
        );

    \I__8511\ : Odrv4
    port map (
            O => \N__40152\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\
        );

    \I__8510\ : InMux
    port map (
            O => \N__40149\,
            I => \N__40146\
        );

    \I__8509\ : LocalMux
    port map (
            O => \N__40146\,
            I => \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\
        );

    \I__8508\ : CascadeMux
    port map (
            O => \N__40143\,
            I => \N__40140\
        );

    \I__8507\ : InMux
    port map (
            O => \N__40140\,
            I => \N__40137\
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__40137\,
            I => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\
        );

    \I__8505\ : CascadeMux
    port map (
            O => \N__40134\,
            I => \N__40131\
        );

    \I__8504\ : InMux
    port map (
            O => \N__40131\,
            I => \N__40127\
        );

    \I__8503\ : CascadeMux
    port map (
            O => \N__40130\,
            I => \N__40124\
        );

    \I__8502\ : LocalMux
    port map (
            O => \N__40127\,
            I => \N__40120\
        );

    \I__8501\ : InMux
    port map (
            O => \N__40124\,
            I => \N__40117\
        );

    \I__8500\ : InMux
    port map (
            O => \N__40123\,
            I => \N__40114\
        );

    \I__8499\ : Span4Mux_v
    port map (
            O => \N__40120\,
            I => \N__40110\
        );

    \I__8498\ : LocalMux
    port map (
            O => \N__40117\,
            I => \N__40107\
        );

    \I__8497\ : LocalMux
    port map (
            O => \N__40114\,
            I => \N__40104\
        );

    \I__8496\ : InMux
    port map (
            O => \N__40113\,
            I => \N__40101\
        );

    \I__8495\ : Span4Mux_v
    port map (
            O => \N__40110\,
            I => \N__40092\
        );

    \I__8494\ : Span4Mux_v
    port map (
            O => \N__40107\,
            I => \N__40092\
        );

    \I__8493\ : Span4Mux_h
    port map (
            O => \N__40104\,
            I => \N__40092\
        );

    \I__8492\ : LocalMux
    port map (
            O => \N__40101\,
            I => \N__40092\
        );

    \I__8491\ : Odrv4
    port map (
            O => \N__40092\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__8490\ : InMux
    port map (
            O => \N__40089\,
            I => \N__40086\
        );

    \I__8489\ : LocalMux
    port map (
            O => \N__40086\,
            I => \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\
        );

    \I__8488\ : CascadeMux
    port map (
            O => \N__40083\,
            I => \N__40080\
        );

    \I__8487\ : InMux
    port map (
            O => \N__40080\,
            I => \N__40077\
        );

    \I__8486\ : LocalMux
    port map (
            O => \N__40077\,
            I => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\
        );

    \I__8485\ : CascadeMux
    port map (
            O => \N__40074\,
            I => \N__40069\
        );

    \I__8484\ : CascadeMux
    port map (
            O => \N__40073\,
            I => \N__40066\
        );

    \I__8483\ : InMux
    port map (
            O => \N__40072\,
            I => \N__40063\
        );

    \I__8482\ : InMux
    port map (
            O => \N__40069\,
            I => \N__40059\
        );

    \I__8481\ : InMux
    port map (
            O => \N__40066\,
            I => \N__40056\
        );

    \I__8480\ : LocalMux
    port map (
            O => \N__40063\,
            I => \N__40053\
        );

    \I__8479\ : CascadeMux
    port map (
            O => \N__40062\,
            I => \N__40050\
        );

    \I__8478\ : LocalMux
    port map (
            O => \N__40059\,
            I => \N__40046\
        );

    \I__8477\ : LocalMux
    port map (
            O => \N__40056\,
            I => \N__40043\
        );

    \I__8476\ : Span4Mux_h
    port map (
            O => \N__40053\,
            I => \N__40040\
        );

    \I__8475\ : InMux
    port map (
            O => \N__40050\,
            I => \N__40035\
        );

    \I__8474\ : InMux
    port map (
            O => \N__40049\,
            I => \N__40035\
        );

    \I__8473\ : Span4Mux_h
    port map (
            O => \N__40046\,
            I => \N__40030\
        );

    \I__8472\ : Span4Mux_v
    port map (
            O => \N__40043\,
            I => \N__40030\
        );

    \I__8471\ : Span4Mux_h
    port map (
            O => \N__40040\,
            I => \N__40027\
        );

    \I__8470\ : LocalMux
    port map (
            O => \N__40035\,
            I => \N__40024\
        );

    \I__8469\ : Odrv4
    port map (
            O => \N__40030\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__8468\ : Odrv4
    port map (
            O => \N__40027\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__8467\ : Odrv4
    port map (
            O => \N__40024\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__8466\ : InMux
    port map (
            O => \N__40017\,
            I => \N__40014\
        );

    \I__8465\ : LocalMux
    port map (
            O => \N__40014\,
            I => \N__40011\
        );

    \I__8464\ : Span4Mux_v
    port map (
            O => \N__40011\,
            I => \N__40008\
        );

    \I__8463\ : Span4Mux_h
    port map (
            O => \N__40008\,
            I => \N__40005\
        );

    \I__8462\ : Odrv4
    port map (
            O => \N__40005\,
            I => \current_shift_inst.PI_CTRL.integrator_i_26\
        );

    \I__8461\ : CascadeMux
    port map (
            O => \N__40002\,
            I => \N__39999\
        );

    \I__8460\ : InMux
    port map (
            O => \N__39999\,
            I => \N__39996\
        );

    \I__8459\ : LocalMux
    port map (
            O => \N__39996\,
            I => \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\
        );

    \I__8458\ : InMux
    port map (
            O => \N__39993\,
            I => \N__39990\
        );

    \I__8457\ : LocalMux
    port map (
            O => \N__39990\,
            I => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\
        );

    \I__8456\ : InMux
    port map (
            O => \N__39987\,
            I => \N__39984\
        );

    \I__8455\ : LocalMux
    port map (
            O => \N__39984\,
            I => \N__39981\
        );

    \I__8454\ : Span4Mux_v
    port map (
            O => \N__39981\,
            I => \N__39977\
        );

    \I__8453\ : InMux
    port map (
            O => \N__39980\,
            I => \N__39974\
        );

    \I__8452\ : Sp12to4
    port map (
            O => \N__39977\,
            I => \N__39968\
        );

    \I__8451\ : LocalMux
    port map (
            O => \N__39974\,
            I => \N__39968\
        );

    \I__8450\ : InMux
    port map (
            O => \N__39973\,
            I => \N__39965\
        );

    \I__8449\ : Odrv12
    port map (
            O => \N__39968\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__39965\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__8447\ : CascadeMux
    port map (
            O => \N__39960\,
            I => \N__39957\
        );

    \I__8446\ : InMux
    port map (
            O => \N__39957\,
            I => \N__39954\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__39954\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\
        );

    \I__8444\ : CascadeMux
    port map (
            O => \N__39951\,
            I => \N__39948\
        );

    \I__8443\ : InMux
    port map (
            O => \N__39948\,
            I => \N__39942\
        );

    \I__8442\ : InMux
    port map (
            O => \N__39947\,
            I => \N__39942\
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__39942\,
            I => \N__39937\
        );

    \I__8440\ : InMux
    port map (
            O => \N__39941\,
            I => \N__39932\
        );

    \I__8439\ : InMux
    port map (
            O => \N__39940\,
            I => \N__39932\
        );

    \I__8438\ : Span4Mux_v
    port map (
            O => \N__39937\,
            I => \N__39927\
        );

    \I__8437\ : LocalMux
    port map (
            O => \N__39932\,
            I => \N__39927\
        );

    \I__8436\ : Odrv4
    port map (
            O => \N__39927\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__8435\ : CascadeMux
    port map (
            O => \N__39924\,
            I => \N__39921\
        );

    \I__8434\ : InMux
    port map (
            O => \N__39921\,
            I => \N__39918\
        );

    \I__8433\ : LocalMux
    port map (
            O => \N__39918\,
            I => \current_shift_inst.un38_control_input_cry_0_s0_sf\
        );

    \I__8432\ : InMux
    port map (
            O => \N__39915\,
            I => \N__39912\
        );

    \I__8431\ : LocalMux
    port map (
            O => \N__39912\,
            I => \current_shift_inst.un4_control_input1_1\
        );

    \I__8430\ : CascadeMux
    port map (
            O => \N__39909\,
            I => \current_shift_inst.un4_control_input1_1_cascade_\
        );

    \I__8429\ : CascadeMux
    port map (
            O => \N__39906\,
            I => \N__39903\
        );

    \I__8428\ : InMux
    port map (
            O => \N__39903\,
            I => \N__39900\
        );

    \I__8427\ : LocalMux
    port map (
            O => \N__39900\,
            I => \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\
        );

    \I__8426\ : CascadeMux
    port map (
            O => \N__39897\,
            I => \N__39894\
        );

    \I__8425\ : InMux
    port map (
            O => \N__39894\,
            I => \N__39891\
        );

    \I__8424\ : LocalMux
    port map (
            O => \N__39891\,
            I => \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\
        );

    \I__8423\ : InMux
    port map (
            O => \N__39888\,
            I => \N__39885\
        );

    \I__8422\ : LocalMux
    port map (
            O => \N__39885\,
            I => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\
        );

    \I__8421\ : CascadeMux
    port map (
            O => \N__39882\,
            I => \N__39879\
        );

    \I__8420\ : InMux
    port map (
            O => \N__39879\,
            I => \N__39876\
        );

    \I__8419\ : LocalMux
    port map (
            O => \N__39876\,
            I => \N__39873\
        );

    \I__8418\ : Span4Mux_h
    port map (
            O => \N__39873\,
            I => \N__39870\
        );

    \I__8417\ : Span4Mux_v
    port map (
            O => \N__39870\,
            I => \N__39867\
        );

    \I__8416\ : Odrv4
    port map (
            O => \N__39867\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\
        );

    \I__8415\ : CascadeMux
    port map (
            O => \N__39864\,
            I => \N__39860\
        );

    \I__8414\ : InMux
    port map (
            O => \N__39863\,
            I => \N__39852\
        );

    \I__8413\ : InMux
    port map (
            O => \N__39860\,
            I => \N__39852\
        );

    \I__8412\ : InMux
    port map (
            O => \N__39859\,
            I => \N__39852\
        );

    \I__8411\ : LocalMux
    port map (
            O => \N__39852\,
            I => \N__39848\
        );

    \I__8410\ : InMux
    port map (
            O => \N__39851\,
            I => \N__39845\
        );

    \I__8409\ : Odrv4
    port map (
            O => \N__39848\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__8408\ : LocalMux
    port map (
            O => \N__39845\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__8407\ : CascadeMux
    port map (
            O => \N__39840\,
            I => \N__39837\
        );

    \I__8406\ : InMux
    port map (
            O => \N__39837\,
            I => \N__39834\
        );

    \I__8405\ : LocalMux
    port map (
            O => \N__39834\,
            I => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\
        );

    \I__8404\ : InMux
    port map (
            O => \N__39831\,
            I => \N__39828\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__39828\,
            I => \N__39825\
        );

    \I__8402\ : Span4Mux_v
    port map (
            O => \N__39825\,
            I => \N__39822\
        );

    \I__8401\ : Odrv4
    port map (
            O => \N__39822\,
            I => \current_shift_inst.un38_control_input_axb_31_s0\
        );

    \I__8400\ : InMux
    port map (
            O => \N__39819\,
            I => \N__39816\
        );

    \I__8399\ : LocalMux
    port map (
            O => \N__39816\,
            I => \N__39813\
        );

    \I__8398\ : Span4Mux_v
    port map (
            O => \N__39813\,
            I => \N__39810\
        );

    \I__8397\ : Odrv4
    port map (
            O => \N__39810\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\
        );

    \I__8396\ : CascadeMux
    port map (
            O => \N__39807\,
            I => \N__39803\
        );

    \I__8395\ : InMux
    port map (
            O => \N__39806\,
            I => \N__39795\
        );

    \I__8394\ : InMux
    port map (
            O => \N__39803\,
            I => \N__39795\
        );

    \I__8393\ : InMux
    port map (
            O => \N__39802\,
            I => \N__39795\
        );

    \I__8392\ : LocalMux
    port map (
            O => \N__39795\,
            I => \N__39792\
        );

    \I__8391\ : Span4Mux_h
    port map (
            O => \N__39792\,
            I => \N__39788\
        );

    \I__8390\ : InMux
    port map (
            O => \N__39791\,
            I => \N__39785\
        );

    \I__8389\ : Odrv4
    port map (
            O => \N__39788\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__8388\ : LocalMux
    port map (
            O => \N__39785\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__8387\ : InMux
    port map (
            O => \N__39780\,
            I => \N__39777\
        );

    \I__8386\ : LocalMux
    port map (
            O => \N__39777\,
            I => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\
        );

    \I__8385\ : CascadeMux
    port map (
            O => \N__39774\,
            I => \N__39771\
        );

    \I__8384\ : InMux
    port map (
            O => \N__39771\,
            I => \N__39768\
        );

    \I__8383\ : LocalMux
    port map (
            O => \N__39768\,
            I => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\
        );

    \I__8382\ : CascadeMux
    port map (
            O => \N__39765\,
            I => \N__39762\
        );

    \I__8381\ : InMux
    port map (
            O => \N__39762\,
            I => \N__39759\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__39759\,
            I => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\
        );

    \I__8379\ : CascadeMux
    port map (
            O => \N__39756\,
            I => \N__39753\
        );

    \I__8378\ : InMux
    port map (
            O => \N__39753\,
            I => \N__39750\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__39750\,
            I => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\
        );

    \I__8376\ : CascadeMux
    port map (
            O => \N__39747\,
            I => \N__39744\
        );

    \I__8375\ : InMux
    port map (
            O => \N__39744\,
            I => \N__39741\
        );

    \I__8374\ : LocalMux
    port map (
            O => \N__39741\,
            I => \N__39738\
        );

    \I__8373\ : Span4Mux_v
    port map (
            O => \N__39738\,
            I => \N__39735\
        );

    \I__8372\ : Odrv4
    port map (
            O => \N__39735\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\
        );

    \I__8371\ : CascadeMux
    port map (
            O => \N__39732\,
            I => \N__39729\
        );

    \I__8370\ : InMux
    port map (
            O => \N__39729\,
            I => \N__39726\
        );

    \I__8369\ : LocalMux
    port map (
            O => \N__39726\,
            I => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\
        );

    \I__8368\ : CascadeMux
    port map (
            O => \N__39723\,
            I => \N__39720\
        );

    \I__8367\ : InMux
    port map (
            O => \N__39720\,
            I => \N__39717\
        );

    \I__8366\ : LocalMux
    port map (
            O => \N__39717\,
            I => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\
        );

    \I__8365\ : InMux
    port map (
            O => \N__39714\,
            I => \N__39711\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__39711\,
            I => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\
        );

    \I__8363\ : InMux
    port map (
            O => \N__39708\,
            I => \N__39705\
        );

    \I__8362\ : LocalMux
    port map (
            O => \N__39705\,
            I => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\
        );

    \I__8361\ : InMux
    port map (
            O => \N__39702\,
            I => \N__39699\
        );

    \I__8360\ : LocalMux
    port map (
            O => \N__39699\,
            I => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\
        );

    \I__8359\ : InMux
    port map (
            O => \N__39696\,
            I => \N__39693\
        );

    \I__8358\ : LocalMux
    port map (
            O => \N__39693\,
            I => \N__39690\
        );

    \I__8357\ : Span12Mux_h
    port map (
            O => \N__39690\,
            I => \N__39687\
        );

    \I__8356\ : Odrv12
    port map (
            O => \N__39687\,
            I => \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\
        );

    \I__8355\ : CascadeMux
    port map (
            O => \N__39684\,
            I => \N__39678\
        );

    \I__8354\ : InMux
    port map (
            O => \N__39683\,
            I => \N__39673\
        );

    \I__8353\ : InMux
    port map (
            O => \N__39682\,
            I => \N__39673\
        );

    \I__8352\ : InMux
    port map (
            O => \N__39681\,
            I => \N__39668\
        );

    \I__8351\ : InMux
    port map (
            O => \N__39678\,
            I => \N__39668\
        );

    \I__8350\ : LocalMux
    port map (
            O => \N__39673\,
            I => \N__39665\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__39668\,
            I => \N__39662\
        );

    \I__8348\ : Span4Mux_v
    port map (
            O => \N__39665\,
            I => \N__39659\
        );

    \I__8347\ : Odrv12
    port map (
            O => \N__39662\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__8346\ : Odrv4
    port map (
            O => \N__39659\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__8345\ : CascadeMux
    port map (
            O => \N__39654\,
            I => \N__39651\
        );

    \I__8344\ : InMux
    port map (
            O => \N__39651\,
            I => \N__39648\
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__39648\,
            I => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\
        );

    \I__8342\ : CascadeMux
    port map (
            O => \N__39645\,
            I => \N__39642\
        );

    \I__8341\ : InMux
    port map (
            O => \N__39642\,
            I => \N__39639\
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__39639\,
            I => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\
        );

    \I__8339\ : InMux
    port map (
            O => \N__39636\,
            I => \N__39633\
        );

    \I__8338\ : LocalMux
    port map (
            O => \N__39633\,
            I => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\
        );

    \I__8337\ : InMux
    port map (
            O => \N__39630\,
            I => \N__39627\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__39627\,
            I => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\
        );

    \I__8335\ : CascadeMux
    port map (
            O => \N__39624\,
            I => \N__39621\
        );

    \I__8334\ : InMux
    port map (
            O => \N__39621\,
            I => \N__39618\
        );

    \I__8333\ : LocalMux
    port map (
            O => \N__39618\,
            I => \N__39615\
        );

    \I__8332\ : Odrv4
    port map (
            O => \N__39615\,
            I => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\
        );

    \I__8331\ : InMux
    port map (
            O => \N__39612\,
            I => \N__39608\
        );

    \I__8330\ : InMux
    port map (
            O => \N__39611\,
            I => \N__39605\
        );

    \I__8329\ : LocalMux
    port map (
            O => \N__39608\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__8328\ : LocalMux
    port map (
            O => \N__39605\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__8327\ : InMux
    port map (
            O => \N__39600\,
            I => \N__39596\
        );

    \I__8326\ : InMux
    port map (
            O => \N__39599\,
            I => \N__39593\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__39596\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__39593\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__8323\ : InMux
    port map (
            O => \N__39588\,
            I => \N__39585\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__39585\,
            I => \N__39582\
        );

    \I__8321\ : Odrv4
    port map (
            O => \N__39582\,
            I => \phase_controller_inst1.stoper_tr.un4_running_df26\
        );

    \I__8320\ : InMux
    port map (
            O => \N__39579\,
            I => \N__39574\
        );

    \I__8319\ : InMux
    port map (
            O => \N__39578\,
            I => \N__39571\
        );

    \I__8318\ : InMux
    port map (
            O => \N__39577\,
            I => \N__39568\
        );

    \I__8317\ : LocalMux
    port map (
            O => \N__39574\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__39571\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__8315\ : LocalMux
    port map (
            O => \N__39568\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__8314\ : InMux
    port map (
            O => \N__39561\,
            I => \N__39556\
        );

    \I__8313\ : InMux
    port map (
            O => \N__39560\,
            I => \N__39553\
        );

    \I__8312\ : InMux
    port map (
            O => \N__39559\,
            I => \N__39550\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__39556\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__8310\ : LocalMux
    port map (
            O => \N__39553\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__8309\ : LocalMux
    port map (
            O => \N__39550\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__8308\ : CascadeMux
    port map (
            O => \N__39543\,
            I => \N__39540\
        );

    \I__8307\ : InMux
    port map (
            O => \N__39540\,
            I => \N__39537\
        );

    \I__8306\ : LocalMux
    port map (
            O => \N__39537\,
            I => \N__39534\
        );

    \I__8305\ : Odrv4
    port map (
            O => \N__39534\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt18\
        );

    \I__8304\ : InMux
    port map (
            O => \N__39531\,
            I => \N__39528\
        );

    \I__8303\ : LocalMux
    port map (
            O => \N__39528\,
            I => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\
        );

    \I__8302\ : InMux
    port map (
            O => \N__39525\,
            I => \N__39520\
        );

    \I__8301\ : InMux
    port map (
            O => \N__39524\,
            I => \N__39515\
        );

    \I__8300\ : InMux
    port map (
            O => \N__39523\,
            I => \N__39515\
        );

    \I__8299\ : LocalMux
    port map (
            O => \N__39520\,
            I => \N__39511\
        );

    \I__8298\ : LocalMux
    port map (
            O => \N__39515\,
            I => \N__39508\
        );

    \I__8297\ : InMux
    port map (
            O => \N__39514\,
            I => \N__39505\
        );

    \I__8296\ : Span4Mux_v
    port map (
            O => \N__39511\,
            I => \N__39498\
        );

    \I__8295\ : Span4Mux_h
    port map (
            O => \N__39508\,
            I => \N__39498\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__39505\,
            I => \N__39498\
        );

    \I__8293\ : Odrv4
    port map (
            O => \N__39498\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__8292\ : InMux
    port map (
            O => \N__39495\,
            I => \N__39492\
        );

    \I__8291\ : LocalMux
    port map (
            O => \N__39492\,
            I => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\
        );

    \I__8290\ : CascadeMux
    port map (
            O => \N__39489\,
            I => \N__39486\
        );

    \I__8289\ : InMux
    port map (
            O => \N__39486\,
            I => \N__39483\
        );

    \I__8288\ : LocalMux
    port map (
            O => \N__39483\,
            I => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\
        );

    \I__8287\ : CascadeMux
    port map (
            O => \N__39480\,
            I => \N__39477\
        );

    \I__8286\ : InMux
    port map (
            O => \N__39477\,
            I => \N__39474\
        );

    \I__8285\ : LocalMux
    port map (
            O => \N__39474\,
            I => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\
        );

    \I__8284\ : InMux
    port map (
            O => \N__39471\,
            I => \N__39468\
        );

    \I__8283\ : LocalMux
    port map (
            O => \N__39468\,
            I => \N__39465\
        );

    \I__8282\ : Odrv4
    port map (
            O => \N__39465\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO\
        );

    \I__8281\ : InMux
    port map (
            O => \N__39462\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_28\
        );

    \I__8280\ : InMux
    port map (
            O => \N__39459\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30\
        );

    \I__8279\ : InMux
    port map (
            O => \N__39456\,
            I => \N__39452\
        );

    \I__8278\ : InMux
    port map (
            O => \N__39455\,
            I => \N__39449\
        );

    \I__8277\ : LocalMux
    port map (
            O => \N__39452\,
            I => \N__39446\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__39449\,
            I => \N__39443\
        );

    \I__8275\ : Span4Mux_h
    port map (
            O => \N__39446\,
            I => \N__39440\
        );

    \I__8274\ : Odrv4
    port map (
            O => \N__39443\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__8273\ : Odrv4
    port map (
            O => \N__39440\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__8272\ : InMux
    port map (
            O => \N__39435\,
            I => \N__39432\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__39432\,
            I => \N__39429\
        );

    \I__8270\ : Odrv4
    port map (
            O => \N__39429\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt16\
        );

    \I__8269\ : InMux
    port map (
            O => \N__39426\,
            I => \N__39419\
        );

    \I__8268\ : InMux
    port map (
            O => \N__39425\,
            I => \N__39419\
        );

    \I__8267\ : InMux
    port map (
            O => \N__39424\,
            I => \N__39416\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__39419\,
            I => \N__39413\
        );

    \I__8265\ : LocalMux
    port map (
            O => \N__39416\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__8264\ : Odrv4
    port map (
            O => \N__39413\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__8263\ : InMux
    port map (
            O => \N__39408\,
            I => \N__39403\
        );

    \I__8262\ : InMux
    port map (
            O => \N__39407\,
            I => \N__39398\
        );

    \I__8261\ : InMux
    port map (
            O => \N__39406\,
            I => \N__39398\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__39403\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__8259\ : LocalMux
    port map (
            O => \N__39398\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__8258\ : CascadeMux
    port map (
            O => \N__39393\,
            I => \N__39390\
        );

    \I__8257\ : InMux
    port map (
            O => \N__39390\,
            I => \N__39387\
        );

    \I__8256\ : LocalMux
    port map (
            O => \N__39387\,
            I => \N__39384\
        );

    \I__8255\ : Span4Mux_h
    port map (
            O => \N__39384\,
            I => \N__39381\
        );

    \I__8254\ : Odrv4
    port map (
            O => \N__39381\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\
        );

    \I__8253\ : CascadeMux
    port map (
            O => \N__39378\,
            I => \N__39375\
        );

    \I__8252\ : InMux
    port map (
            O => \N__39375\,
            I => \N__39369\
        );

    \I__8251\ : InMux
    port map (
            O => \N__39374\,
            I => \N__39369\
        );

    \I__8250\ : LocalMux
    port map (
            O => \N__39369\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__8249\ : InMux
    port map (
            O => \N__39366\,
            I => \N__39363\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__39363\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\
        );

    \I__8247\ : InMux
    port map (
            O => \N__39360\,
            I => \N__39355\
        );

    \I__8246\ : InMux
    port map (
            O => \N__39359\,
            I => \N__39351\
        );

    \I__8245\ : InMux
    port map (
            O => \N__39358\,
            I => \N__39348\
        );

    \I__8244\ : LocalMux
    port map (
            O => \N__39355\,
            I => \N__39345\
        );

    \I__8243\ : InMux
    port map (
            O => \N__39354\,
            I => \N__39342\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__39351\,
            I => \N__39339\
        );

    \I__8241\ : LocalMux
    port map (
            O => \N__39348\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__8240\ : Odrv4
    port map (
            O => \N__39345\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__8239\ : LocalMux
    port map (
            O => \N__39342\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__8238\ : Odrv12
    port map (
            O => \N__39339\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__8237\ : CascadeMux
    port map (
            O => \N__39330\,
            I => \N__39327\
        );

    \I__8236\ : InMux
    port map (
            O => \N__39327\,
            I => \N__39324\
        );

    \I__8235\ : LocalMux
    port map (
            O => \N__39324\,
            I => \N__39319\
        );

    \I__8234\ : InMux
    port map (
            O => \N__39323\,
            I => \N__39316\
        );

    \I__8233\ : InMux
    port map (
            O => \N__39322\,
            I => \N__39313\
        );

    \I__8232\ : Span4Mux_h
    port map (
            O => \N__39319\,
            I => \N__39310\
        );

    \I__8231\ : LocalMux
    port map (
            O => \N__39316\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__8230\ : LocalMux
    port map (
            O => \N__39313\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__8229\ : Odrv4
    port map (
            O => \N__39310\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__8228\ : CascadeMux
    port map (
            O => \N__39303\,
            I => \N__39300\
        );

    \I__8227\ : InMux
    port map (
            O => \N__39300\,
            I => \N__39297\
        );

    \I__8226\ : LocalMux
    port map (
            O => \N__39297\,
            I => \N__39294\
        );

    \I__8225\ : Odrv4
    port map (
            O => \N__39294\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30\
        );

    \I__8224\ : InMux
    port map (
            O => \N__39291\,
            I => \N__39287\
        );

    \I__8223\ : InMux
    port map (
            O => \N__39290\,
            I => \N__39284\
        );

    \I__8222\ : LocalMux
    port map (
            O => \N__39287\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__8221\ : LocalMux
    port map (
            O => \N__39284\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__8220\ : InMux
    port map (
            O => \N__39279\,
            I => \N__39275\
        );

    \I__8219\ : InMux
    port map (
            O => \N__39278\,
            I => \N__39272\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__39275\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__8217\ : LocalMux
    port map (
            O => \N__39272\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__8216\ : InMux
    port map (
            O => \N__39267\,
            I => \N__39264\
        );

    \I__8215\ : LocalMux
    port map (
            O => \N__39264\,
            I => \N__39261\
        );

    \I__8214\ : Odrv12
    port map (
            O => \N__39261\,
            I => \phase_controller_inst1.stoper_tr.un4_running_df28\
        );

    \I__8213\ : InMux
    port map (
            O => \N__39258\,
            I => \N__39255\
        );

    \I__8212\ : LocalMux
    port map (
            O => \N__39255\,
            I => \N__39252\
        );

    \I__8211\ : Odrv4
    port map (
            O => \N__39252\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\
        );

    \I__8210\ : InMux
    port map (
            O => \N__39249\,
            I => \N__39245\
        );

    \I__8209\ : InMux
    port map (
            O => \N__39248\,
            I => \N__39242\
        );

    \I__8208\ : LocalMux
    port map (
            O => \N__39245\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__8207\ : LocalMux
    port map (
            O => \N__39242\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__8206\ : CascadeMux
    port map (
            O => \N__39237\,
            I => \N__39234\
        );

    \I__8205\ : InMux
    port map (
            O => \N__39234\,
            I => \N__39231\
        );

    \I__8204\ : LocalMux
    port map (
            O => \N__39231\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__8203\ : CascadeMux
    port map (
            O => \N__39228\,
            I => \N__39225\
        );

    \I__8202\ : InMux
    port map (
            O => \N__39225\,
            I => \N__39222\
        );

    \I__8201\ : LocalMux
    port map (
            O => \N__39222\,
            I => \N__39219\
        );

    \I__8200\ : Odrv12
    port map (
            O => \N__39219\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\
        );

    \I__8199\ : InMux
    port map (
            O => \N__39216\,
            I => \N__39212\
        );

    \I__8198\ : InMux
    port map (
            O => \N__39215\,
            I => \N__39209\
        );

    \I__8197\ : LocalMux
    port map (
            O => \N__39212\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__39209\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__8195\ : InMux
    port map (
            O => \N__39204\,
            I => \N__39201\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__39201\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__8193\ : InMux
    port map (
            O => \N__39198\,
            I => \N__39195\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__39195\,
            I => \N__39192\
        );

    \I__8191\ : Odrv4
    port map (
            O => \N__39192\,
            I => \phase_controller_inst1.stoper_tr.un4_running_df20\
        );

    \I__8190\ : InMux
    port map (
            O => \N__39189\,
            I => \N__39186\
        );

    \I__8189\ : LocalMux
    port map (
            O => \N__39186\,
            I => \N__39183\
        );

    \I__8188\ : Span4Mux_v
    port map (
            O => \N__39183\,
            I => \N__39180\
        );

    \I__8187\ : Odrv4
    port map (
            O => \N__39180\,
            I => \phase_controller_inst1.stoper_tr.un4_running_df22\
        );

    \I__8186\ : InMux
    port map (
            O => \N__39177\,
            I => \N__39174\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__39174\,
            I => \N__39171\
        );

    \I__8184\ : Odrv4
    port map (
            O => \N__39171\,
            I => \phase_controller_inst1.stoper_tr.un4_running_df24\
        );

    \I__8183\ : InMux
    port map (
            O => \N__39168\,
            I => \N__39164\
        );

    \I__8182\ : InMux
    port map (
            O => \N__39167\,
            I => \N__39161\
        );

    \I__8181\ : LocalMux
    port map (
            O => \N__39164\,
            I => \N__39158\
        );

    \I__8180\ : LocalMux
    port map (
            O => \N__39161\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__8179\ : Odrv4
    port map (
            O => \N__39158\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__8178\ : CascadeMux
    port map (
            O => \N__39153\,
            I => \N__39150\
        );

    \I__8177\ : InMux
    port map (
            O => \N__39150\,
            I => \N__39147\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__39147\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__8175\ : CascadeMux
    port map (
            O => \N__39144\,
            I => \N__39141\
        );

    \I__8174\ : InMux
    port map (
            O => \N__39141\,
            I => \N__39138\
        );

    \I__8173\ : LocalMux
    port map (
            O => \N__39138\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\
        );

    \I__8172\ : InMux
    port map (
            O => \N__39135\,
            I => \N__39131\
        );

    \I__8171\ : InMux
    port map (
            O => \N__39134\,
            I => \N__39128\
        );

    \I__8170\ : LocalMux
    port map (
            O => \N__39131\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__8169\ : LocalMux
    port map (
            O => \N__39128\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__8168\ : InMux
    port map (
            O => \N__39123\,
            I => \N__39120\
        );

    \I__8167\ : LocalMux
    port map (
            O => \N__39120\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__8166\ : InMux
    port map (
            O => \N__39117\,
            I => \N__39113\
        );

    \I__8165\ : InMux
    port map (
            O => \N__39116\,
            I => \N__39110\
        );

    \I__8164\ : LocalMux
    port map (
            O => \N__39113\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__8163\ : LocalMux
    port map (
            O => \N__39110\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__8162\ : CascadeMux
    port map (
            O => \N__39105\,
            I => \N__39102\
        );

    \I__8161\ : InMux
    port map (
            O => \N__39102\,
            I => \N__39099\
        );

    \I__8160\ : LocalMux
    port map (
            O => \N__39099\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\
        );

    \I__8159\ : InMux
    port map (
            O => \N__39096\,
            I => \N__39093\
        );

    \I__8158\ : LocalMux
    port map (
            O => \N__39093\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__8157\ : InMux
    port map (
            O => \N__39090\,
            I => \N__39086\
        );

    \I__8156\ : InMux
    port map (
            O => \N__39089\,
            I => \N__39083\
        );

    \I__8155\ : LocalMux
    port map (
            O => \N__39086\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__39083\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__8153\ : CascadeMux
    port map (
            O => \N__39078\,
            I => \N__39075\
        );

    \I__8152\ : InMux
    port map (
            O => \N__39075\,
            I => \N__39072\
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__39072\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__8150\ : InMux
    port map (
            O => \N__39069\,
            I => \N__39065\
        );

    \I__8149\ : InMux
    port map (
            O => \N__39068\,
            I => \N__39062\
        );

    \I__8148\ : LocalMux
    port map (
            O => \N__39065\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__8147\ : LocalMux
    port map (
            O => \N__39062\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__8146\ : InMux
    port map (
            O => \N__39057\,
            I => \N__39054\
        );

    \I__8145\ : LocalMux
    port map (
            O => \N__39054\,
            I => \N__39051\
        );

    \I__8144\ : Span4Mux_h
    port map (
            O => \N__39051\,
            I => \N__39048\
        );

    \I__8143\ : Odrv4
    port map (
            O => \N__39048\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\
        );

    \I__8142\ : CascadeMux
    port map (
            O => \N__39045\,
            I => \N__39042\
        );

    \I__8141\ : InMux
    port map (
            O => \N__39042\,
            I => \N__39039\
        );

    \I__8140\ : LocalMux
    port map (
            O => \N__39039\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__8139\ : InMux
    port map (
            O => \N__39036\,
            I => \N__39033\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__39033\,
            I => \N__39030\
        );

    \I__8137\ : Span4Mux_v
    port map (
            O => \N__39030\,
            I => \N__39027\
        );

    \I__8136\ : Span4Mux_v
    port map (
            O => \N__39027\,
            I => \N__39024\
        );

    \I__8135\ : Odrv4
    port map (
            O => \N__39024\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\
        );

    \I__8134\ : InMux
    port map (
            O => \N__39021\,
            I => \N__39017\
        );

    \I__8133\ : InMux
    port map (
            O => \N__39020\,
            I => \N__39014\
        );

    \I__8132\ : LocalMux
    port map (
            O => \N__39017\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__39014\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__8130\ : CascadeMux
    port map (
            O => \N__39009\,
            I => \N__39006\
        );

    \I__8129\ : InMux
    port map (
            O => \N__39006\,
            I => \N__39003\
        );

    \I__8128\ : LocalMux
    port map (
            O => \N__39003\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__8127\ : InMux
    port map (
            O => \N__39000\,
            I => \N__38996\
        );

    \I__8126\ : InMux
    port map (
            O => \N__38999\,
            I => \N__38993\
        );

    \I__8125\ : LocalMux
    port map (
            O => \N__38996\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__38993\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__8123\ : CascadeMux
    port map (
            O => \N__38988\,
            I => \N__38985\
        );

    \I__8122\ : InMux
    port map (
            O => \N__38985\,
            I => \N__38982\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__38982\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__8120\ : InMux
    port map (
            O => \N__38979\,
            I => \N__38975\
        );

    \I__8119\ : InMux
    port map (
            O => \N__38978\,
            I => \N__38972\
        );

    \I__8118\ : LocalMux
    port map (
            O => \N__38975\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__8117\ : LocalMux
    port map (
            O => \N__38972\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__8116\ : CascadeMux
    port map (
            O => \N__38967\,
            I => \N__38964\
        );

    \I__8115\ : InMux
    port map (
            O => \N__38964\,
            I => \N__38961\
        );

    \I__8114\ : LocalMux
    port map (
            O => \N__38961\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__8113\ : CascadeMux
    port map (
            O => \N__38958\,
            I => \N__38954\
        );

    \I__8112\ : CascadeMux
    port map (
            O => \N__38957\,
            I => \N__38951\
        );

    \I__8111\ : InMux
    port map (
            O => \N__38954\,
            I => \N__38948\
        );

    \I__8110\ : InMux
    port map (
            O => \N__38951\,
            I => \N__38944\
        );

    \I__8109\ : LocalMux
    port map (
            O => \N__38948\,
            I => \N__38941\
        );

    \I__8108\ : InMux
    port map (
            O => \N__38947\,
            I => \N__38938\
        );

    \I__8107\ : LocalMux
    port map (
            O => \N__38944\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8106\ : Odrv4
    port map (
            O => \N__38941\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8105\ : LocalMux
    port map (
            O => \N__38938\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8104\ : CascadeMux
    port map (
            O => \N__38931\,
            I => \N__38928\
        );

    \I__8103\ : InMux
    port map (
            O => \N__38928\,
            I => \N__38925\
        );

    \I__8102\ : LocalMux
    port map (
            O => \N__38925\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__8101\ : InMux
    port map (
            O => \N__38922\,
            I => \N__38918\
        );

    \I__8100\ : InMux
    port map (
            O => \N__38921\,
            I => \N__38915\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__38918\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__8098\ : LocalMux
    port map (
            O => \N__38915\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__8097\ : CascadeMux
    port map (
            O => \N__38910\,
            I => \N__38907\
        );

    \I__8096\ : InMux
    port map (
            O => \N__38907\,
            I => \N__38904\
        );

    \I__8095\ : LocalMux
    port map (
            O => \N__38904\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__8094\ : InMux
    port map (
            O => \N__38901\,
            I => \N__38897\
        );

    \I__8093\ : InMux
    port map (
            O => \N__38900\,
            I => \N__38894\
        );

    \I__8092\ : LocalMux
    port map (
            O => \N__38897\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__38894\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__8090\ : CascadeMux
    port map (
            O => \N__38889\,
            I => \N__38886\
        );

    \I__8089\ : InMux
    port map (
            O => \N__38886\,
            I => \N__38883\
        );

    \I__8088\ : LocalMux
    port map (
            O => \N__38883\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__8087\ : InMux
    port map (
            O => \N__38880\,
            I => \N__38876\
        );

    \I__8086\ : InMux
    port map (
            O => \N__38879\,
            I => \N__38873\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__38876\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__8084\ : LocalMux
    port map (
            O => \N__38873\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__8083\ : CascadeMux
    port map (
            O => \N__38868\,
            I => \N__38865\
        );

    \I__8082\ : InMux
    port map (
            O => \N__38865\,
            I => \N__38862\
        );

    \I__8081\ : LocalMux
    port map (
            O => \N__38862\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__8080\ : InMux
    port map (
            O => \N__38859\,
            I => \N__38855\
        );

    \I__8079\ : InMux
    port map (
            O => \N__38858\,
            I => \N__38852\
        );

    \I__8078\ : LocalMux
    port map (
            O => \N__38855\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__8077\ : LocalMux
    port map (
            O => \N__38852\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__8076\ : InMux
    port map (
            O => \N__38847\,
            I => \N__38844\
        );

    \I__8075\ : LocalMux
    port map (
            O => \N__38844\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\
        );

    \I__8074\ : CascadeMux
    port map (
            O => \N__38841\,
            I => \N__38838\
        );

    \I__8073\ : InMux
    port map (
            O => \N__38838\,
            I => \N__38835\
        );

    \I__8072\ : LocalMux
    port map (
            O => \N__38835\,
            I => \N__38832\
        );

    \I__8071\ : Odrv4
    port map (
            O => \N__38832\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__8070\ : InMux
    port map (
            O => \N__38829\,
            I => \N__38826\
        );

    \I__8069\ : LocalMux
    port map (
            O => \N__38826\,
            I => \N__38823\
        );

    \I__8068\ : Span4Mux_h
    port map (
            O => \N__38823\,
            I => \N__38820\
        );

    \I__8067\ : Span4Mux_h
    port map (
            O => \N__38820\,
            I => \N__38817\
        );

    \I__8066\ : Odrv4
    port map (
            O => \N__38817\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\
        );

    \I__8065\ : InMux
    port map (
            O => \N__38814\,
            I => \N__38807\
        );

    \I__8064\ : InMux
    port map (
            O => \N__38813\,
            I => \N__38807\
        );

    \I__8063\ : InMux
    port map (
            O => \N__38812\,
            I => \N__38804\
        );

    \I__8062\ : LocalMux
    port map (
            O => \N__38807\,
            I => \N__38801\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__38804\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__8060\ : Odrv4
    port map (
            O => \N__38801\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__8059\ : CascadeMux
    port map (
            O => \N__38796\,
            I => \N__38793\
        );

    \I__8058\ : InMux
    port map (
            O => \N__38793\,
            I => \N__38787\
        );

    \I__8057\ : InMux
    port map (
            O => \N__38792\,
            I => \N__38787\
        );

    \I__8056\ : LocalMux
    port map (
            O => \N__38787\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\
        );

    \I__8055\ : InMux
    port map (
            O => \N__38784\,
            I => \N__38779\
        );

    \I__8054\ : InMux
    port map (
            O => \N__38783\,
            I => \N__38774\
        );

    \I__8053\ : InMux
    port map (
            O => \N__38782\,
            I => \N__38774\
        );

    \I__8052\ : LocalMux
    port map (
            O => \N__38779\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__8051\ : LocalMux
    port map (
            O => \N__38774\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__8050\ : CascadeMux
    port map (
            O => \N__38769\,
            I => \N__38766\
        );

    \I__8049\ : InMux
    port map (
            O => \N__38766\,
            I => \N__38763\
        );

    \I__8048\ : LocalMux
    port map (
            O => \N__38763\,
            I => \N__38760\
        );

    \I__8047\ : Odrv12
    port map (
            O => \N__38760\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt16\
        );

    \I__8046\ : CascadeMux
    port map (
            O => \N__38757\,
            I => \elapsed_time_ns_1_RNIQENQL1_0_9_cascade_\
        );

    \I__8045\ : InMux
    port map (
            O => \N__38754\,
            I => \N__38751\
        );

    \I__8044\ : LocalMux
    port map (
            O => \N__38751\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9\
        );

    \I__8043\ : CascadeMux
    port map (
            O => \N__38748\,
            I => \phase_controller_inst1.stoper_tr.N_242_cascade_\
        );

    \I__8042\ : InMux
    port map (
            O => \N__38745\,
            I => \N__38742\
        );

    \I__8041\ : LocalMux
    port map (
            O => \N__38742\,
            I => \N__38739\
        );

    \I__8040\ : Span4Mux_h
    port map (
            O => \N__38739\,
            I => \N__38736\
        );

    \I__8039\ : Odrv4
    port map (
            O => \N__38736\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\
        );

    \I__8038\ : InMux
    port map (
            O => \N__38733\,
            I => \N__38730\
        );

    \I__8037\ : LocalMux
    port map (
            O => \N__38730\,
            I => \N__38727\
        );

    \I__8036\ : Span4Mux_v
    port map (
            O => \N__38727\,
            I => \N__38724\
        );

    \I__8035\ : Span4Mux_h
    port map (
            O => \N__38724\,
            I => \N__38721\
        );

    \I__8034\ : Sp12to4
    port map (
            O => \N__38721\,
            I => \N__38718\
        );

    \I__8033\ : Odrv12
    port map (
            O => \N__38718\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\
        );

    \I__8032\ : InMux
    port map (
            O => \N__38715\,
            I => \N__38712\
        );

    \I__8031\ : LocalMux
    port map (
            O => \N__38712\,
            I => \N__38709\
        );

    \I__8030\ : Span4Mux_h
    port map (
            O => \N__38709\,
            I => \N__38706\
        );

    \I__8029\ : Odrv4
    port map (
            O => \N__38706\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9\
        );

    \I__8028\ : CascadeMux
    port map (
            O => \N__38703\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_\
        );

    \I__8027\ : InMux
    port map (
            O => \N__38700\,
            I => \N__38697\
        );

    \I__8026\ : LocalMux
    port map (
            O => \N__38697\,
            I => \N__38694\
        );

    \I__8025\ : Span4Mux_h
    port map (
            O => \N__38694\,
            I => \N__38691\
        );

    \I__8024\ : Odrv4
    port map (
            O => \N__38691\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\
        );

    \I__8023\ : InMux
    port map (
            O => \N__38688\,
            I => \N__38685\
        );

    \I__8022\ : LocalMux
    port map (
            O => \N__38685\,
            I => \N__38682\
        );

    \I__8021\ : Span4Mux_h
    port map (
            O => \N__38682\,
            I => \N__38679\
        );

    \I__8020\ : Odrv4
    port map (
            O => \N__38679\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\
        );

    \I__8019\ : CascadeMux
    port map (
            O => \N__38676\,
            I => \N__38673\
        );

    \I__8018\ : InMux
    port map (
            O => \N__38673\,
            I => \N__38669\
        );

    \I__8017\ : InMux
    port map (
            O => \N__38672\,
            I => \N__38666\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__38669\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\
        );

    \I__8015\ : LocalMux
    port map (
            O => \N__38666\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\
        );

    \I__8014\ : CascadeMux
    port map (
            O => \N__38661\,
            I => \N__38656\
        );

    \I__8013\ : InMux
    port map (
            O => \N__38660\,
            I => \N__38653\
        );

    \I__8012\ : InMux
    port map (
            O => \N__38659\,
            I => \N__38648\
        );

    \I__8011\ : InMux
    port map (
            O => \N__38656\,
            I => \N__38648\
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__38653\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__8009\ : LocalMux
    port map (
            O => \N__38648\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__8008\ : InMux
    port map (
            O => \N__38643\,
            I => \N__38638\
        );

    \I__8007\ : InMux
    port map (
            O => \N__38642\,
            I => \N__38635\
        );

    \I__8006\ : InMux
    port map (
            O => \N__38641\,
            I => \N__38632\
        );

    \I__8005\ : LocalMux
    port map (
            O => \N__38638\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__8004\ : LocalMux
    port map (
            O => \N__38635\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__8003\ : LocalMux
    port map (
            O => \N__38632\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__8002\ : CascadeMux
    port map (
            O => \N__38625\,
            I => \N__38622\
        );

    \I__8001\ : InMux
    port map (
            O => \N__38622\,
            I => \N__38619\
        );

    \I__8000\ : LocalMux
    port map (
            O => \N__38619\,
            I => \N__38616\
        );

    \I__7999\ : Span4Mux_h
    port map (
            O => \N__38616\,
            I => \N__38613\
        );

    \I__7998\ : Odrv4
    port map (
            O => \N__38613\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt18\
        );

    \I__7997\ : InMux
    port map (
            O => \N__38610\,
            I => \N__38604\
        );

    \I__7996\ : InMux
    port map (
            O => \N__38609\,
            I => \N__38604\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__38604\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\
        );

    \I__7994\ : InMux
    port map (
            O => \N__38601\,
            I => \N__38598\
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__38598\,
            I => \N__38595\
        );

    \I__7992\ : Odrv4
    port map (
            O => \N__38595\,
            I => \current_shift_inst.un38_control_input_0_s0_25\
        );

    \I__7991\ : InMux
    port map (
            O => \N__38592\,
            I => \current_shift_inst.un38_control_input_cry_24_s0\
        );

    \I__7990\ : InMux
    port map (
            O => \N__38589\,
            I => \N__38586\
        );

    \I__7989\ : LocalMux
    port map (
            O => \N__38586\,
            I => \N__38583\
        );

    \I__7988\ : Odrv4
    port map (
            O => \N__38583\,
            I => \current_shift_inst.un38_control_input_0_s0_26\
        );

    \I__7987\ : InMux
    port map (
            O => \N__38580\,
            I => \current_shift_inst.un38_control_input_cry_25_s0\
        );

    \I__7986\ : InMux
    port map (
            O => \N__38577\,
            I => \N__38574\
        );

    \I__7985\ : LocalMux
    port map (
            O => \N__38574\,
            I => \N__38571\
        );

    \I__7984\ : Odrv4
    port map (
            O => \N__38571\,
            I => \current_shift_inst.un38_control_input_0_s0_27\
        );

    \I__7983\ : InMux
    port map (
            O => \N__38568\,
            I => \current_shift_inst.un38_control_input_cry_26_s0\
        );

    \I__7982\ : InMux
    port map (
            O => \N__38565\,
            I => \N__38562\
        );

    \I__7981\ : LocalMux
    port map (
            O => \N__38562\,
            I => \N__38559\
        );

    \I__7980\ : Odrv4
    port map (
            O => \N__38559\,
            I => \current_shift_inst.un38_control_input_0_s0_28\
        );

    \I__7979\ : InMux
    port map (
            O => \N__38556\,
            I => \current_shift_inst.un38_control_input_cry_27_s0\
        );

    \I__7978\ : InMux
    port map (
            O => \N__38553\,
            I => \N__38550\
        );

    \I__7977\ : LocalMux
    port map (
            O => \N__38550\,
            I => \N__38547\
        );

    \I__7976\ : Odrv4
    port map (
            O => \N__38547\,
            I => \current_shift_inst.un38_control_input_0_s0_29\
        );

    \I__7975\ : InMux
    port map (
            O => \N__38544\,
            I => \current_shift_inst.un38_control_input_cry_28_s0\
        );

    \I__7974\ : InMux
    port map (
            O => \N__38541\,
            I => \N__38538\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__38538\,
            I => \N__38535\
        );

    \I__7972\ : Odrv4
    port map (
            O => \N__38535\,
            I => \current_shift_inst.un38_control_input_0_s0_30\
        );

    \I__7971\ : InMux
    port map (
            O => \N__38532\,
            I => \current_shift_inst.un38_control_input_cry_29_s0\
        );

    \I__7970\ : InMux
    port map (
            O => \N__38529\,
            I => \N__38525\
        );

    \I__7969\ : InMux
    port map (
            O => \N__38528\,
            I => \N__38522\
        );

    \I__7968\ : LocalMux
    port map (
            O => \N__38525\,
            I => \N__38515\
        );

    \I__7967\ : LocalMux
    port map (
            O => \N__38522\,
            I => \N__38509\
        );

    \I__7966\ : InMux
    port map (
            O => \N__38521\,
            I => \N__38500\
        );

    \I__7965\ : InMux
    port map (
            O => \N__38520\,
            I => \N__38500\
        );

    \I__7964\ : InMux
    port map (
            O => \N__38519\,
            I => \N__38500\
        );

    \I__7963\ : InMux
    port map (
            O => \N__38518\,
            I => \N__38500\
        );

    \I__7962\ : Span4Mux_h
    port map (
            O => \N__38515\,
            I => \N__38491\
        );

    \I__7961\ : InMux
    port map (
            O => \N__38514\,
            I => \N__38484\
        );

    \I__7960\ : InMux
    port map (
            O => \N__38513\,
            I => \N__38484\
        );

    \I__7959\ : InMux
    port map (
            O => \N__38512\,
            I => \N__38484\
        );

    \I__7958\ : Span4Mux_v
    port map (
            O => \N__38509\,
            I => \N__38479\
        );

    \I__7957\ : LocalMux
    port map (
            O => \N__38500\,
            I => \N__38479\
        );

    \I__7956\ : InMux
    port map (
            O => \N__38499\,
            I => \N__38468\
        );

    \I__7955\ : InMux
    port map (
            O => \N__38498\,
            I => \N__38468\
        );

    \I__7954\ : InMux
    port map (
            O => \N__38497\,
            I => \N__38468\
        );

    \I__7953\ : InMux
    port map (
            O => \N__38496\,
            I => \N__38468\
        );

    \I__7952\ : InMux
    port map (
            O => \N__38495\,
            I => \N__38468\
        );

    \I__7951\ : InMux
    port map (
            O => \N__38494\,
            I => \N__38465\
        );

    \I__7950\ : Odrv4
    port map (
            O => \N__38491\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__7949\ : LocalMux
    port map (
            O => \N__38484\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__7948\ : Odrv4
    port map (
            O => \N__38479\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__7947\ : LocalMux
    port map (
            O => \N__38468\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__7946\ : LocalMux
    port map (
            O => \N__38465\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__7945\ : InMux
    port map (
            O => \N__38454\,
            I => \current_shift_inst.un38_control_input_cry_30_s0\
        );

    \I__7944\ : InMux
    port map (
            O => \N__38451\,
            I => \N__38448\
        );

    \I__7943\ : LocalMux
    port map (
            O => \N__38448\,
            I => \N__38445\
        );

    \I__7942\ : Span4Mux_h
    port map (
            O => \N__38445\,
            I => \N__38442\
        );

    \I__7941\ : Odrv4
    port map (
            O => \N__38442\,
            I => \current_shift_inst.control_input_axb_11\
        );

    \I__7940\ : InMux
    port map (
            O => \N__38439\,
            I => \N__38436\
        );

    \I__7939\ : LocalMux
    port map (
            O => \N__38436\,
            I => \N__38433\
        );

    \I__7938\ : Span4Mux_h
    port map (
            O => \N__38433\,
            I => \N__38430\
        );

    \I__7937\ : Odrv4
    port map (
            O => \N__38430\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\
        );

    \I__7936\ : InMux
    port map (
            O => \N__38427\,
            I => \N__38424\
        );

    \I__7935\ : LocalMux
    port map (
            O => \N__38424\,
            I => \N__38421\
        );

    \I__7934\ : Odrv12
    port map (
            O => \N__38421\,
            I => \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\
        );

    \I__7933\ : InMux
    port map (
            O => \N__38418\,
            I => \N__38415\
        );

    \I__7932\ : LocalMux
    port map (
            O => \N__38415\,
            I => \N__38412\
        );

    \I__7931\ : Span4Mux_h
    port map (
            O => \N__38412\,
            I => \N__38409\
        );

    \I__7930\ : Odrv4
    port map (
            O => \N__38409\,
            I => \current_shift_inst.un38_control_input_0_s0_20\
        );

    \I__7929\ : InMux
    port map (
            O => \N__38406\,
            I => \current_shift_inst.un38_control_input_cry_19_s0\
        );

    \I__7928\ : InMux
    port map (
            O => \N__38403\,
            I => \N__38400\
        );

    \I__7927\ : LocalMux
    port map (
            O => \N__38400\,
            I => \N__38397\
        );

    \I__7926\ : Odrv4
    port map (
            O => \N__38397\,
            I => \current_shift_inst.un38_control_input_0_s0_21\
        );

    \I__7925\ : InMux
    port map (
            O => \N__38394\,
            I => \current_shift_inst.un38_control_input_cry_20_s0\
        );

    \I__7924\ : InMux
    port map (
            O => \N__38391\,
            I => \N__38388\
        );

    \I__7923\ : LocalMux
    port map (
            O => \N__38388\,
            I => \N__38385\
        );

    \I__7922\ : Odrv4
    port map (
            O => \N__38385\,
            I => \current_shift_inst.un38_control_input_0_s0_22\
        );

    \I__7921\ : InMux
    port map (
            O => \N__38382\,
            I => \current_shift_inst.un38_control_input_cry_21_s0\
        );

    \I__7920\ : InMux
    port map (
            O => \N__38379\,
            I => \N__38376\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__38376\,
            I => \N__38373\
        );

    \I__7918\ : Odrv4
    port map (
            O => \N__38373\,
            I => \current_shift_inst.un38_control_input_0_s0_23\
        );

    \I__7917\ : InMux
    port map (
            O => \N__38370\,
            I => \current_shift_inst.un38_control_input_cry_22_s0\
        );

    \I__7916\ : InMux
    port map (
            O => \N__38367\,
            I => \N__38364\
        );

    \I__7915\ : LocalMux
    port map (
            O => \N__38364\,
            I => \N__38361\
        );

    \I__7914\ : Odrv4
    port map (
            O => \N__38361\,
            I => \current_shift_inst.un38_control_input_0_s0_24\
        );

    \I__7913\ : InMux
    port map (
            O => \N__38358\,
            I => \bfn_15_15_0_\
        );

    \I__7912\ : CascadeMux
    port map (
            O => \N__38355\,
            I => \N__38352\
        );

    \I__7911\ : InMux
    port map (
            O => \N__38352\,
            I => \N__38349\
        );

    \I__7910\ : LocalMux
    port map (
            O => \N__38349\,
            I => \N__38346\
        );

    \I__7909\ : Span4Mux_v
    port map (
            O => \N__38346\,
            I => \N__38343\
        );

    \I__7908\ : Odrv4
    port map (
            O => \N__38343\,
            I => \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\
        );

    \I__7907\ : InMux
    port map (
            O => \N__38340\,
            I => \N__38337\
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__38337\,
            I => \N__38334\
        );

    \I__7905\ : Span4Mux_v
    port map (
            O => \N__38334\,
            I => \N__38331\
        );

    \I__7904\ : Odrv4
    port map (
            O => \N__38331\,
            I => \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\
        );

    \I__7903\ : InMux
    port map (
            O => \N__38328\,
            I => \current_shift_inst.un10_control_input_cry_30\
        );

    \I__7902\ : CascadeMux
    port map (
            O => \N__38325\,
            I => \N__38322\
        );

    \I__7901\ : InMux
    port map (
            O => \N__38322\,
            I => \N__38319\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__38319\,
            I => \N__38316\
        );

    \I__7899\ : Odrv12
    port map (
            O => \N__38316\,
            I => \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\
        );

    \I__7898\ : InMux
    port map (
            O => \N__38313\,
            I => \N__38310\
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__38310\,
            I => \N__38307\
        );

    \I__7896\ : Span4Mux_v
    port map (
            O => \N__38307\,
            I => \N__38304\
        );

    \I__7895\ : Odrv4
    port map (
            O => \N__38304\,
            I => \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\
        );

    \I__7894\ : InMux
    port map (
            O => \N__38301\,
            I => \N__38298\
        );

    \I__7893\ : LocalMux
    port map (
            O => \N__38298\,
            I => \N__38295\
        );

    \I__7892\ : Span4Mux_v
    port map (
            O => \N__38295\,
            I => \N__38292\
        );

    \I__7891\ : Odrv4
    port map (
            O => \N__38292\,
            I => \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\
        );

    \I__7890\ : InMux
    port map (
            O => \N__38289\,
            I => \N__38286\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__38286\,
            I => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\
        );

    \I__7888\ : InMux
    port map (
            O => \N__38283\,
            I => \N__38271\
        );

    \I__7887\ : InMux
    port map (
            O => \N__38282\,
            I => \N__38267\
        );

    \I__7886\ : InMux
    port map (
            O => \N__38281\,
            I => \N__38260\
        );

    \I__7885\ : InMux
    port map (
            O => \N__38280\,
            I => \N__38260\
        );

    \I__7884\ : InMux
    port map (
            O => \N__38279\,
            I => \N__38260\
        );

    \I__7883\ : InMux
    port map (
            O => \N__38278\,
            I => \N__38251\
        );

    \I__7882\ : InMux
    port map (
            O => \N__38277\,
            I => \N__38251\
        );

    \I__7881\ : InMux
    port map (
            O => \N__38276\,
            I => \N__38251\
        );

    \I__7880\ : InMux
    port map (
            O => \N__38275\,
            I => \N__38251\
        );

    \I__7879\ : InMux
    port map (
            O => \N__38274\,
            I => \N__38240\
        );

    \I__7878\ : LocalMux
    port map (
            O => \N__38271\,
            I => \N__38237\
        );

    \I__7877\ : InMux
    port map (
            O => \N__38270\,
            I => \N__38233\
        );

    \I__7876\ : LocalMux
    port map (
            O => \N__38267\,
            I => \N__38226\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__38260\,
            I => \N__38226\
        );

    \I__7874\ : LocalMux
    port map (
            O => \N__38251\,
            I => \N__38226\
        );

    \I__7873\ : InMux
    port map (
            O => \N__38250\,
            I => \N__38223\
        );

    \I__7872\ : InMux
    port map (
            O => \N__38249\,
            I => \N__38216\
        );

    \I__7871\ : InMux
    port map (
            O => \N__38248\,
            I => \N__38216\
        );

    \I__7870\ : InMux
    port map (
            O => \N__38247\,
            I => \N__38216\
        );

    \I__7869\ : InMux
    port map (
            O => \N__38246\,
            I => \N__38207\
        );

    \I__7868\ : InMux
    port map (
            O => \N__38245\,
            I => \N__38207\
        );

    \I__7867\ : InMux
    port map (
            O => \N__38244\,
            I => \N__38207\
        );

    \I__7866\ : InMux
    port map (
            O => \N__38243\,
            I => \N__38207\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__38240\,
            I => \N__38204\
        );

    \I__7864\ : Span4Mux_s2_h
    port map (
            O => \N__38237\,
            I => \N__38201\
        );

    \I__7863\ : InMux
    port map (
            O => \N__38236\,
            I => \N__38195\
        );

    \I__7862\ : LocalMux
    port map (
            O => \N__38233\,
            I => \N__38189\
        );

    \I__7861\ : Span4Mux_v
    port map (
            O => \N__38226\,
            I => \N__38180\
        );

    \I__7860\ : LocalMux
    port map (
            O => \N__38223\,
            I => \N__38180\
        );

    \I__7859\ : LocalMux
    port map (
            O => \N__38216\,
            I => \N__38180\
        );

    \I__7858\ : LocalMux
    port map (
            O => \N__38207\,
            I => \N__38180\
        );

    \I__7857\ : Span12Mux_s2_h
    port map (
            O => \N__38204\,
            I => \N__38175\
        );

    \I__7856\ : Sp12to4
    port map (
            O => \N__38201\,
            I => \N__38175\
        );

    \I__7855\ : InMux
    port map (
            O => \N__38200\,
            I => \N__38172\
        );

    \I__7854\ : InMux
    port map (
            O => \N__38199\,
            I => \N__38167\
        );

    \I__7853\ : InMux
    port map (
            O => \N__38198\,
            I => \N__38167\
        );

    \I__7852\ : LocalMux
    port map (
            O => \N__38195\,
            I => \N__38164\
        );

    \I__7851\ : CascadeMux
    port map (
            O => \N__38194\,
            I => \N__38158\
        );

    \I__7850\ : CascadeMux
    port map (
            O => \N__38193\,
            I => \N__38154\
        );

    \I__7849\ : CascadeMux
    port map (
            O => \N__38192\,
            I => \N__38150\
        );

    \I__7848\ : Span12Mux_s6_h
    port map (
            O => \N__38189\,
            I => \N__38135\
        );

    \I__7847\ : Span4Mux_v
    port map (
            O => \N__38180\,
            I => \N__38132\
        );

    \I__7846\ : Span12Mux_v
    port map (
            O => \N__38175\,
            I => \N__38125\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__38172\,
            I => \N__38125\
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__38167\,
            I => \N__38125\
        );

    \I__7843\ : Span12Mux_s11_h
    port map (
            O => \N__38164\,
            I => \N__38122\
        );

    \I__7842\ : InMux
    port map (
            O => \N__38163\,
            I => \N__38117\
        );

    \I__7841\ : InMux
    port map (
            O => \N__38162\,
            I => \N__38117\
        );

    \I__7840\ : InMux
    port map (
            O => \N__38161\,
            I => \N__38102\
        );

    \I__7839\ : InMux
    port map (
            O => \N__38158\,
            I => \N__38102\
        );

    \I__7838\ : InMux
    port map (
            O => \N__38157\,
            I => \N__38102\
        );

    \I__7837\ : InMux
    port map (
            O => \N__38154\,
            I => \N__38102\
        );

    \I__7836\ : InMux
    port map (
            O => \N__38153\,
            I => \N__38102\
        );

    \I__7835\ : InMux
    port map (
            O => \N__38150\,
            I => \N__38102\
        );

    \I__7834\ : InMux
    port map (
            O => \N__38149\,
            I => \N__38102\
        );

    \I__7833\ : CascadeMux
    port map (
            O => \N__38148\,
            I => \N__38099\
        );

    \I__7832\ : CascadeMux
    port map (
            O => \N__38147\,
            I => \N__38095\
        );

    \I__7831\ : CascadeMux
    port map (
            O => \N__38146\,
            I => \N__38091\
        );

    \I__7830\ : CascadeMux
    port map (
            O => \N__38145\,
            I => \N__38087\
        );

    \I__7829\ : CascadeMux
    port map (
            O => \N__38144\,
            I => \N__38083\
        );

    \I__7828\ : CascadeMux
    port map (
            O => \N__38143\,
            I => \N__38079\
        );

    \I__7827\ : CascadeMux
    port map (
            O => \N__38142\,
            I => \N__38075\
        );

    \I__7826\ : CascadeMux
    port map (
            O => \N__38141\,
            I => \N__38071\
        );

    \I__7825\ : CascadeMux
    port map (
            O => \N__38140\,
            I => \N__38066\
        );

    \I__7824\ : CascadeMux
    port map (
            O => \N__38139\,
            I => \N__38062\
        );

    \I__7823\ : CascadeMux
    port map (
            O => \N__38138\,
            I => \N__38058\
        );

    \I__7822\ : Span12Mux_v
    port map (
            O => \N__38135\,
            I => \N__38054\
        );

    \I__7821\ : Sp12to4
    port map (
            O => \N__38132\,
            I => \N__38051\
        );

    \I__7820\ : Span12Mux_v
    port map (
            O => \N__38125\,
            I => \N__38048\
        );

    \I__7819\ : Span12Mux_v
    port map (
            O => \N__38122\,
            I => \N__38043\
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__38117\,
            I => \N__38043\
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__38102\,
            I => \N__38040\
        );

    \I__7816\ : InMux
    port map (
            O => \N__38099\,
            I => \N__38023\
        );

    \I__7815\ : InMux
    port map (
            O => \N__38098\,
            I => \N__38023\
        );

    \I__7814\ : InMux
    port map (
            O => \N__38095\,
            I => \N__38023\
        );

    \I__7813\ : InMux
    port map (
            O => \N__38094\,
            I => \N__38023\
        );

    \I__7812\ : InMux
    port map (
            O => \N__38091\,
            I => \N__38023\
        );

    \I__7811\ : InMux
    port map (
            O => \N__38090\,
            I => \N__38023\
        );

    \I__7810\ : InMux
    port map (
            O => \N__38087\,
            I => \N__38023\
        );

    \I__7809\ : InMux
    port map (
            O => \N__38086\,
            I => \N__38023\
        );

    \I__7808\ : InMux
    port map (
            O => \N__38083\,
            I => \N__38006\
        );

    \I__7807\ : InMux
    port map (
            O => \N__38082\,
            I => \N__38006\
        );

    \I__7806\ : InMux
    port map (
            O => \N__38079\,
            I => \N__38006\
        );

    \I__7805\ : InMux
    port map (
            O => \N__38078\,
            I => \N__38006\
        );

    \I__7804\ : InMux
    port map (
            O => \N__38075\,
            I => \N__38006\
        );

    \I__7803\ : InMux
    port map (
            O => \N__38074\,
            I => \N__38006\
        );

    \I__7802\ : InMux
    port map (
            O => \N__38071\,
            I => \N__38006\
        );

    \I__7801\ : InMux
    port map (
            O => \N__38070\,
            I => \N__38006\
        );

    \I__7800\ : InMux
    port map (
            O => \N__38069\,
            I => \N__37991\
        );

    \I__7799\ : InMux
    port map (
            O => \N__38066\,
            I => \N__37991\
        );

    \I__7798\ : InMux
    port map (
            O => \N__38065\,
            I => \N__37991\
        );

    \I__7797\ : InMux
    port map (
            O => \N__38062\,
            I => \N__37991\
        );

    \I__7796\ : InMux
    port map (
            O => \N__38061\,
            I => \N__37991\
        );

    \I__7795\ : InMux
    port map (
            O => \N__38058\,
            I => \N__37991\
        );

    \I__7794\ : InMux
    port map (
            O => \N__38057\,
            I => \N__37991\
        );

    \I__7793\ : Span12Mux_v
    port map (
            O => \N__38054\,
            I => \N__37986\
        );

    \I__7792\ : Span12Mux_s6_h
    port map (
            O => \N__38051\,
            I => \N__37986\
        );

    \I__7791\ : Span12Mux_h
    port map (
            O => \N__38048\,
            I => \N__37981\
        );

    \I__7790\ : Span12Mux_v
    port map (
            O => \N__38043\,
            I => \N__37981\
        );

    \I__7789\ : Span12Mux_v
    port map (
            O => \N__38040\,
            I => \N__37972\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__38023\,
            I => \N__37972\
        );

    \I__7787\ : LocalMux
    port map (
            O => \N__38006\,
            I => \N__37972\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__37991\,
            I => \N__37972\
        );

    \I__7785\ : Odrv12
    port map (
            O => \N__37986\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7784\ : Odrv12
    port map (
            O => \N__37981\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7783\ : Odrv12
    port map (
            O => \N__37972\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7782\ : InMux
    port map (
            O => \N__37965\,
            I => \N__37962\
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__37962\,
            I => \N__37959\
        );

    \I__7780\ : Odrv4
    port map (
            O => \N__37959\,
            I => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\
        );

    \I__7779\ : CascadeMux
    port map (
            O => \N__37956\,
            I => \N__37953\
        );

    \I__7778\ : InMux
    port map (
            O => \N__37953\,
            I => \N__37950\
        );

    \I__7777\ : LocalMux
    port map (
            O => \N__37950\,
            I => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\
        );

    \I__7776\ : InMux
    port map (
            O => \N__37947\,
            I => \N__37944\
        );

    \I__7775\ : LocalMux
    port map (
            O => \N__37944\,
            I => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\
        );

    \I__7774\ : InMux
    port map (
            O => \N__37941\,
            I => \N__37938\
        );

    \I__7773\ : LocalMux
    port map (
            O => \N__37938\,
            I => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\
        );

    \I__7772\ : CascadeMux
    port map (
            O => \N__37935\,
            I => \N__37932\
        );

    \I__7771\ : InMux
    port map (
            O => \N__37932\,
            I => \N__37929\
        );

    \I__7770\ : LocalMux
    port map (
            O => \N__37929\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__7769\ : InMux
    port map (
            O => \N__37926\,
            I => \N__37923\
        );

    \I__7768\ : LocalMux
    port map (
            O => \N__37923\,
            I => \N__37919\
        );

    \I__7767\ : InMux
    port map (
            O => \N__37922\,
            I => \N__37916\
        );

    \I__7766\ : Sp12to4
    port map (
            O => \N__37919\,
            I => \N__37910\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__37916\,
            I => \N__37910\
        );

    \I__7764\ : InMux
    port map (
            O => \N__37915\,
            I => \N__37907\
        );

    \I__7763\ : Span12Mux_v
    port map (
            O => \N__37910\,
            I => \N__37904\
        );

    \I__7762\ : LocalMux
    port map (
            O => \N__37907\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\
        );

    \I__7761\ : Odrv12
    port map (
            O => \N__37904\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\
        );

    \I__7760\ : CascadeMux
    port map (
            O => \N__37899\,
            I => \N__37896\
        );

    \I__7759\ : InMux
    port map (
            O => \N__37896\,
            I => \N__37892\
        );

    \I__7758\ : InMux
    port map (
            O => \N__37895\,
            I => \N__37888\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__37892\,
            I => \N__37885\
        );

    \I__7756\ : CascadeMux
    port map (
            O => \N__37891\,
            I => \N__37882\
        );

    \I__7755\ : LocalMux
    port map (
            O => \N__37888\,
            I => \N__37878\
        );

    \I__7754\ : Span4Mux_v
    port map (
            O => \N__37885\,
            I => \N__37874\
        );

    \I__7753\ : InMux
    port map (
            O => \N__37882\,
            I => \N__37869\
        );

    \I__7752\ : InMux
    port map (
            O => \N__37881\,
            I => \N__37869\
        );

    \I__7751\ : Span4Mux_v
    port map (
            O => \N__37878\,
            I => \N__37866\
        );

    \I__7750\ : InMux
    port map (
            O => \N__37877\,
            I => \N__37863\
        );

    \I__7749\ : Span4Mux_h
    port map (
            O => \N__37874\,
            I => \N__37860\
        );

    \I__7748\ : LocalMux
    port map (
            O => \N__37869\,
            I => \N__37855\
        );

    \I__7747\ : Span4Mux_h
    port map (
            O => \N__37866\,
            I => \N__37855\
        );

    \I__7746\ : LocalMux
    port map (
            O => \N__37863\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__7745\ : Odrv4
    port map (
            O => \N__37860\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__7744\ : Odrv4
    port map (
            O => \N__37855\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__7743\ : InMux
    port map (
            O => \N__37848\,
            I => \N__37845\
        );

    \I__7742\ : LocalMux
    port map (
            O => \N__37845\,
            I => \N__37842\
        );

    \I__7741\ : Span4Mux_h
    port map (
            O => \N__37842\,
            I => \N__37839\
        );

    \I__7740\ : Span4Mux_v
    port map (
            O => \N__37839\,
            I => \N__37836\
        );

    \I__7739\ : Odrv4
    port map (
            O => \N__37836\,
            I => \current_shift_inst.PI_CTRL.integrator_i_11\
        );

    \I__7738\ : InMux
    port map (
            O => \N__37833\,
            I => \N__37829\
        );

    \I__7737\ : InMux
    port map (
            O => \N__37832\,
            I => \N__37826\
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__37829\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__7735\ : LocalMux
    port map (
            O => \N__37826\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__7734\ : InMux
    port map (
            O => \N__37821\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\
        );

    \I__7733\ : InMux
    port map (
            O => \N__37818\,
            I => \N__37814\
        );

    \I__7732\ : InMux
    port map (
            O => \N__37817\,
            I => \N__37811\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__37814\,
            I => \N__37808\
        );

    \I__7730\ : LocalMux
    port map (
            O => \N__37811\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__7729\ : Odrv4
    port map (
            O => \N__37808\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__7728\ : InMux
    port map (
            O => \N__37803\,
            I => \bfn_14_24_0_\
        );

    \I__7727\ : InMux
    port map (
            O => \N__37800\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\
        );

    \I__7726\ : InMux
    port map (
            O => \N__37797\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\
        );

    \I__7725\ : InMux
    port map (
            O => \N__37794\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\
        );

    \I__7724\ : InMux
    port map (
            O => \N__37791\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\
        );

    \I__7723\ : InMux
    port map (
            O => \N__37788\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\
        );

    \I__7722\ : InMux
    port map (
            O => \N__37785\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\
        );

    \I__7721\ : InMux
    port map (
            O => \N__37782\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__7720\ : InMux
    port map (
            O => \N__37779\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__7719\ : InMux
    port map (
            O => \N__37776\,
            I => \bfn_14_23_0_\
        );

    \I__7718\ : InMux
    port map (
            O => \N__37773\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__7717\ : InMux
    port map (
            O => \N__37770\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__7716\ : InMux
    port map (
            O => \N__37767\,
            I => \N__37763\
        );

    \I__7715\ : InMux
    port map (
            O => \N__37766\,
            I => \N__37760\
        );

    \I__7714\ : LocalMux
    port map (
            O => \N__37763\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__37760\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__7712\ : InMux
    port map (
            O => \N__37755\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\
        );

    \I__7711\ : InMux
    port map (
            O => \N__37752\,
            I => \N__37748\
        );

    \I__7710\ : InMux
    port map (
            O => \N__37751\,
            I => \N__37745\
        );

    \I__7709\ : LocalMux
    port map (
            O => \N__37748\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__37745\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__7707\ : InMux
    port map (
            O => \N__37740\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__7706\ : InMux
    port map (
            O => \N__37737\,
            I => \N__37733\
        );

    \I__7705\ : InMux
    port map (
            O => \N__37736\,
            I => \N__37730\
        );

    \I__7704\ : LocalMux
    port map (
            O => \N__37733\,
            I => \N__37727\
        );

    \I__7703\ : LocalMux
    port map (
            O => \N__37730\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__7702\ : Odrv4
    port map (
            O => \N__37727\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__7701\ : InMux
    port map (
            O => \N__37722\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\
        );

    \I__7700\ : InMux
    port map (
            O => \N__37719\,
            I => \N__37716\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__37716\,
            I => \N__37712\
        );

    \I__7698\ : InMux
    port map (
            O => \N__37715\,
            I => \N__37709\
        );

    \I__7697\ : Span4Mux_h
    port map (
            O => \N__37712\,
            I => \N__37706\
        );

    \I__7696\ : LocalMux
    port map (
            O => \N__37709\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__7695\ : Odrv4
    port map (
            O => \N__37706\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__7694\ : InMux
    port map (
            O => \N__37701\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\
        );

    \I__7693\ : InMux
    port map (
            O => \N__37698\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__7692\ : InMux
    port map (
            O => \N__37695\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__7691\ : InMux
    port map (
            O => \N__37692\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__7690\ : InMux
    port map (
            O => \N__37689\,
            I => \bfn_14_22_0_\
        );

    \I__7689\ : InMux
    port map (
            O => \N__37686\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__7688\ : InMux
    port map (
            O => \N__37683\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__7687\ : InMux
    port map (
            O => \N__37680\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__7686\ : InMux
    port map (
            O => \N__37677\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__7685\ : InMux
    port map (
            O => \N__37674\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__7684\ : CascadeMux
    port map (
            O => \N__37671\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\
        );

    \I__7683\ : InMux
    port map (
            O => \N__37668\,
            I => \N__37662\
        );

    \I__7682\ : InMux
    port map (
            O => \N__37667\,
            I => \N__37662\
        );

    \I__7681\ : LocalMux
    port map (
            O => \N__37662\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__7680\ : CascadeMux
    port map (
            O => \N__37659\,
            I => \N__37656\
        );

    \I__7679\ : InMux
    port map (
            O => \N__37656\,
            I => \N__37649\
        );

    \I__7678\ : InMux
    port map (
            O => \N__37655\,
            I => \N__37644\
        );

    \I__7677\ : InMux
    port map (
            O => \N__37654\,
            I => \N__37644\
        );

    \I__7676\ : InMux
    port map (
            O => \N__37653\,
            I => \N__37639\
        );

    \I__7675\ : InMux
    port map (
            O => \N__37652\,
            I => \N__37639\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__37649\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__7673\ : LocalMux
    port map (
            O => \N__37644\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__7672\ : LocalMux
    port map (
            O => \N__37639\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__7671\ : CascadeMux
    port map (
            O => \N__37632\,
            I => \N__37627\
        );

    \I__7670\ : InMux
    port map (
            O => \N__37631\,
            I => \N__37622\
        );

    \I__7669\ : InMux
    port map (
            O => \N__37630\,
            I => \N__37613\
        );

    \I__7668\ : InMux
    port map (
            O => \N__37627\,
            I => \N__37613\
        );

    \I__7667\ : InMux
    port map (
            O => \N__37626\,
            I => \N__37613\
        );

    \I__7666\ : InMux
    port map (
            O => \N__37625\,
            I => \N__37613\
        );

    \I__7665\ : LocalMux
    port map (
            O => \N__37622\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__37613\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__7663\ : InMux
    port map (
            O => \N__37608\,
            I => \N__37604\
        );

    \I__7662\ : InMux
    port map (
            O => \N__37607\,
            I => \N__37601\
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__37604\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__7660\ : LocalMux
    port map (
            O => \N__37601\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__7659\ : InMux
    port map (
            O => \N__37596\,
            I => \N__37593\
        );

    \I__7658\ : LocalMux
    port map (
            O => \N__37593\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\
        );

    \I__7657\ : InMux
    port map (
            O => \N__37590\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__7656\ : CascadeMux
    port map (
            O => \N__37587\,
            I => \N__37584\
        );

    \I__7655\ : InMux
    port map (
            O => \N__37584\,
            I => \N__37581\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__37581\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIJF7V2Z0Z_28\
        );

    \I__7653\ : InMux
    port map (
            O => \N__37578\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__7652\ : InMux
    port map (
            O => \N__37575\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__7651\ : InMux
    port map (
            O => \N__37572\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__7650\ : InMux
    port map (
            O => \N__37569\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\
        );

    \I__7649\ : InMux
    port map (
            O => \N__37566\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\
        );

    \I__7648\ : InMux
    port map (
            O => \N__37563\,
            I => \N__37560\
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__37560\,
            I => \N__37556\
        );

    \I__7646\ : InMux
    port map (
            O => \N__37559\,
            I => \N__37553\
        );

    \I__7645\ : Span4Mux_h
    port map (
            O => \N__37556\,
            I => \N__37550\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__37553\,
            I => \N__37547\
        );

    \I__7643\ : Sp12to4
    port map (
            O => \N__37550\,
            I => \N__37540\
        );

    \I__7642\ : Sp12to4
    port map (
            O => \N__37547\,
            I => \N__37540\
        );

    \I__7641\ : InMux
    port map (
            O => \N__37546\,
            I => \N__37535\
        );

    \I__7640\ : InMux
    port map (
            O => \N__37545\,
            I => \N__37535\
        );

    \I__7639\ : Span12Mux_v
    port map (
            O => \N__37540\,
            I => \N__37532\
        );

    \I__7638\ : LocalMux
    port map (
            O => \N__37535\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__7637\ : Odrv12
    port map (
            O => \N__37532\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__7636\ : InMux
    port map (
            O => \N__37527\,
            I => \N__37524\
        );

    \I__7635\ : LocalMux
    port map (
            O => \N__37524\,
            I => \N__37520\
        );

    \I__7634\ : InMux
    port map (
            O => \N__37523\,
            I => \N__37517\
        );

    \I__7633\ : Span4Mux_v
    port map (
            O => \N__37520\,
            I => \N__37514\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__37517\,
            I => \N__37511\
        );

    \I__7631\ : Span4Mux_v
    port map (
            O => \N__37514\,
            I => \N__37508\
        );

    \I__7630\ : Span12Mux_v
    port map (
            O => \N__37511\,
            I => \N__37504\
        );

    \I__7629\ : Span4Mux_v
    port map (
            O => \N__37508\,
            I => \N__37501\
        );

    \I__7628\ : InMux
    port map (
            O => \N__37507\,
            I => \N__37498\
        );

    \I__7627\ : Odrv12
    port map (
            O => \N__37504\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__7626\ : Odrv4
    port map (
            O => \N__37501\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__7625\ : LocalMux
    port map (
            O => \N__37498\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__7624\ : CascadeMux
    port map (
            O => \N__37491\,
            I => \N__37488\
        );

    \I__7623\ : InMux
    port map (
            O => \N__37488\,
            I => \N__37485\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__37485\,
            I => \N__37479\
        );

    \I__7621\ : InMux
    port map (
            O => \N__37484\,
            I => \N__37476\
        );

    \I__7620\ : InMux
    port map (
            O => \N__37483\,
            I => \N__37473\
        );

    \I__7619\ : InMux
    port map (
            O => \N__37482\,
            I => \N__37470\
        );

    \I__7618\ : Span4Mux_h
    port map (
            O => \N__37479\,
            I => \N__37467\
        );

    \I__7617\ : LocalMux
    port map (
            O => \N__37476\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__37473\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__37470\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__7614\ : Odrv4
    port map (
            O => \N__37467\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__7613\ : InMux
    port map (
            O => \N__37458\,
            I => \N__37453\
        );

    \I__7612\ : InMux
    port map (
            O => \N__37457\,
            I => \N__37450\
        );

    \I__7611\ : InMux
    port map (
            O => \N__37456\,
            I => \N__37447\
        );

    \I__7610\ : LocalMux
    port map (
            O => \N__37453\,
            I => \N__37444\
        );

    \I__7609\ : LocalMux
    port map (
            O => \N__37450\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__7608\ : LocalMux
    port map (
            O => \N__37447\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__7607\ : Odrv4
    port map (
            O => \N__37444\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__7606\ : CascadeMux
    port map (
            O => \N__37437\,
            I => \N__37434\
        );

    \I__7605\ : InMux
    port map (
            O => \N__37434\,
            I => \N__37431\
        );

    \I__7604\ : LocalMux
    port map (
            O => \N__37431\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\
        );

    \I__7603\ : InMux
    port map (
            O => \N__37428\,
            I => \N__37424\
        );

    \I__7602\ : InMux
    port map (
            O => \N__37427\,
            I => \N__37421\
        );

    \I__7601\ : LocalMux
    port map (
            O => \N__37424\,
            I => \N__37418\
        );

    \I__7600\ : LocalMux
    port map (
            O => \N__37421\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__7599\ : Odrv4
    port map (
            O => \N__37418\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__7598\ : InMux
    port map (
            O => \N__37413\,
            I => \N__37409\
        );

    \I__7597\ : InMux
    port map (
            O => \N__37412\,
            I => \N__37406\
        );

    \I__7596\ : LocalMux
    port map (
            O => \N__37409\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__7595\ : LocalMux
    port map (
            O => \N__37406\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__7594\ : InMux
    port map (
            O => \N__37401\,
            I => \N__37398\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__37398\,
            I => \phase_controller_inst2.stoper_tr.un4_running_df24\
        );

    \I__7592\ : CascadeMux
    port map (
            O => \N__37395\,
            I => \N__37392\
        );

    \I__7591\ : InMux
    port map (
            O => \N__37392\,
            I => \N__37389\
        );

    \I__7590\ : LocalMux
    port map (
            O => \N__37389\,
            I => \N__37386\
        );

    \I__7589\ : Span4Mux_v
    port map (
            O => \N__37386\,
            I => \N__37383\
        );

    \I__7588\ : Odrv4
    port map (
            O => \N__37383\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\
        );

    \I__7587\ : InMux
    port map (
            O => \N__37380\,
            I => \N__37377\
        );

    \I__7586\ : LocalMux
    port map (
            O => \N__37377\,
            I => \N__37374\
        );

    \I__7585\ : Odrv4
    port map (
            O => \N__37374\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\
        );

    \I__7584\ : InMux
    port map (
            O => \N__37371\,
            I => \N__37368\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__37368\,
            I => \N__37365\
        );

    \I__7582\ : Span4Mux_h
    port map (
            O => \N__37365\,
            I => \N__37362\
        );

    \I__7581\ : Odrv4
    port map (
            O => \N__37362\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\
        );

    \I__7580\ : InMux
    port map (
            O => \N__37359\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__7579\ : InMux
    port map (
            O => \N__37356\,
            I => \N__37352\
        );

    \I__7578\ : InMux
    port map (
            O => \N__37355\,
            I => \N__37349\
        );

    \I__7577\ : LocalMux
    port map (
            O => \N__37352\,
            I => \N__37346\
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__37349\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__7575\ : Odrv4
    port map (
            O => \N__37346\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__7574\ : InMux
    port map (
            O => \N__37341\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\
        );

    \I__7573\ : InMux
    port map (
            O => \N__37338\,
            I => \N__37334\
        );

    \I__7572\ : InMux
    port map (
            O => \N__37337\,
            I => \N__37331\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__37334\,
            I => \N__37328\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__37331\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__7569\ : Odrv4
    port map (
            O => \N__37328\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__7568\ : InMux
    port map (
            O => \N__37323\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\
        );

    \I__7567\ : InMux
    port map (
            O => \N__37320\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\
        );

    \I__7566\ : InMux
    port map (
            O => \N__37317\,
            I => \bfn_14_17_0_\
        );

    \I__7565\ : InMux
    port map (
            O => \N__37314\,
            I => \N__37311\
        );

    \I__7564\ : LocalMux
    port map (
            O => \N__37311\,
            I => \N__37308\
        );

    \I__7563\ : Span4Mux_v
    port map (
            O => \N__37308\,
            I => \N__37304\
        );

    \I__7562\ : InMux
    port map (
            O => \N__37307\,
            I => \N__37301\
        );

    \I__7561\ : Span4Mux_v
    port map (
            O => \N__37304\,
            I => \N__37298\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__37301\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__7559\ : Odrv4
    port map (
            O => \N__37298\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__7558\ : InMux
    port map (
            O => \N__37293\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\
        );

    \I__7557\ : InMux
    port map (
            O => \N__37290\,
            I => \N__37287\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__37287\,
            I => \N__37284\
        );

    \I__7555\ : Span4Mux_h
    port map (
            O => \N__37284\,
            I => \N__37280\
        );

    \I__7554\ : InMux
    port map (
            O => \N__37283\,
            I => \N__37277\
        );

    \I__7553\ : Span4Mux_v
    port map (
            O => \N__37280\,
            I => \N__37274\
        );

    \I__7552\ : LocalMux
    port map (
            O => \N__37277\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__7551\ : Odrv4
    port map (
            O => \N__37274\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__7550\ : InMux
    port map (
            O => \N__37269\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\
        );

    \I__7549\ : InMux
    port map (
            O => \N__37266\,
            I => \N__37263\
        );

    \I__7548\ : LocalMux
    port map (
            O => \N__37263\,
            I => \N__37260\
        );

    \I__7547\ : Span4Mux_h
    port map (
            O => \N__37260\,
            I => \N__37256\
        );

    \I__7546\ : InMux
    port map (
            O => \N__37259\,
            I => \N__37253\
        );

    \I__7545\ : Span4Mux_v
    port map (
            O => \N__37256\,
            I => \N__37250\
        );

    \I__7544\ : LocalMux
    port map (
            O => \N__37253\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__7543\ : Odrv4
    port map (
            O => \N__37250\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__7542\ : InMux
    port map (
            O => \N__37245\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\
        );

    \I__7541\ : InMux
    port map (
            O => \N__37242\,
            I => \N__37239\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__37239\,
            I => \N__37236\
        );

    \I__7539\ : Span4Mux_h
    port map (
            O => \N__37236\,
            I => \N__37232\
        );

    \I__7538\ : InMux
    port map (
            O => \N__37235\,
            I => \N__37229\
        );

    \I__7537\ : Span4Mux_v
    port map (
            O => \N__37232\,
            I => \N__37226\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__37229\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__7535\ : Odrv4
    port map (
            O => \N__37226\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__7534\ : InMux
    port map (
            O => \N__37221\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\
        );

    \I__7533\ : InMux
    port map (
            O => \N__37218\,
            I => \N__37214\
        );

    \I__7532\ : InMux
    port map (
            O => \N__37217\,
            I => \N__37211\
        );

    \I__7531\ : LocalMux
    port map (
            O => \N__37214\,
            I => \N__37208\
        );

    \I__7530\ : LocalMux
    port map (
            O => \N__37211\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__7529\ : Odrv4
    port map (
            O => \N__37208\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__7528\ : InMux
    port map (
            O => \N__37203\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__7527\ : InMux
    port map (
            O => \N__37200\,
            I => \N__37196\
        );

    \I__7526\ : InMux
    port map (
            O => \N__37199\,
            I => \N__37193\
        );

    \I__7525\ : LocalMux
    port map (
            O => \N__37196\,
            I => \N__37190\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__37193\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__7523\ : Odrv4
    port map (
            O => \N__37190\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__7522\ : InMux
    port map (
            O => \N__37185\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__7521\ : InMux
    port map (
            O => \N__37182\,
            I => \N__37178\
        );

    \I__7520\ : InMux
    port map (
            O => \N__37181\,
            I => \N__37175\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__37178\,
            I => \N__37172\
        );

    \I__7518\ : LocalMux
    port map (
            O => \N__37175\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__7517\ : Odrv4
    port map (
            O => \N__37172\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__7516\ : InMux
    port map (
            O => \N__37167\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__7515\ : InMux
    port map (
            O => \N__37164\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__7514\ : InMux
    port map (
            O => \N__37161\,
            I => \bfn_14_16_0_\
        );

    \I__7513\ : InMux
    port map (
            O => \N__37158\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__7512\ : InMux
    port map (
            O => \N__37155\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__7511\ : InMux
    port map (
            O => \N__37152\,
            I => \N__37148\
        );

    \I__7510\ : InMux
    port map (
            O => \N__37151\,
            I => \N__37145\
        );

    \I__7509\ : LocalMux
    port map (
            O => \N__37148\,
            I => \N__37142\
        );

    \I__7508\ : LocalMux
    port map (
            O => \N__37145\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__7507\ : Odrv4
    port map (
            O => \N__37142\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__7506\ : InMux
    port map (
            O => \N__37137\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\
        );

    \I__7505\ : InMux
    port map (
            O => \N__37134\,
            I => \N__37130\
        );

    \I__7504\ : InMux
    port map (
            O => \N__37133\,
            I => \N__37127\
        );

    \I__7503\ : LocalMux
    port map (
            O => \N__37130\,
            I => \N__37124\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__37127\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__7501\ : Odrv4
    port map (
            O => \N__37124\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__7500\ : InMux
    port map (
            O => \N__37119\,
            I => \N__37115\
        );

    \I__7499\ : InMux
    port map (
            O => \N__37118\,
            I => \N__37112\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__37115\,
            I => \N__37109\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__37112\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__7496\ : Odrv4
    port map (
            O => \N__37109\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__7495\ : InMux
    port map (
            O => \N__37104\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__7494\ : InMux
    port map (
            O => \N__37101\,
            I => \N__37097\
        );

    \I__7493\ : InMux
    port map (
            O => \N__37100\,
            I => \N__37094\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__37097\,
            I => \N__37091\
        );

    \I__7491\ : LocalMux
    port map (
            O => \N__37094\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__7490\ : Odrv4
    port map (
            O => \N__37091\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__7489\ : InMux
    port map (
            O => \N__37086\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__7488\ : InMux
    port map (
            O => \N__37083\,
            I => \N__37079\
        );

    \I__7487\ : InMux
    port map (
            O => \N__37082\,
            I => \N__37076\
        );

    \I__7486\ : LocalMux
    port map (
            O => \N__37079\,
            I => \N__37073\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__37076\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__7484\ : Odrv4
    port map (
            O => \N__37073\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__7483\ : InMux
    port map (
            O => \N__37068\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__7482\ : InMux
    port map (
            O => \N__37065\,
            I => \N__37061\
        );

    \I__7481\ : InMux
    port map (
            O => \N__37064\,
            I => \N__37058\
        );

    \I__7480\ : LocalMux
    port map (
            O => \N__37061\,
            I => \N__37055\
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__37058\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__7478\ : Odrv4
    port map (
            O => \N__37055\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__7477\ : InMux
    port map (
            O => \N__37050\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__7476\ : InMux
    port map (
            O => \N__37047\,
            I => \N__37043\
        );

    \I__7475\ : InMux
    port map (
            O => \N__37046\,
            I => \N__37040\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__37043\,
            I => \N__37037\
        );

    \I__7473\ : LocalMux
    port map (
            O => \N__37040\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__7472\ : Odrv4
    port map (
            O => \N__37037\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__7471\ : InMux
    port map (
            O => \N__37032\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__7470\ : InMux
    port map (
            O => \N__37029\,
            I => \N__37025\
        );

    \I__7469\ : InMux
    port map (
            O => \N__37028\,
            I => \N__37022\
        );

    \I__7468\ : LocalMux
    port map (
            O => \N__37025\,
            I => \N__37019\
        );

    \I__7467\ : LocalMux
    port map (
            O => \N__37022\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__7466\ : Odrv4
    port map (
            O => \N__37019\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__7465\ : InMux
    port map (
            O => \N__37014\,
            I => \bfn_14_15_0_\
        );

    \I__7464\ : InMux
    port map (
            O => \N__37011\,
            I => \N__37008\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__37008\,
            I => \N__37004\
        );

    \I__7462\ : InMux
    port map (
            O => \N__37007\,
            I => \N__37001\
        );

    \I__7461\ : Span4Mux_v
    port map (
            O => \N__37004\,
            I => \N__36998\
        );

    \I__7460\ : LocalMux
    port map (
            O => \N__37001\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__7459\ : Odrv4
    port map (
            O => \N__36998\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__7458\ : InMux
    port map (
            O => \N__36993\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__7457\ : InMux
    port map (
            O => \N__36990\,
            I => \N__36986\
        );

    \I__7456\ : InMux
    port map (
            O => \N__36989\,
            I => \N__36983\
        );

    \I__7455\ : LocalMux
    port map (
            O => \N__36986\,
            I => \N__36980\
        );

    \I__7454\ : LocalMux
    port map (
            O => \N__36983\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__7453\ : Odrv4
    port map (
            O => \N__36980\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__7452\ : InMux
    port map (
            O => \N__36975\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__7451\ : InMux
    port map (
            O => \N__36972\,
            I => \N__36968\
        );

    \I__7450\ : InMux
    port map (
            O => \N__36971\,
            I => \N__36965\
        );

    \I__7449\ : LocalMux
    port map (
            O => \N__36968\,
            I => \N__36962\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__36965\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__7447\ : Odrv4
    port map (
            O => \N__36962\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__7446\ : InMux
    port map (
            O => \N__36957\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__7445\ : InMux
    port map (
            O => \N__36954\,
            I => \N__36951\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__36951\,
            I => \current_shift_inst.control_input_axb_6\
        );

    \I__7443\ : InMux
    port map (
            O => \N__36948\,
            I => \N__36945\
        );

    \I__7442\ : LocalMux
    port map (
            O => \N__36945\,
            I => \N__36942\
        );

    \I__7441\ : Odrv4
    port map (
            O => \N__36942\,
            I => \current_shift_inst.control_input_axb_7\
        );

    \I__7440\ : InMux
    port map (
            O => \N__36939\,
            I => \N__36936\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__36936\,
            I => \N__36933\
        );

    \I__7438\ : Odrv4
    port map (
            O => \N__36933\,
            I => \current_shift_inst.control_input_axb_8\
        );

    \I__7437\ : InMux
    port map (
            O => \N__36930\,
            I => \N__36927\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__36927\,
            I => \current_shift_inst.control_input_axb_9\
        );

    \I__7435\ : InMux
    port map (
            O => \N__36924\,
            I => \N__36921\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__36921\,
            I => \current_shift_inst.control_input_axb_10\
        );

    \I__7433\ : CascadeMux
    port map (
            O => \N__36918\,
            I => \N__36915\
        );

    \I__7432\ : InMux
    port map (
            O => \N__36915\,
            I => \N__36910\
        );

    \I__7431\ : InMux
    port map (
            O => \N__36914\,
            I => \N__36907\
        );

    \I__7430\ : InMux
    port map (
            O => \N__36913\,
            I => \N__36904\
        );

    \I__7429\ : LocalMux
    port map (
            O => \N__36910\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__7428\ : LocalMux
    port map (
            O => \N__36907\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__7427\ : LocalMux
    port map (
            O => \N__36904\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__7426\ : CascadeMux
    port map (
            O => \N__36897\,
            I => \N__36894\
        );

    \I__7425\ : InMux
    port map (
            O => \N__36894\,
            I => \N__36891\
        );

    \I__7424\ : LocalMux
    port map (
            O => \N__36891\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\
        );

    \I__7423\ : InMux
    port map (
            O => \N__36888\,
            I => \N__36884\
        );

    \I__7422\ : InMux
    port map (
            O => \N__36887\,
            I => \N__36881\
        );

    \I__7421\ : LocalMux
    port map (
            O => \N__36884\,
            I => \N__36878\
        );

    \I__7420\ : LocalMux
    port map (
            O => \N__36881\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__7419\ : Odrv4
    port map (
            O => \N__36878\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__7418\ : InMux
    port map (
            O => \N__36873\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__7417\ : CascadeMux
    port map (
            O => \N__36870\,
            I => \N__36867\
        );

    \I__7416\ : InMux
    port map (
            O => \N__36867\,
            I => \N__36864\
        );

    \I__7415\ : LocalMux
    port map (
            O => \N__36864\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIQU8A2Z0Z_28\
        );

    \I__7414\ : InMux
    port map (
            O => \N__36861\,
            I => \N__36857\
        );

    \I__7413\ : InMux
    port map (
            O => \N__36860\,
            I => \N__36854\
        );

    \I__7412\ : LocalMux
    port map (
            O => \N__36857\,
            I => \N__36851\
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__36854\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__7410\ : Odrv4
    port map (
            O => \N__36851\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__7409\ : InMux
    port map (
            O => \N__36846\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__7408\ : CascadeMux
    port map (
            O => \N__36843\,
            I => \current_shift_inst.control_input_axb_0_cascade_\
        );

    \I__7407\ : InMux
    port map (
            O => \N__36840\,
            I => \N__36837\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__36837\,
            I => \N__36833\
        );

    \I__7405\ : InMux
    port map (
            O => \N__36836\,
            I => \N__36830\
        );

    \I__7404\ : Span4Mux_h
    port map (
            O => \N__36833\,
            I => \N__36827\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__36830\,
            I => \N__36824\
        );

    \I__7402\ : Span4Mux_h
    port map (
            O => \N__36827\,
            I => \N__36821\
        );

    \I__7401\ : Span4Mux_h
    port map (
            O => \N__36824\,
            I => \N__36818\
        );

    \I__7400\ : Odrv4
    port map (
            O => \N__36821\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__7399\ : Odrv4
    port map (
            O => \N__36818\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__7398\ : InMux
    port map (
            O => \N__36813\,
            I => \N__36810\
        );

    \I__7397\ : LocalMux
    port map (
            O => \N__36810\,
            I => \N__36807\
        );

    \I__7396\ : Odrv4
    port map (
            O => \N__36807\,
            I => \current_shift_inst.elapsed_time_ns_s1_fast_31\
        );

    \I__7395\ : InMux
    port map (
            O => \N__36804\,
            I => \N__36801\
        );

    \I__7394\ : LocalMux
    port map (
            O => \N__36801\,
            I => \current_shift_inst.control_input_axb_1\
        );

    \I__7393\ : InMux
    port map (
            O => \N__36798\,
            I => \N__36795\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__36795\,
            I => \current_shift_inst.control_input_axb_12\
        );

    \I__7391\ : InMux
    port map (
            O => \N__36792\,
            I => \N__36788\
        );

    \I__7390\ : CascadeMux
    port map (
            O => \N__36791\,
            I => \N__36784\
        );

    \I__7389\ : LocalMux
    port map (
            O => \N__36788\,
            I => \N__36781\
        );

    \I__7388\ : InMux
    port map (
            O => \N__36787\,
            I => \N__36778\
        );

    \I__7387\ : InMux
    port map (
            O => \N__36784\,
            I => \N__36775\
        );

    \I__7386\ : Odrv4
    port map (
            O => \N__36781\,
            I => \current_shift_inst.N_1460_i\
        );

    \I__7385\ : LocalMux
    port map (
            O => \N__36778\,
            I => \current_shift_inst.N_1460_i\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__36775\,
            I => \current_shift_inst.N_1460_i\
        );

    \I__7383\ : InMux
    port map (
            O => \N__36768\,
            I => \N__36765\
        );

    \I__7382\ : LocalMux
    port map (
            O => \N__36765\,
            I => \current_shift_inst.control_input_axb_2\
        );

    \I__7381\ : InMux
    port map (
            O => \N__36762\,
            I => \N__36759\
        );

    \I__7380\ : LocalMux
    port map (
            O => \N__36759\,
            I => \current_shift_inst.control_input_axb_3\
        );

    \I__7379\ : InMux
    port map (
            O => \N__36756\,
            I => \N__36753\
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__36753\,
            I => \current_shift_inst.control_input_axb_4\
        );

    \I__7377\ : InMux
    port map (
            O => \N__36750\,
            I => \N__36747\
        );

    \I__7376\ : LocalMux
    port map (
            O => \N__36747\,
            I => \current_shift_inst.control_input_axb_5\
        );

    \I__7375\ : InMux
    port map (
            O => \N__36744\,
            I => \N__36741\
        );

    \I__7374\ : LocalMux
    port map (
            O => \N__36741\,
            I => \current_shift_inst.control_input_axb_0\
        );

    \I__7373\ : CascadeMux
    port map (
            O => \N__36738\,
            I => \N__36734\
        );

    \I__7372\ : CascadeMux
    port map (
            O => \N__36737\,
            I => \N__36731\
        );

    \I__7371\ : InMux
    port map (
            O => \N__36734\,
            I => \N__36725\
        );

    \I__7370\ : InMux
    port map (
            O => \N__36731\,
            I => \N__36725\
        );

    \I__7369\ : InMux
    port map (
            O => \N__36730\,
            I => \N__36722\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__36725\,
            I => \N__36719\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__36722\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__7366\ : Odrv4
    port map (
            O => \N__36719\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__7365\ : InMux
    port map (
            O => \N__36714\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__7364\ : InMux
    port map (
            O => \N__36711\,
            I => \N__36704\
        );

    \I__7363\ : InMux
    port map (
            O => \N__36710\,
            I => \N__36704\
        );

    \I__7362\ : InMux
    port map (
            O => \N__36709\,
            I => \N__36701\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__36704\,
            I => \N__36698\
        );

    \I__7360\ : LocalMux
    port map (
            O => \N__36701\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__7359\ : Odrv4
    port map (
            O => \N__36698\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__7358\ : InMux
    port map (
            O => \N__36693\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__7357\ : InMux
    port map (
            O => \N__36690\,
            I => \N__36686\
        );

    \I__7356\ : InMux
    port map (
            O => \N__36689\,
            I => \N__36683\
        );

    \I__7355\ : LocalMux
    port map (
            O => \N__36686\,
            I => \N__36680\
        );

    \I__7354\ : LocalMux
    port map (
            O => \N__36683\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__7353\ : Odrv4
    port map (
            O => \N__36680\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__7352\ : InMux
    port map (
            O => \N__36675\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__7351\ : InMux
    port map (
            O => \N__36672\,
            I => \N__36658\
        );

    \I__7350\ : InMux
    port map (
            O => \N__36671\,
            I => \N__36658\
        );

    \I__7349\ : InMux
    port map (
            O => \N__36670\,
            I => \N__36637\
        );

    \I__7348\ : InMux
    port map (
            O => \N__36669\,
            I => \N__36637\
        );

    \I__7347\ : InMux
    port map (
            O => \N__36668\,
            I => \N__36637\
        );

    \I__7346\ : InMux
    port map (
            O => \N__36667\,
            I => \N__36637\
        );

    \I__7345\ : InMux
    port map (
            O => \N__36666\,
            I => \N__36620\
        );

    \I__7344\ : InMux
    port map (
            O => \N__36665\,
            I => \N__36620\
        );

    \I__7343\ : InMux
    port map (
            O => \N__36664\,
            I => \N__36620\
        );

    \I__7342\ : InMux
    port map (
            O => \N__36663\,
            I => \N__36620\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__36658\,
            I => \N__36617\
        );

    \I__7340\ : InMux
    port map (
            O => \N__36657\,
            I => \N__36608\
        );

    \I__7339\ : InMux
    port map (
            O => \N__36656\,
            I => \N__36608\
        );

    \I__7338\ : InMux
    port map (
            O => \N__36655\,
            I => \N__36608\
        );

    \I__7337\ : InMux
    port map (
            O => \N__36654\,
            I => \N__36608\
        );

    \I__7336\ : InMux
    port map (
            O => \N__36653\,
            I => \N__36599\
        );

    \I__7335\ : InMux
    port map (
            O => \N__36652\,
            I => \N__36599\
        );

    \I__7334\ : InMux
    port map (
            O => \N__36651\,
            I => \N__36599\
        );

    \I__7333\ : InMux
    port map (
            O => \N__36650\,
            I => \N__36599\
        );

    \I__7332\ : InMux
    port map (
            O => \N__36649\,
            I => \N__36590\
        );

    \I__7331\ : InMux
    port map (
            O => \N__36648\,
            I => \N__36590\
        );

    \I__7330\ : InMux
    port map (
            O => \N__36647\,
            I => \N__36590\
        );

    \I__7329\ : InMux
    port map (
            O => \N__36646\,
            I => \N__36590\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__36637\,
            I => \N__36587\
        );

    \I__7327\ : InMux
    port map (
            O => \N__36636\,
            I => \N__36578\
        );

    \I__7326\ : InMux
    port map (
            O => \N__36635\,
            I => \N__36578\
        );

    \I__7325\ : InMux
    port map (
            O => \N__36634\,
            I => \N__36578\
        );

    \I__7324\ : InMux
    port map (
            O => \N__36633\,
            I => \N__36578\
        );

    \I__7323\ : InMux
    port map (
            O => \N__36632\,
            I => \N__36569\
        );

    \I__7322\ : InMux
    port map (
            O => \N__36631\,
            I => \N__36569\
        );

    \I__7321\ : InMux
    port map (
            O => \N__36630\,
            I => \N__36569\
        );

    \I__7320\ : InMux
    port map (
            O => \N__36629\,
            I => \N__36569\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__36620\,
            I => \N__36558\
        );

    \I__7318\ : Span4Mux_h
    port map (
            O => \N__36617\,
            I => \N__36558\
        );

    \I__7317\ : LocalMux
    port map (
            O => \N__36608\,
            I => \N__36558\
        );

    \I__7316\ : LocalMux
    port map (
            O => \N__36599\,
            I => \N__36558\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__36590\,
            I => \N__36558\
        );

    \I__7314\ : Odrv4
    port map (
            O => \N__36587\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__36578\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__36569\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__7311\ : Odrv4
    port map (
            O => \N__36558\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__7310\ : InMux
    port map (
            O => \N__36549\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__7309\ : CascadeMux
    port map (
            O => \N__36546\,
            I => \N__36543\
        );

    \I__7308\ : InMux
    port map (
            O => \N__36543\,
            I => \N__36539\
        );

    \I__7307\ : InMux
    port map (
            O => \N__36542\,
            I => \N__36536\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__36539\,
            I => \N__36533\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__36536\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__7304\ : Odrv4
    port map (
            O => \N__36533\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__7303\ : CEMux
    port map (
            O => \N__36528\,
            I => \N__36525\
        );

    \I__7302\ : LocalMux
    port map (
            O => \N__36525\,
            I => \N__36520\
        );

    \I__7301\ : CEMux
    port map (
            O => \N__36524\,
            I => \N__36517\
        );

    \I__7300\ : CEMux
    port map (
            O => \N__36523\,
            I => \N__36513\
        );

    \I__7299\ : Span4Mux_v
    port map (
            O => \N__36520\,
            I => \N__36508\
        );

    \I__7298\ : LocalMux
    port map (
            O => \N__36517\,
            I => \N__36508\
        );

    \I__7297\ : CEMux
    port map (
            O => \N__36516\,
            I => \N__36505\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__36513\,
            I => \N__36502\
        );

    \I__7295\ : Span4Mux_v
    port map (
            O => \N__36508\,
            I => \N__36497\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__36505\,
            I => \N__36497\
        );

    \I__7293\ : Span4Mux_v
    port map (
            O => \N__36502\,
            I => \N__36494\
        );

    \I__7292\ : Span4Mux_v
    port map (
            O => \N__36497\,
            I => \N__36489\
        );

    \I__7291\ : Span4Mux_s1_v
    port map (
            O => \N__36494\,
            I => \N__36489\
        );

    \I__7290\ : Odrv4
    port map (
            O => \N__36489\,
            I => \current_shift_inst.timer_s1.N_167_i\
        );

    \I__7289\ : CascadeMux
    port map (
            O => \N__36486\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1_cascade_\
        );

    \I__7288\ : CascadeMux
    port map (
            O => \N__36483\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\
        );

    \I__7287\ : CascadeMux
    port map (
            O => \N__36480\,
            I => \N__36477\
        );

    \I__7286\ : InMux
    port map (
            O => \N__36477\,
            I => \N__36474\
        );

    \I__7285\ : LocalMux
    port map (
            O => \N__36474\,
            I => \N__36470\
        );

    \I__7284\ : InMux
    port map (
            O => \N__36473\,
            I => \N__36466\
        );

    \I__7283\ : Span4Mux_h
    port map (
            O => \N__36470\,
            I => \N__36463\
        );

    \I__7282\ : InMux
    port map (
            O => \N__36469\,
            I => \N__36460\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__36466\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__7280\ : Odrv4
    port map (
            O => \N__36463\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__7279\ : LocalMux
    port map (
            O => \N__36460\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__7278\ : InMux
    port map (
            O => \N__36453\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__7277\ : InMux
    port map (
            O => \N__36450\,
            I => \N__36444\
        );

    \I__7276\ : InMux
    port map (
            O => \N__36449\,
            I => \N__36444\
        );

    \I__7275\ : LocalMux
    port map (
            O => \N__36444\,
            I => \N__36440\
        );

    \I__7274\ : InMux
    port map (
            O => \N__36443\,
            I => \N__36437\
        );

    \I__7273\ : Span4Mux_v
    port map (
            O => \N__36440\,
            I => \N__36434\
        );

    \I__7272\ : LocalMux
    port map (
            O => \N__36437\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__7271\ : Odrv4
    port map (
            O => \N__36434\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__7270\ : InMux
    port map (
            O => \N__36429\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__7269\ : InMux
    port map (
            O => \N__36426\,
            I => \N__36419\
        );

    \I__7268\ : InMux
    port map (
            O => \N__36425\,
            I => \N__36419\
        );

    \I__7267\ : InMux
    port map (
            O => \N__36424\,
            I => \N__36416\
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__36419\,
            I => \N__36413\
        );

    \I__7265\ : LocalMux
    port map (
            O => \N__36416\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__7264\ : Odrv4
    port map (
            O => \N__36413\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__7263\ : InMux
    port map (
            O => \N__36408\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__7262\ : CascadeMux
    port map (
            O => \N__36405\,
            I => \N__36401\
        );

    \I__7261\ : CascadeMux
    port map (
            O => \N__36404\,
            I => \N__36398\
        );

    \I__7260\ : InMux
    port map (
            O => \N__36401\,
            I => \N__36393\
        );

    \I__7259\ : InMux
    port map (
            O => \N__36398\,
            I => \N__36393\
        );

    \I__7258\ : LocalMux
    port map (
            O => \N__36393\,
            I => \N__36389\
        );

    \I__7257\ : InMux
    port map (
            O => \N__36392\,
            I => \N__36386\
        );

    \I__7256\ : Span4Mux_h
    port map (
            O => \N__36389\,
            I => \N__36383\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__36386\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__7254\ : Odrv4
    port map (
            O => \N__36383\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__7253\ : InMux
    port map (
            O => \N__36378\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__7252\ : CascadeMux
    port map (
            O => \N__36375\,
            I => \N__36371\
        );

    \I__7251\ : CascadeMux
    port map (
            O => \N__36374\,
            I => \N__36368\
        );

    \I__7250\ : InMux
    port map (
            O => \N__36371\,
            I => \N__36362\
        );

    \I__7249\ : InMux
    port map (
            O => \N__36368\,
            I => \N__36362\
        );

    \I__7248\ : InMux
    port map (
            O => \N__36367\,
            I => \N__36359\
        );

    \I__7247\ : LocalMux
    port map (
            O => \N__36362\,
            I => \N__36356\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__36359\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__7245\ : Odrv4
    port map (
            O => \N__36356\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__7244\ : InMux
    port map (
            O => \N__36351\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__7243\ : InMux
    port map (
            O => \N__36348\,
            I => \N__36341\
        );

    \I__7242\ : InMux
    port map (
            O => \N__36347\,
            I => \N__36341\
        );

    \I__7241\ : InMux
    port map (
            O => \N__36346\,
            I => \N__36338\
        );

    \I__7240\ : LocalMux
    port map (
            O => \N__36341\,
            I => \N__36335\
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__36338\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__7238\ : Odrv4
    port map (
            O => \N__36335\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__7237\ : InMux
    port map (
            O => \N__36330\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__7236\ : CascadeMux
    port map (
            O => \N__36327\,
            I => \N__36323\
        );

    \I__7235\ : InMux
    port map (
            O => \N__36326\,
            I => \N__36320\
        );

    \I__7234\ : InMux
    port map (
            O => \N__36323\,
            I => \N__36316\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__36320\,
            I => \N__36313\
        );

    \I__7232\ : InMux
    port map (
            O => \N__36319\,
            I => \N__36310\
        );

    \I__7231\ : LocalMux
    port map (
            O => \N__36316\,
            I => \N__36305\
        );

    \I__7230\ : Span4Mux_h
    port map (
            O => \N__36313\,
            I => \N__36305\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__36310\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__7228\ : Odrv4
    port map (
            O => \N__36305\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__7227\ : InMux
    port map (
            O => \N__36300\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__7226\ : InMux
    port map (
            O => \N__36297\,
            I => \N__36294\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__36294\,
            I => \N__36289\
        );

    \I__7224\ : CascadeMux
    port map (
            O => \N__36293\,
            I => \N__36286\
        );

    \I__7223\ : InMux
    port map (
            O => \N__36292\,
            I => \N__36283\
        );

    \I__7222\ : Span4Mux_h
    port map (
            O => \N__36289\,
            I => \N__36280\
        );

    \I__7221\ : InMux
    port map (
            O => \N__36286\,
            I => \N__36277\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__36283\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__7219\ : Odrv4
    port map (
            O => \N__36280\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__7218\ : LocalMux
    port map (
            O => \N__36277\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__7217\ : InMux
    port map (
            O => \N__36270\,
            I => \bfn_14_8_0_\
        );

    \I__7216\ : CascadeMux
    port map (
            O => \N__36267\,
            I => \N__36264\
        );

    \I__7215\ : InMux
    port map (
            O => \N__36264\,
            I => \N__36261\
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__36261\,
            I => \N__36257\
        );

    \I__7213\ : InMux
    port map (
            O => \N__36260\,
            I => \N__36253\
        );

    \I__7212\ : Span4Mux_h
    port map (
            O => \N__36257\,
            I => \N__36250\
        );

    \I__7211\ : InMux
    port map (
            O => \N__36256\,
            I => \N__36247\
        );

    \I__7210\ : LocalMux
    port map (
            O => \N__36253\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__7209\ : Odrv4
    port map (
            O => \N__36250\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__36247\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__7207\ : InMux
    port map (
            O => \N__36240\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__7206\ : CascadeMux
    port map (
            O => \N__36237\,
            I => \N__36234\
        );

    \I__7205\ : InMux
    port map (
            O => \N__36234\,
            I => \N__36231\
        );

    \I__7204\ : LocalMux
    port map (
            O => \N__36231\,
            I => \N__36227\
        );

    \I__7203\ : InMux
    port map (
            O => \N__36230\,
            I => \N__36223\
        );

    \I__7202\ : Span4Mux_h
    port map (
            O => \N__36227\,
            I => \N__36220\
        );

    \I__7201\ : InMux
    port map (
            O => \N__36226\,
            I => \N__36217\
        );

    \I__7200\ : LocalMux
    port map (
            O => \N__36223\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__7199\ : Odrv4
    port map (
            O => \N__36220\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__36217\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__7197\ : InMux
    port map (
            O => \N__36210\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__7196\ : InMux
    port map (
            O => \N__36207\,
            I => \N__36201\
        );

    \I__7195\ : InMux
    port map (
            O => \N__36206\,
            I => \N__36201\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__36201\,
            I => \N__36197\
        );

    \I__7193\ : InMux
    port map (
            O => \N__36200\,
            I => \N__36194\
        );

    \I__7192\ : Span4Mux_v
    port map (
            O => \N__36197\,
            I => \N__36191\
        );

    \I__7191\ : LocalMux
    port map (
            O => \N__36194\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__7190\ : Odrv4
    port map (
            O => \N__36191\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__7189\ : InMux
    port map (
            O => \N__36186\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__7188\ : InMux
    port map (
            O => \N__36183\,
            I => \N__36176\
        );

    \I__7187\ : InMux
    port map (
            O => \N__36182\,
            I => \N__36176\
        );

    \I__7186\ : InMux
    port map (
            O => \N__36181\,
            I => \N__36173\
        );

    \I__7185\ : LocalMux
    port map (
            O => \N__36176\,
            I => \N__36170\
        );

    \I__7184\ : LocalMux
    port map (
            O => \N__36173\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__7183\ : Odrv4
    port map (
            O => \N__36170\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__7182\ : InMux
    port map (
            O => \N__36165\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__7181\ : CascadeMux
    port map (
            O => \N__36162\,
            I => \N__36158\
        );

    \I__7180\ : CascadeMux
    port map (
            O => \N__36161\,
            I => \N__36155\
        );

    \I__7179\ : InMux
    port map (
            O => \N__36158\,
            I => \N__36150\
        );

    \I__7178\ : InMux
    port map (
            O => \N__36155\,
            I => \N__36150\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__36150\,
            I => \N__36146\
        );

    \I__7176\ : InMux
    port map (
            O => \N__36149\,
            I => \N__36143\
        );

    \I__7175\ : Span4Mux_h
    port map (
            O => \N__36146\,
            I => \N__36140\
        );

    \I__7174\ : LocalMux
    port map (
            O => \N__36143\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__7173\ : Odrv4
    port map (
            O => \N__36140\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__7172\ : InMux
    port map (
            O => \N__36135\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__7171\ : CascadeMux
    port map (
            O => \N__36132\,
            I => \N__36128\
        );

    \I__7170\ : CascadeMux
    port map (
            O => \N__36131\,
            I => \N__36125\
        );

    \I__7169\ : InMux
    port map (
            O => \N__36128\,
            I => \N__36119\
        );

    \I__7168\ : InMux
    port map (
            O => \N__36125\,
            I => \N__36119\
        );

    \I__7167\ : InMux
    port map (
            O => \N__36124\,
            I => \N__36116\
        );

    \I__7166\ : LocalMux
    port map (
            O => \N__36119\,
            I => \N__36113\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__36116\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__7164\ : Odrv4
    port map (
            O => \N__36113\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__7163\ : InMux
    port map (
            O => \N__36108\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__7162\ : InMux
    port map (
            O => \N__36105\,
            I => \N__36098\
        );

    \I__7161\ : InMux
    port map (
            O => \N__36104\,
            I => \N__36098\
        );

    \I__7160\ : InMux
    port map (
            O => \N__36103\,
            I => \N__36095\
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__36098\,
            I => \N__36092\
        );

    \I__7158\ : LocalMux
    port map (
            O => \N__36095\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__7157\ : Odrv4
    port map (
            O => \N__36092\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__7156\ : InMux
    port map (
            O => \N__36087\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__7155\ : CascadeMux
    port map (
            O => \N__36084\,
            I => \N__36081\
        );

    \I__7154\ : InMux
    port map (
            O => \N__36081\,
            I => \N__36077\
        );

    \I__7153\ : InMux
    port map (
            O => \N__36080\,
            I => \N__36074\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__36077\,
            I => \N__36068\
        );

    \I__7151\ : LocalMux
    port map (
            O => \N__36074\,
            I => \N__36068\
        );

    \I__7150\ : InMux
    port map (
            O => \N__36073\,
            I => \N__36065\
        );

    \I__7149\ : Span4Mux_h
    port map (
            O => \N__36068\,
            I => \N__36062\
        );

    \I__7148\ : LocalMux
    port map (
            O => \N__36065\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__7147\ : Odrv4
    port map (
            O => \N__36062\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__7146\ : InMux
    port map (
            O => \N__36057\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__7145\ : CascadeMux
    port map (
            O => \N__36054\,
            I => \N__36051\
        );

    \I__7144\ : InMux
    port map (
            O => \N__36051\,
            I => \N__36046\
        );

    \I__7143\ : CascadeMux
    port map (
            O => \N__36050\,
            I => \N__36043\
        );

    \I__7142\ : InMux
    port map (
            O => \N__36049\,
            I => \N__36040\
        );

    \I__7141\ : LocalMux
    port map (
            O => \N__36046\,
            I => \N__36037\
        );

    \I__7140\ : InMux
    port map (
            O => \N__36043\,
            I => \N__36034\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__36040\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__7138\ : Odrv4
    port map (
            O => \N__36037\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__7137\ : LocalMux
    port map (
            O => \N__36034\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__7136\ : InMux
    port map (
            O => \N__36027\,
            I => \bfn_14_7_0_\
        );

    \I__7135\ : InMux
    port map (
            O => \N__36024\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__7134\ : CascadeMux
    port map (
            O => \N__36021\,
            I => \N__36017\
        );

    \I__7133\ : CascadeMux
    port map (
            O => \N__36020\,
            I => \N__36014\
        );

    \I__7132\ : InMux
    port map (
            O => \N__36017\,
            I => \N__36008\
        );

    \I__7131\ : InMux
    port map (
            O => \N__36014\,
            I => \N__36008\
        );

    \I__7130\ : InMux
    port map (
            O => \N__36013\,
            I => \N__36005\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__36008\,
            I => \N__36002\
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__36005\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__7127\ : Odrv4
    port map (
            O => \N__36002\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__7126\ : InMux
    port map (
            O => \N__35997\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__7125\ : CascadeMux
    port map (
            O => \N__35994\,
            I => \N__35991\
        );

    \I__7124\ : InMux
    port map (
            O => \N__35991\,
            I => \N__35987\
        );

    \I__7123\ : InMux
    port map (
            O => \N__35990\,
            I => \N__35983\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__35987\,
            I => \N__35980\
        );

    \I__7121\ : InMux
    port map (
            O => \N__35986\,
            I => \N__35977\
        );

    \I__7120\ : LocalMux
    port map (
            O => \N__35983\,
            I => \N__35974\
        );

    \I__7119\ : Span4Mux_v
    port map (
            O => \N__35980\,
            I => \N__35971\
        );

    \I__7118\ : LocalMux
    port map (
            O => \N__35977\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__7117\ : Odrv4
    port map (
            O => \N__35974\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__7116\ : Odrv4
    port map (
            O => \N__35971\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__7115\ : InMux
    port map (
            O => \N__35964\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__7114\ : InMux
    port map (
            O => \N__35961\,
            I => \N__35954\
        );

    \I__7113\ : InMux
    port map (
            O => \N__35960\,
            I => \N__35954\
        );

    \I__7112\ : InMux
    port map (
            O => \N__35959\,
            I => \N__35951\
        );

    \I__7111\ : LocalMux
    port map (
            O => \N__35954\,
            I => \N__35948\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__35951\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__7109\ : Odrv4
    port map (
            O => \N__35948\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__7108\ : InMux
    port map (
            O => \N__35943\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__7107\ : CascadeMux
    port map (
            O => \N__35940\,
            I => \N__35936\
        );

    \I__7106\ : CascadeMux
    port map (
            O => \N__35939\,
            I => \N__35933\
        );

    \I__7105\ : InMux
    port map (
            O => \N__35936\,
            I => \N__35927\
        );

    \I__7104\ : InMux
    port map (
            O => \N__35933\,
            I => \N__35927\
        );

    \I__7103\ : InMux
    port map (
            O => \N__35932\,
            I => \N__35924\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__35927\,
            I => \N__35921\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__35924\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__7100\ : Odrv4
    port map (
            O => \N__35921\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__7099\ : InMux
    port map (
            O => \N__35916\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__7098\ : CascadeMux
    port map (
            O => \N__35913\,
            I => \N__35909\
        );

    \I__7097\ : CascadeMux
    port map (
            O => \N__35912\,
            I => \N__35906\
        );

    \I__7096\ : InMux
    port map (
            O => \N__35909\,
            I => \N__35901\
        );

    \I__7095\ : InMux
    port map (
            O => \N__35906\,
            I => \N__35901\
        );

    \I__7094\ : LocalMux
    port map (
            O => \N__35901\,
            I => \N__35897\
        );

    \I__7093\ : InMux
    port map (
            O => \N__35900\,
            I => \N__35894\
        );

    \I__7092\ : Span4Mux_h
    port map (
            O => \N__35897\,
            I => \N__35891\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__35894\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__7090\ : Odrv4
    port map (
            O => \N__35891\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__7089\ : InMux
    port map (
            O => \N__35886\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__7088\ : CascadeMux
    port map (
            O => \N__35883\,
            I => \N__35879\
        );

    \I__7087\ : InMux
    port map (
            O => \N__35882\,
            I => \N__35876\
        );

    \I__7086\ : InMux
    port map (
            O => \N__35879\,
            I => \N__35872\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__35876\,
            I => \N__35869\
        );

    \I__7084\ : InMux
    port map (
            O => \N__35875\,
            I => \N__35866\
        );

    \I__7083\ : LocalMux
    port map (
            O => \N__35872\,
            I => \N__35861\
        );

    \I__7082\ : Span4Mux_h
    port map (
            O => \N__35869\,
            I => \N__35861\
        );

    \I__7081\ : LocalMux
    port map (
            O => \N__35866\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__7080\ : Odrv4
    port map (
            O => \N__35861\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__7079\ : InMux
    port map (
            O => \N__35856\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__7078\ : CascadeMux
    port map (
            O => \N__35853\,
            I => \N__35850\
        );

    \I__7077\ : InMux
    port map (
            O => \N__35850\,
            I => \N__35846\
        );

    \I__7076\ : InMux
    port map (
            O => \N__35849\,
            I => \N__35842\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__35846\,
            I => \N__35839\
        );

    \I__7074\ : InMux
    port map (
            O => \N__35845\,
            I => \N__35836\
        );

    \I__7073\ : LocalMux
    port map (
            O => \N__35842\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__7072\ : Odrv4
    port map (
            O => \N__35839\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__7071\ : LocalMux
    port map (
            O => \N__35836\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__7070\ : InMux
    port map (
            O => \N__35829\,
            I => \bfn_14_6_0_\
        );

    \I__7069\ : IoInMux
    port map (
            O => \N__35826\,
            I => \N__35823\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__35823\,
            I => \N__35820\
        );

    \I__7067\ : Span12Mux_s1_v
    port map (
            O => \N__35820\,
            I => \N__35817\
        );

    \I__7066\ : Odrv12
    port map (
            O => \N__35817\,
            I => \current_shift_inst.timer_s1.N_166_i\
        );

    \I__7065\ : InMux
    port map (
            O => \N__35814\,
            I => \N__35810\
        );

    \I__7064\ : InMux
    port map (
            O => \N__35813\,
            I => \N__35807\
        );

    \I__7063\ : LocalMux
    port map (
            O => \N__35810\,
            I => \N__35801\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__35807\,
            I => \N__35801\
        );

    \I__7061\ : InMux
    port map (
            O => \N__35806\,
            I => \N__35797\
        );

    \I__7060\ : Span12Mux_s10_v
    port map (
            O => \N__35801\,
            I => \N__35794\
        );

    \I__7059\ : InMux
    port map (
            O => \N__35800\,
            I => \N__35791\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__35797\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7057\ : Odrv12
    port map (
            O => \N__35794\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7056\ : LocalMux
    port map (
            O => \N__35791\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7055\ : InMux
    port map (
            O => \N__35784\,
            I => \N__35781\
        );

    \I__7054\ : LocalMux
    port map (
            O => \N__35781\,
            I => \N__35776\
        );

    \I__7053\ : InMux
    port map (
            O => \N__35780\,
            I => \N__35770\
        );

    \I__7052\ : InMux
    port map (
            O => \N__35779\,
            I => \N__35770\
        );

    \I__7051\ : Span12Mux_s11_v
    port map (
            O => \N__35776\,
            I => \N__35767\
        );

    \I__7050\ : InMux
    port map (
            O => \N__35775\,
            I => \N__35764\
        );

    \I__7049\ : LocalMux
    port map (
            O => \N__35770\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7048\ : Odrv12
    port map (
            O => \N__35767\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7047\ : LocalMux
    port map (
            O => \N__35764\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7046\ : InMux
    port map (
            O => \N__35757\,
            I => \N__35754\
        );

    \I__7045\ : LocalMux
    port map (
            O => \N__35754\,
            I => \N__35751\
        );

    \I__7044\ : Span12Mux_s9_v
    port map (
            O => \N__35751\,
            I => \N__35745\
        );

    \I__7043\ : InMux
    port map (
            O => \N__35750\,
            I => \N__35740\
        );

    \I__7042\ : InMux
    port map (
            O => \N__35749\,
            I => \N__35740\
        );

    \I__7041\ : InMux
    port map (
            O => \N__35748\,
            I => \N__35737\
        );

    \I__7040\ : Span12Mux_v
    port map (
            O => \N__35745\,
            I => \N__35734\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__35740\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__7038\ : LocalMux
    port map (
            O => \N__35737\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__7037\ : Odrv12
    port map (
            O => \N__35734\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__7036\ : IoInMux
    port map (
            O => \N__35727\,
            I => \N__35724\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__35724\,
            I => \N__35720\
        );

    \I__7034\ : InMux
    port map (
            O => \N__35723\,
            I => \N__35717\
        );

    \I__7033\ : Span12Mux_s5_v
    port map (
            O => \N__35720\,
            I => \N__35713\
        );

    \I__7032\ : LocalMux
    port map (
            O => \N__35717\,
            I => \N__35710\
        );

    \I__7031\ : InMux
    port map (
            O => \N__35716\,
            I => \N__35707\
        );

    \I__7030\ : Odrv12
    port map (
            O => \N__35713\,
            I => s1_phy_c
        );

    \I__7029\ : Odrv4
    port map (
            O => \N__35710\,
            I => s1_phy_c
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__35707\,
            I => s1_phy_c
        );

    \I__7027\ : IoInMux
    port map (
            O => \N__35700\,
            I => \N__35697\
        );

    \I__7026\ : LocalMux
    port map (
            O => \N__35697\,
            I => \N__35694\
        );

    \I__7025\ : Span4Mux_s2_v
    port map (
            O => \N__35694\,
            I => \N__35691\
        );

    \I__7024\ : Span4Mux_h
    port map (
            O => \N__35691\,
            I => \N__35687\
        );

    \I__7023\ : InMux
    port map (
            O => \N__35690\,
            I => \N__35684\
        );

    \I__7022\ : Odrv4
    port map (
            O => \N__35687\,
            I => \T23_c\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__35684\,
            I => \T23_c\
        );

    \I__7020\ : InMux
    port map (
            O => \N__35679\,
            I => \N__35673\
        );

    \I__7019\ : InMux
    port map (
            O => \N__35678\,
            I => \N__35673\
        );

    \I__7018\ : LocalMux
    port map (
            O => \N__35673\,
            I => \N__35670\
        );

    \I__7017\ : Span4Mux_v
    port map (
            O => \N__35670\,
            I => \N__35665\
        );

    \I__7016\ : InMux
    port map (
            O => \N__35669\,
            I => \N__35662\
        );

    \I__7015\ : InMux
    port map (
            O => \N__35668\,
            I => \N__35659\
        );

    \I__7014\ : Odrv4
    port map (
            O => \N__35665\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__35662\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__7012\ : LocalMux
    port map (
            O => \N__35659\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__7011\ : CascadeMux
    port map (
            O => \N__35652\,
            I => \N__35646\
        );

    \I__7010\ : InMux
    port map (
            O => \N__35651\,
            I => \N__35642\
        );

    \I__7009\ : InMux
    port map (
            O => \N__35650\,
            I => \N__35639\
        );

    \I__7008\ : InMux
    port map (
            O => \N__35649\,
            I => \N__35636\
        );

    \I__7007\ : InMux
    port map (
            O => \N__35646\,
            I => \N__35633\
        );

    \I__7006\ : InMux
    port map (
            O => \N__35645\,
            I => \N__35630\
        );

    \I__7005\ : LocalMux
    port map (
            O => \N__35642\,
            I => \N__35625\
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__35639\,
            I => \N__35616\
        );

    \I__7003\ : LocalMux
    port map (
            O => \N__35636\,
            I => \N__35616\
        );

    \I__7002\ : LocalMux
    port map (
            O => \N__35633\,
            I => \N__35616\
        );

    \I__7001\ : LocalMux
    port map (
            O => \N__35630\,
            I => \N__35616\
        );

    \I__7000\ : InMux
    port map (
            O => \N__35629\,
            I => \N__35612\
        );

    \I__6999\ : InMux
    port map (
            O => \N__35628\,
            I => \N__35609\
        );

    \I__6998\ : Span4Mux_v
    port map (
            O => \N__35625\,
            I => \N__35604\
        );

    \I__6997\ : Span4Mux_v
    port map (
            O => \N__35616\,
            I => \N__35604\
        );

    \I__6996\ : InMux
    port map (
            O => \N__35615\,
            I => \N__35601\
        );

    \I__6995\ : LocalMux
    port map (
            O => \N__35612\,
            I => state_3
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__35609\,
            I => state_3
        );

    \I__6993\ : Odrv4
    port map (
            O => \N__35604\,
            I => state_3
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__35601\,
            I => state_3
        );

    \I__6991\ : IoInMux
    port map (
            O => \N__35592\,
            I => \N__35589\
        );

    \I__6990\ : LocalMux
    port map (
            O => \N__35589\,
            I => \N__35586\
        );

    \I__6989\ : Span4Mux_s0_v
    port map (
            O => \N__35586\,
            I => \N__35583\
        );

    \I__6988\ : Span4Mux_v
    port map (
            O => \N__35583\,
            I => \N__35579\
        );

    \I__6987\ : InMux
    port map (
            O => \N__35582\,
            I => \N__35576\
        );

    \I__6986\ : Odrv4
    port map (
            O => \N__35579\,
            I => \T45_c\
        );

    \I__6985\ : LocalMux
    port map (
            O => \N__35576\,
            I => \T45_c\
        );

    \I__6984\ : CascadeMux
    port map (
            O => \N__35571\,
            I => \N__35565\
        );

    \I__6983\ : InMux
    port map (
            O => \N__35570\,
            I => \N__35561\
        );

    \I__6982\ : InMux
    port map (
            O => \N__35569\,
            I => \N__35558\
        );

    \I__6981\ : CascadeMux
    port map (
            O => \N__35568\,
            I => \N__35554\
        );

    \I__6980\ : InMux
    port map (
            O => \N__35565\,
            I => \N__35551\
        );

    \I__6979\ : InMux
    port map (
            O => \N__35564\,
            I => \N__35548\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__35561\,
            I => \N__35545\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__35558\,
            I => \N__35542\
        );

    \I__6976\ : InMux
    port map (
            O => \N__35557\,
            I => \N__35539\
        );

    \I__6975\ : InMux
    port map (
            O => \N__35554\,
            I => \N__35536\
        );

    \I__6974\ : LocalMux
    port map (
            O => \N__35551\,
            I => \N__35533\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__35548\,
            I => \N__35530\
        );

    \I__6972\ : Span4Mux_h
    port map (
            O => \N__35545\,
            I => \N__35527\
        );

    \I__6971\ : Span4Mux_h
    port map (
            O => \N__35542\,
            I => \N__35524\
        );

    \I__6970\ : LocalMux
    port map (
            O => \N__35539\,
            I => \N__35521\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__35536\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__6968\ : Odrv4
    port map (
            O => \N__35533\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__6967\ : Odrv4
    port map (
            O => \N__35530\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__6966\ : Odrv4
    port map (
            O => \N__35527\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__6965\ : Odrv4
    port map (
            O => \N__35524\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__6964\ : Odrv4
    port map (
            O => \N__35521\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__6963\ : IoInMux
    port map (
            O => \N__35508\,
            I => \N__35505\
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__35505\,
            I => \N__35502\
        );

    \I__6961\ : Odrv12
    port map (
            O => \N__35502\,
            I => s2_phy_c
        );

    \I__6960\ : InMux
    port map (
            O => \N__35499\,
            I => \bfn_14_5_0_\
        );

    \I__6959\ : CascadeMux
    port map (
            O => \N__35496\,
            I => \N__35493\
        );

    \I__6958\ : InMux
    port map (
            O => \N__35493\,
            I => \N__35490\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__35490\,
            I => \phase_controller_inst2.stoper_tr.un4_running_df22\
        );

    \I__6956\ : InMux
    port map (
            O => \N__35487\,
            I => \N__35483\
        );

    \I__6955\ : InMux
    port map (
            O => \N__35486\,
            I => \N__35480\
        );

    \I__6954\ : LocalMux
    port map (
            O => \N__35483\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__35480\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__6952\ : InMux
    port map (
            O => \N__35475\,
            I => \N__35471\
        );

    \I__6951\ : InMux
    port map (
            O => \N__35474\,
            I => \N__35468\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__35471\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__35468\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__6948\ : InMux
    port map (
            O => \N__35463\,
            I => \N__35460\
        );

    \I__6947\ : LocalMux
    port map (
            O => \N__35460\,
            I => \N__35457\
        );

    \I__6946\ : Span4Mux_v
    port map (
            O => \N__35457\,
            I => \N__35454\
        );

    \I__6945\ : Odrv4
    port map (
            O => \N__35454\,
            I => \phase_controller_inst2.stoper_hc.un4_running_df20\
        );

    \I__6944\ : InMux
    port map (
            O => \N__35451\,
            I => \N__35446\
        );

    \I__6943\ : InMux
    port map (
            O => \N__35450\,
            I => \N__35443\
        );

    \I__6942\ : InMux
    port map (
            O => \N__35449\,
            I => \N__35440\
        );

    \I__6941\ : LocalMux
    port map (
            O => \N__35446\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__35443\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__35440\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__6938\ : InMux
    port map (
            O => \N__35433\,
            I => \N__35430\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__35430\,
            I => \N__35427\
        );

    \I__6936\ : Odrv12
    port map (
            O => \N__35427\,
            I => \phase_controller_inst1.start_timer_tr_0_sqmuxa\
        );

    \I__6935\ : InMux
    port map (
            O => \N__35424\,
            I => \N__35420\
        );

    \I__6934\ : InMux
    port map (
            O => \N__35423\,
            I => \N__35417\
        );

    \I__6933\ : LocalMux
    port map (
            O => \N__35420\,
            I => \phase_controller_inst1.time_passed_RNI7NN7\
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__35417\,
            I => \phase_controller_inst1.time_passed_RNI7NN7\
        );

    \I__6931\ : CascadeMux
    port map (
            O => \N__35412\,
            I => \N__35409\
        );

    \I__6930\ : InMux
    port map (
            O => \N__35409\,
            I => \N__35404\
        );

    \I__6929\ : InMux
    port map (
            O => \N__35408\,
            I => \N__35401\
        );

    \I__6928\ : InMux
    port map (
            O => \N__35407\,
            I => \N__35397\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__35404\,
            I => \N__35393\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__35401\,
            I => \N__35390\
        );

    \I__6925\ : InMux
    port map (
            O => \N__35400\,
            I => \N__35387\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__35397\,
            I => \N__35384\
        );

    \I__6923\ : InMux
    port map (
            O => \N__35396\,
            I => \N__35380\
        );

    \I__6922\ : Span4Mux_h
    port map (
            O => \N__35393\,
            I => \N__35377\
        );

    \I__6921\ : Span4Mux_h
    port map (
            O => \N__35390\,
            I => \N__35374\
        );

    \I__6920\ : LocalMux
    port map (
            O => \N__35387\,
            I => \N__35369\
        );

    \I__6919\ : Span12Mux_v
    port map (
            O => \N__35384\,
            I => \N__35369\
        );

    \I__6918\ : InMux
    port map (
            O => \N__35383\,
            I => \N__35366\
        );

    \I__6917\ : LocalMux
    port map (
            O => \N__35380\,
            I => phase_controller_inst1_state_4
        );

    \I__6916\ : Odrv4
    port map (
            O => \N__35377\,
            I => phase_controller_inst1_state_4
        );

    \I__6915\ : Odrv4
    port map (
            O => \N__35374\,
            I => phase_controller_inst1_state_4
        );

    \I__6914\ : Odrv12
    port map (
            O => \N__35369\,
            I => phase_controller_inst1_state_4
        );

    \I__6913\ : LocalMux
    port map (
            O => \N__35366\,
            I => phase_controller_inst1_state_4
        );

    \I__6912\ : InMux
    port map (
            O => \N__35355\,
            I => \N__35347\
        );

    \I__6911\ : InMux
    port map (
            O => \N__35354\,
            I => \N__35347\
        );

    \I__6910\ : InMux
    port map (
            O => \N__35353\,
            I => \N__35342\
        );

    \I__6909\ : InMux
    port map (
            O => \N__35352\,
            I => \N__35342\
        );

    \I__6908\ : LocalMux
    port map (
            O => \N__35347\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6907\ : LocalMux
    port map (
            O => \N__35342\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6906\ : InMux
    port map (
            O => \N__35337\,
            I => \N__35334\
        );

    \I__6905\ : LocalMux
    port map (
            O => \N__35334\,
            I => \N__35331\
        );

    \I__6904\ : Odrv12
    port map (
            O => \N__35331\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO\
        );

    \I__6903\ : InMux
    port map (
            O => \N__35328\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_28\
        );

    \I__6902\ : InMux
    port map (
            O => \N__35325\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30\
        );

    \I__6901\ : InMux
    port map (
            O => \N__35322\,
            I => \N__35316\
        );

    \I__6900\ : InMux
    port map (
            O => \N__35321\,
            I => \N__35316\
        );

    \I__6899\ : LocalMux
    port map (
            O => \N__35316\,
            I => \N__35313\
        );

    \I__6898\ : Odrv12
    port map (
            O => \N__35313\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__6897\ : InMux
    port map (
            O => \N__35310\,
            I => \N__35306\
        );

    \I__6896\ : InMux
    port map (
            O => \N__35309\,
            I => \N__35303\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__35306\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__6894\ : LocalMux
    port map (
            O => \N__35303\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__6893\ : InMux
    port map (
            O => \N__35298\,
            I => \N__35294\
        );

    \I__6892\ : InMux
    port map (
            O => \N__35297\,
            I => \N__35291\
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__35294\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__6890\ : LocalMux
    port map (
            O => \N__35291\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__6889\ : InMux
    port map (
            O => \N__35286\,
            I => \N__35283\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__35283\,
            I => \N__35280\
        );

    \I__6887\ : Odrv4
    port map (
            O => \N__35280\,
            I => \phase_controller_inst2.stoper_hc.un4_running_df22\
        );

    \I__6886\ : InMux
    port map (
            O => \N__35277\,
            I => \N__35273\
        );

    \I__6885\ : InMux
    port map (
            O => \N__35276\,
            I => \N__35270\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__35273\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__35270\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__6882\ : InMux
    port map (
            O => \N__35265\,
            I => \N__35261\
        );

    \I__6881\ : InMux
    port map (
            O => \N__35264\,
            I => \N__35258\
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__35261\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__35258\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__6878\ : CascadeMux
    port map (
            O => \N__35253\,
            I => \N__35250\
        );

    \I__6877\ : InMux
    port map (
            O => \N__35250\,
            I => \N__35247\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__35247\,
            I => \N__35244\
        );

    \I__6875\ : Odrv4
    port map (
            O => \N__35244\,
            I => \phase_controller_inst2.stoper_hc.un4_running_df24\
        );

    \I__6874\ : InMux
    port map (
            O => \N__35241\,
            I => \N__35237\
        );

    \I__6873\ : InMux
    port map (
            O => \N__35240\,
            I => \N__35234\
        );

    \I__6872\ : LocalMux
    port map (
            O => \N__35237\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__35234\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__6870\ : InMux
    port map (
            O => \N__35229\,
            I => \N__35225\
        );

    \I__6869\ : InMux
    port map (
            O => \N__35228\,
            I => \N__35222\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__35225\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__35222\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__6866\ : CascadeMux
    port map (
            O => \N__35217\,
            I => \N__35214\
        );

    \I__6865\ : InMux
    port map (
            O => \N__35214\,
            I => \N__35211\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__35211\,
            I => \N__35208\
        );

    \I__6863\ : Odrv4
    port map (
            O => \N__35208\,
            I => \phase_controller_inst2.stoper_hc.un4_running_df26\
        );

    \I__6862\ : InMux
    port map (
            O => \N__35205\,
            I => \N__35201\
        );

    \I__6861\ : InMux
    port map (
            O => \N__35204\,
            I => \N__35198\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__35201\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__35198\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__6858\ : InMux
    port map (
            O => \N__35193\,
            I => \N__35189\
        );

    \I__6857\ : InMux
    port map (
            O => \N__35192\,
            I => \N__35186\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__35189\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__35186\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__6854\ : InMux
    port map (
            O => \N__35181\,
            I => \N__35178\
        );

    \I__6853\ : LocalMux
    port map (
            O => \N__35178\,
            I => \N__35175\
        );

    \I__6852\ : Odrv4
    port map (
            O => \N__35175\,
            I => \phase_controller_inst2.stoper_hc.un4_running_df28\
        );

    \I__6851\ : InMux
    port map (
            O => \N__35172\,
            I => \N__35168\
        );

    \I__6850\ : InMux
    port map (
            O => \N__35171\,
            I => \N__35165\
        );

    \I__6849\ : LocalMux
    port map (
            O => \N__35168\,
            I => \N__35158\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__35165\,
            I => \N__35158\
        );

    \I__6847\ : InMux
    port map (
            O => \N__35164\,
            I => \N__35155\
        );

    \I__6846\ : InMux
    port map (
            O => \N__35163\,
            I => \N__35152\
        );

    \I__6845\ : Span4Mux_v
    port map (
            O => \N__35158\,
            I => \N__35149\
        );

    \I__6844\ : LocalMux
    port map (
            O => \N__35155\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__35152\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__6842\ : Odrv4
    port map (
            O => \N__35149\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__6841\ : InMux
    port map (
            O => \N__35142\,
            I => \N__35139\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__35139\,
            I => \N__35134\
        );

    \I__6839\ : InMux
    port map (
            O => \N__35138\,
            I => \N__35131\
        );

    \I__6838\ : InMux
    port map (
            O => \N__35137\,
            I => \N__35128\
        );

    \I__6837\ : Span4Mux_h
    port map (
            O => \N__35134\,
            I => \N__35125\
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__35131\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__35128\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__6834\ : Odrv4
    port map (
            O => \N__35125\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__6833\ : CascadeMux
    port map (
            O => \N__35118\,
            I => \N__35115\
        );

    \I__6832\ : InMux
    port map (
            O => \N__35115\,
            I => \N__35112\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__35112\,
            I => \N__35109\
        );

    \I__6830\ : Odrv4
    port map (
            O => \N__35109\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\
        );

    \I__6829\ : InMux
    port map (
            O => \N__35106\,
            I => \N__35103\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__35103\,
            I => \phase_controller_inst2.stoper_tr.un4_running_df20\
        );

    \I__6827\ : CascadeMux
    port map (
            O => \N__35100\,
            I => \N__35097\
        );

    \I__6826\ : InMux
    port map (
            O => \N__35097\,
            I => \N__35094\
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__35094\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\
        );

    \I__6824\ : InMux
    port map (
            O => \N__35091\,
            I => \N__35088\
        );

    \I__6823\ : LocalMux
    port map (
            O => \N__35088\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\
        );

    \I__6822\ : InMux
    port map (
            O => \N__35085\,
            I => \N__35082\
        );

    \I__6821\ : LocalMux
    port map (
            O => \N__35082\,
            I => \N__35079\
        );

    \I__6820\ : Span4Mux_v
    port map (
            O => \N__35079\,
            I => \N__35076\
        );

    \I__6819\ : Odrv4
    port map (
            O => \N__35076\,
            I => \phase_controller_inst2.stoper_tr.un4_running_df26\
        );

    \I__6818\ : InMux
    port map (
            O => \N__35073\,
            I => \N__35070\
        );

    \I__6817\ : LocalMux
    port map (
            O => \N__35070\,
            I => \N__35067\
        );

    \I__6816\ : Span4Mux_v
    port map (
            O => \N__35067\,
            I => \N__35064\
        );

    \I__6815\ : Odrv4
    port map (
            O => \N__35064\,
            I => \phase_controller_inst2.stoper_tr.un4_running_df28\
        );

    \I__6814\ : InMux
    port map (
            O => \N__35061\,
            I => \N__35058\
        );

    \I__6813\ : LocalMux
    port map (
            O => \N__35058\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\
        );

    \I__6812\ : CascadeMux
    port map (
            O => \N__35055\,
            I => \N__35052\
        );

    \I__6811\ : InMux
    port map (
            O => \N__35052\,
            I => \N__35049\
        );

    \I__6810\ : LocalMux
    port map (
            O => \N__35049\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\
        );

    \I__6809\ : CascadeMux
    port map (
            O => \N__35046\,
            I => \N__35043\
        );

    \I__6808\ : InMux
    port map (
            O => \N__35043\,
            I => \N__35040\
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__35040\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\
        );

    \I__6806\ : CascadeMux
    port map (
            O => \N__35037\,
            I => \N__35034\
        );

    \I__6805\ : InMux
    port map (
            O => \N__35034\,
            I => \N__35031\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__35031\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\
        );

    \I__6803\ : CascadeMux
    port map (
            O => \N__35028\,
            I => \N__35025\
        );

    \I__6802\ : InMux
    port map (
            O => \N__35025\,
            I => \N__35022\
        );

    \I__6801\ : LocalMux
    port map (
            O => \N__35022\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\
        );

    \I__6800\ : CascadeMux
    port map (
            O => \N__35019\,
            I => \N__35016\
        );

    \I__6799\ : InMux
    port map (
            O => \N__35016\,
            I => \N__35013\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__35013\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\
        );

    \I__6797\ : CascadeMux
    port map (
            O => \N__35010\,
            I => \N__35007\
        );

    \I__6796\ : InMux
    port map (
            O => \N__35007\,
            I => \N__35004\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__35004\,
            I => \N__35001\
        );

    \I__6794\ : Odrv4
    port map (
            O => \N__35001\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\
        );

    \I__6793\ : CascadeMux
    port map (
            O => \N__34998\,
            I => \N__34995\
        );

    \I__6792\ : InMux
    port map (
            O => \N__34995\,
            I => \N__34992\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__34992\,
            I => \N__34989\
        );

    \I__6790\ : Odrv4
    port map (
            O => \N__34989\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\
        );

    \I__6789\ : InMux
    port map (
            O => \N__34986\,
            I => \N__34981\
        );

    \I__6788\ : InMux
    port map (
            O => \N__34985\,
            I => \N__34978\
        );

    \I__6787\ : InMux
    port map (
            O => \N__34984\,
            I => \N__34975\
        );

    \I__6786\ : LocalMux
    port map (
            O => \N__34981\,
            I => \N__34970\
        );

    \I__6785\ : LocalMux
    port map (
            O => \N__34978\,
            I => \N__34970\
        );

    \I__6784\ : LocalMux
    port map (
            O => \N__34975\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__6783\ : Odrv12
    port map (
            O => \N__34970\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__6782\ : InMux
    port map (
            O => \N__34965\,
            I => \N__34959\
        );

    \I__6781\ : InMux
    port map (
            O => \N__34964\,
            I => \N__34959\
        );

    \I__6780\ : LocalMux
    port map (
            O => \N__34959\,
            I => \N__34954\
        );

    \I__6779\ : CascadeMux
    port map (
            O => \N__34958\,
            I => \N__34951\
        );

    \I__6778\ : InMux
    port map (
            O => \N__34957\,
            I => \N__34948\
        );

    \I__6777\ : Span4Mux_h
    port map (
            O => \N__34954\,
            I => \N__34945\
        );

    \I__6776\ : InMux
    port map (
            O => \N__34951\,
            I => \N__34942\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__34948\,
            I => \N__34939\
        );

    \I__6774\ : Span4Mux_h
    port map (
            O => \N__34945\,
            I => \N__34936\
        );

    \I__6773\ : LocalMux
    port map (
            O => \N__34942\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__6772\ : Odrv4
    port map (
            O => \N__34939\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__6771\ : Odrv4
    port map (
            O => \N__34936\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__6770\ : InMux
    port map (
            O => \N__34929\,
            I => \N__34926\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__34926\,
            I => \N__34923\
        );

    \I__6768\ : Span4Mux_h
    port map (
            O => \N__34923\,
            I => \N__34920\
        );

    \I__6767\ : Span4Mux_h
    port map (
            O => \N__34920\,
            I => \N__34913\
        );

    \I__6766\ : InMux
    port map (
            O => \N__34919\,
            I => \N__34904\
        );

    \I__6765\ : InMux
    port map (
            O => \N__34918\,
            I => \N__34904\
        );

    \I__6764\ : InMux
    port map (
            O => \N__34917\,
            I => \N__34904\
        );

    \I__6763\ : InMux
    port map (
            O => \N__34916\,
            I => \N__34904\
        );

    \I__6762\ : Odrv4
    port map (
            O => \N__34913\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__34904\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__6760\ : CascadeMux
    port map (
            O => \N__34899\,
            I => \N__34895\
        );

    \I__6759\ : CascadeMux
    port map (
            O => \N__34898\,
            I => \N__34892\
        );

    \I__6758\ : InMux
    port map (
            O => \N__34895\,
            I => \N__34884\
        );

    \I__6757\ : InMux
    port map (
            O => \N__34892\,
            I => \N__34884\
        );

    \I__6756\ : InMux
    port map (
            O => \N__34891\,
            I => \N__34881\
        );

    \I__6755\ : InMux
    port map (
            O => \N__34890\,
            I => \N__34876\
        );

    \I__6754\ : InMux
    port map (
            O => \N__34889\,
            I => \N__34876\
        );

    \I__6753\ : LocalMux
    port map (
            O => \N__34884\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__34881\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__34876\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__6750\ : InMux
    port map (
            O => \N__34869\,
            I => \N__34865\
        );

    \I__6749\ : InMux
    port map (
            O => \N__34868\,
            I => \N__34862\
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__34865\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__6747\ : LocalMux
    port map (
            O => \N__34862\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__6746\ : CascadeMux
    port map (
            O => \N__34857\,
            I => \N__34854\
        );

    \I__6745\ : InMux
    port map (
            O => \N__34854\,
            I => \N__34851\
        );

    \I__6744\ : LocalMux
    port map (
            O => \N__34851\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\
        );

    \I__6743\ : CascadeMux
    port map (
            O => \N__34848\,
            I => \N__34845\
        );

    \I__6742\ : InMux
    port map (
            O => \N__34845\,
            I => \N__34842\
        );

    \I__6741\ : LocalMux
    port map (
            O => \N__34842\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\
        );

    \I__6740\ : CascadeMux
    port map (
            O => \N__34839\,
            I => \N__34836\
        );

    \I__6739\ : InMux
    port map (
            O => \N__34836\,
            I => \N__34833\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__34833\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\
        );

    \I__6737\ : CascadeMux
    port map (
            O => \N__34830\,
            I => \N__34827\
        );

    \I__6736\ : InMux
    port map (
            O => \N__34827\,
            I => \N__34824\
        );

    \I__6735\ : LocalMux
    port map (
            O => \N__34824\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\
        );

    \I__6734\ : CascadeMux
    port map (
            O => \N__34821\,
            I => \N__34818\
        );

    \I__6733\ : InMux
    port map (
            O => \N__34818\,
            I => \N__34815\
        );

    \I__6732\ : LocalMux
    port map (
            O => \N__34815\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\
        );

    \I__6731\ : InMux
    port map (
            O => \N__34812\,
            I => \N__34809\
        );

    \I__6730\ : LocalMux
    port map (
            O => \N__34809\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\
        );

    \I__6729\ : InMux
    port map (
            O => \N__34806\,
            I => \current_shift_inst.control_input_cry_10\
        );

    \I__6728\ : InMux
    port map (
            O => \N__34803\,
            I => \N__34800\
        );

    \I__6727\ : LocalMux
    port map (
            O => \N__34800\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\
        );

    \I__6726\ : InMux
    port map (
            O => \N__34797\,
            I => \current_shift_inst.control_input_cry_11\
        );

    \I__6725\ : InMux
    port map (
            O => \N__34794\,
            I => \current_shift_inst.control_input_cry_12\
        );

    \I__6724\ : InMux
    port map (
            O => \N__34791\,
            I => \N__34787\
        );

    \I__6723\ : InMux
    port map (
            O => \N__34790\,
            I => \N__34784\
        );

    \I__6722\ : LocalMux
    port map (
            O => \N__34787\,
            I => \current_shift_inst.control_input_31\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__34784\,
            I => \current_shift_inst.control_input_31\
        );

    \I__6720\ : CascadeMux
    port map (
            O => \N__34779\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\
        );

    \I__6719\ : InMux
    port map (
            O => \N__34776\,
            I => \N__34770\
        );

    \I__6718\ : InMux
    port map (
            O => \N__34775\,
            I => \N__34770\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__34770\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__6716\ : InMux
    port map (
            O => \N__34767\,
            I => \N__34764\
        );

    \I__6715\ : LocalMux
    port map (
            O => \N__34764\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\
        );

    \I__6714\ : InMux
    port map (
            O => \N__34761\,
            I => \current_shift_inst.control_input_cry_2\
        );

    \I__6713\ : InMux
    port map (
            O => \N__34758\,
            I => \N__34755\
        );

    \I__6712\ : LocalMux
    port map (
            O => \N__34755\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\
        );

    \I__6711\ : InMux
    port map (
            O => \N__34752\,
            I => \current_shift_inst.control_input_cry_3\
        );

    \I__6710\ : InMux
    port map (
            O => \N__34749\,
            I => \N__34746\
        );

    \I__6709\ : LocalMux
    port map (
            O => \N__34746\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\
        );

    \I__6708\ : InMux
    port map (
            O => \N__34743\,
            I => \current_shift_inst.control_input_cry_4\
        );

    \I__6707\ : InMux
    port map (
            O => \N__34740\,
            I => \N__34737\
        );

    \I__6706\ : LocalMux
    port map (
            O => \N__34737\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\
        );

    \I__6705\ : InMux
    port map (
            O => \N__34734\,
            I => \current_shift_inst.control_input_cry_5\
        );

    \I__6704\ : InMux
    port map (
            O => \N__34731\,
            I => \N__34728\
        );

    \I__6703\ : LocalMux
    port map (
            O => \N__34728\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\
        );

    \I__6702\ : InMux
    port map (
            O => \N__34725\,
            I => \current_shift_inst.control_input_cry_6\
        );

    \I__6701\ : InMux
    port map (
            O => \N__34722\,
            I => \N__34719\
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__34719\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\
        );

    \I__6699\ : InMux
    port map (
            O => \N__34716\,
            I => \bfn_13_12_0_\
        );

    \I__6698\ : InMux
    port map (
            O => \N__34713\,
            I => \N__34710\
        );

    \I__6697\ : LocalMux
    port map (
            O => \N__34710\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\
        );

    \I__6696\ : InMux
    port map (
            O => \N__34707\,
            I => \current_shift_inst.control_input_cry_8\
        );

    \I__6695\ : InMux
    port map (
            O => \N__34704\,
            I => \N__34701\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__34701\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\
        );

    \I__6693\ : InMux
    port map (
            O => \N__34698\,
            I => \current_shift_inst.control_input_cry_9\
        );

    \I__6692\ : InMux
    port map (
            O => \N__34695\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__6691\ : InMux
    port map (
            O => \N__34692\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__6690\ : InMux
    port map (
            O => \N__34689\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__6689\ : InMux
    port map (
            O => \N__34686\,
            I => \N__34683\
        );

    \I__6688\ : LocalMux
    port map (
            O => \N__34683\,
            I => \current_shift_inst.control_input_18\
        );

    \I__6687\ : InMux
    port map (
            O => \N__34680\,
            I => \N__34677\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__34677\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\
        );

    \I__6685\ : InMux
    port map (
            O => \N__34674\,
            I => \current_shift_inst.control_input_cry_0\
        );

    \I__6684\ : InMux
    port map (
            O => \N__34671\,
            I => \N__34668\
        );

    \I__6683\ : LocalMux
    port map (
            O => \N__34668\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\
        );

    \I__6682\ : InMux
    port map (
            O => \N__34665\,
            I => \current_shift_inst.control_input_cry_1\
        );

    \I__6681\ : InMux
    port map (
            O => \N__34662\,
            I => \bfn_13_9_0_\
        );

    \I__6680\ : InMux
    port map (
            O => \N__34659\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__6679\ : InMux
    port map (
            O => \N__34656\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__6678\ : InMux
    port map (
            O => \N__34653\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__6677\ : InMux
    port map (
            O => \N__34650\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__6676\ : InMux
    port map (
            O => \N__34647\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__6675\ : InMux
    port map (
            O => \N__34644\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__6674\ : InMux
    port map (
            O => \N__34641\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__6673\ : InMux
    port map (
            O => \N__34638\,
            I => \bfn_13_10_0_\
        );

    \I__6672\ : InMux
    port map (
            O => \N__34635\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__6671\ : InMux
    port map (
            O => \N__34632\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__6670\ : InMux
    port map (
            O => \N__34629\,
            I => \bfn_13_8_0_\
        );

    \I__6669\ : InMux
    port map (
            O => \N__34626\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__6668\ : InMux
    port map (
            O => \N__34623\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__6667\ : InMux
    port map (
            O => \N__34620\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__6666\ : InMux
    port map (
            O => \N__34617\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__6665\ : InMux
    port map (
            O => \N__34614\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__6664\ : InMux
    port map (
            O => \N__34611\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__6663\ : InMux
    port map (
            O => \N__34608\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__6662\ : InMux
    port map (
            O => \N__34605\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__6661\ : InMux
    port map (
            O => \N__34602\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__6660\ : InMux
    port map (
            O => \N__34599\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__6659\ : InMux
    port map (
            O => \N__34596\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__6658\ : InMux
    port map (
            O => \N__34593\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__6657\ : InMux
    port map (
            O => \N__34590\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__6656\ : InMux
    port map (
            O => \N__34587\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\
        );

    \I__6655\ : InMux
    port map (
            O => \N__34584\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\
        );

    \I__6654\ : InMux
    port map (
            O => \N__34581\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\
        );

    \I__6653\ : InMux
    port map (
            O => \N__34578\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\
        );

    \I__6652\ : CEMux
    port map (
            O => \N__34575\,
            I => \N__34564\
        );

    \I__6651\ : CEMux
    port map (
            O => \N__34574\,
            I => \N__34548\
        );

    \I__6650\ : InMux
    port map (
            O => \N__34573\,
            I => \N__34541\
        );

    \I__6649\ : InMux
    port map (
            O => \N__34572\,
            I => \N__34541\
        );

    \I__6648\ : InMux
    port map (
            O => \N__34571\,
            I => \N__34541\
        );

    \I__6647\ : InMux
    port map (
            O => \N__34570\,
            I => \N__34532\
        );

    \I__6646\ : InMux
    port map (
            O => \N__34569\,
            I => \N__34532\
        );

    \I__6645\ : InMux
    port map (
            O => \N__34568\,
            I => \N__34532\
        );

    \I__6644\ : InMux
    port map (
            O => \N__34567\,
            I => \N__34532\
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__34564\,
            I => \N__34525\
        );

    \I__6642\ : InMux
    port map (
            O => \N__34563\,
            I => \N__34516\
        );

    \I__6641\ : InMux
    port map (
            O => \N__34562\,
            I => \N__34516\
        );

    \I__6640\ : InMux
    port map (
            O => \N__34561\,
            I => \N__34516\
        );

    \I__6639\ : InMux
    port map (
            O => \N__34560\,
            I => \N__34516\
        );

    \I__6638\ : CEMux
    port map (
            O => \N__34559\,
            I => \N__34503\
        );

    \I__6637\ : CEMux
    port map (
            O => \N__34558\,
            I => \N__34499\
        );

    \I__6636\ : InMux
    port map (
            O => \N__34557\,
            I => \N__34492\
        );

    \I__6635\ : InMux
    port map (
            O => \N__34556\,
            I => \N__34492\
        );

    \I__6634\ : InMux
    port map (
            O => \N__34555\,
            I => \N__34492\
        );

    \I__6633\ : InMux
    port map (
            O => \N__34554\,
            I => \N__34483\
        );

    \I__6632\ : InMux
    port map (
            O => \N__34553\,
            I => \N__34483\
        );

    \I__6631\ : InMux
    port map (
            O => \N__34552\,
            I => \N__34483\
        );

    \I__6630\ : InMux
    port map (
            O => \N__34551\,
            I => \N__34483\
        );

    \I__6629\ : LocalMux
    port map (
            O => \N__34548\,
            I => \N__34480\
        );

    \I__6628\ : LocalMux
    port map (
            O => \N__34541\,
            I => \N__34477\
        );

    \I__6627\ : LocalMux
    port map (
            O => \N__34532\,
            I => \N__34474\
        );

    \I__6626\ : InMux
    port map (
            O => \N__34531\,
            I => \N__34465\
        );

    \I__6625\ : InMux
    port map (
            O => \N__34530\,
            I => \N__34465\
        );

    \I__6624\ : InMux
    port map (
            O => \N__34529\,
            I => \N__34465\
        );

    \I__6623\ : InMux
    port map (
            O => \N__34528\,
            I => \N__34465\
        );

    \I__6622\ : Span4Mux_h
    port map (
            O => \N__34525\,
            I => \N__34460\
        );

    \I__6621\ : LocalMux
    port map (
            O => \N__34516\,
            I => \N__34460\
        );

    \I__6620\ : InMux
    port map (
            O => \N__34515\,
            I => \N__34451\
        );

    \I__6619\ : InMux
    port map (
            O => \N__34514\,
            I => \N__34451\
        );

    \I__6618\ : InMux
    port map (
            O => \N__34513\,
            I => \N__34451\
        );

    \I__6617\ : InMux
    port map (
            O => \N__34512\,
            I => \N__34451\
        );

    \I__6616\ : InMux
    port map (
            O => \N__34511\,
            I => \N__34442\
        );

    \I__6615\ : InMux
    port map (
            O => \N__34510\,
            I => \N__34442\
        );

    \I__6614\ : InMux
    port map (
            O => \N__34509\,
            I => \N__34442\
        );

    \I__6613\ : InMux
    port map (
            O => \N__34508\,
            I => \N__34442\
        );

    \I__6612\ : CEMux
    port map (
            O => \N__34507\,
            I => \N__34438\
        );

    \I__6611\ : CEMux
    port map (
            O => \N__34506\,
            I => \N__34435\
        );

    \I__6610\ : LocalMux
    port map (
            O => \N__34503\,
            I => \N__34432\
        );

    \I__6609\ : CEMux
    port map (
            O => \N__34502\,
            I => \N__34429\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__34499\,
            I => \N__34426\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__34492\,
            I => \N__34407\
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__34483\,
            I => \N__34407\
        );

    \I__6605\ : Span4Mux_v
    port map (
            O => \N__34480\,
            I => \N__34407\
        );

    \I__6604\ : Span4Mux_v
    port map (
            O => \N__34477\,
            I => \N__34407\
        );

    \I__6603\ : Span4Mux_h
    port map (
            O => \N__34474\,
            I => \N__34407\
        );

    \I__6602\ : LocalMux
    port map (
            O => \N__34465\,
            I => \N__34407\
        );

    \I__6601\ : Span4Mux_v
    port map (
            O => \N__34460\,
            I => \N__34407\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__34451\,
            I => \N__34407\
        );

    \I__6599\ : LocalMux
    port map (
            O => \N__34442\,
            I => \N__34407\
        );

    \I__6598\ : InMux
    port map (
            O => \N__34441\,
            I => \N__34404\
        );

    \I__6597\ : LocalMux
    port map (
            O => \N__34438\,
            I => \N__34401\
        );

    \I__6596\ : LocalMux
    port map (
            O => \N__34435\,
            I => \N__34396\
        );

    \I__6595\ : Span4Mux_h
    port map (
            O => \N__34432\,
            I => \N__34396\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__34429\,
            I => \N__34391\
        );

    \I__6593\ : Span4Mux_h
    port map (
            O => \N__34426\,
            I => \N__34391\
        );

    \I__6592\ : Span4Mux_v
    port map (
            O => \N__34407\,
            I => \N__34386\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__34404\,
            I => \N__34386\
        );

    \I__6590\ : Span4Mux_h
    port map (
            O => \N__34401\,
            I => \N__34383\
        );

    \I__6589\ : Span4Mux_h
    port map (
            O => \N__34396\,
            I => \N__34378\
        );

    \I__6588\ : Span4Mux_h
    port map (
            O => \N__34391\,
            I => \N__34378\
        );

    \I__6587\ : Span4Mux_h
    port map (
            O => \N__34386\,
            I => \N__34375\
        );

    \I__6586\ : Odrv4
    port map (
            O => \N__34383\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__6585\ : Odrv4
    port map (
            O => \N__34378\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__6584\ : Odrv4
    port map (
            O => \N__34375\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__6583\ : InMux
    port map (
            O => \N__34368\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\
        );

    \I__6582\ : InMux
    port map (
            O => \N__34365\,
            I => \N__34362\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__34362\,
            I => \N__34358\
        );

    \I__6580\ : InMux
    port map (
            O => \N__34361\,
            I => \N__34354\
        );

    \I__6579\ : Span4Mux_h
    port map (
            O => \N__34358\,
            I => \N__34351\
        );

    \I__6578\ : InMux
    port map (
            O => \N__34357\,
            I => \N__34348\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__34354\,
            I => \N__34341\
        );

    \I__6576\ : Sp12to4
    port map (
            O => \N__34351\,
            I => \N__34341\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__34348\,
            I => \N__34341\
        );

    \I__6574\ : Span12Mux_s10_v
    port map (
            O => \N__34341\,
            I => \N__34338\
        );

    \I__6573\ : Odrv12
    port map (
            O => \N__34338\,
            I => \il_min_comp1_D2\
        );

    \I__6572\ : IoInMux
    port map (
            O => \N__34335\,
            I => \N__34332\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__34332\,
            I => \N__34329\
        );

    \I__6570\ : IoSpan4Mux
    port map (
            O => \N__34329\,
            I => \N__34326\
        );

    \I__6569\ : Span4Mux_s0_v
    port map (
            O => \N__34326\,
            I => \N__34323\
        );

    \I__6568\ : Span4Mux_v
    port map (
            O => \N__34323\,
            I => \N__34319\
        );

    \I__6567\ : InMux
    port map (
            O => \N__34322\,
            I => \N__34316\
        );

    \I__6566\ : Odrv4
    port map (
            O => \N__34319\,
            I => \T12_c\
        );

    \I__6565\ : LocalMux
    port map (
            O => \N__34316\,
            I => \T12_c\
        );

    \I__6564\ : InMux
    port map (
            O => \N__34311\,
            I => \N__34303\
        );

    \I__6563\ : InMux
    port map (
            O => \N__34310\,
            I => \N__34303\
        );

    \I__6562\ : InMux
    port map (
            O => \N__34309\,
            I => \N__34299\
        );

    \I__6561\ : InMux
    port map (
            O => \N__34308\,
            I => \N__34296\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__34303\,
            I => \N__34293\
        );

    \I__6559\ : InMux
    port map (
            O => \N__34302\,
            I => \N__34290\
        );

    \I__6558\ : LocalMux
    port map (
            O => \N__34299\,
            I => \N__34287\
        );

    \I__6557\ : LocalMux
    port map (
            O => \N__34296\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__6556\ : Odrv4
    port map (
            O => \N__34293\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__6555\ : LocalMux
    port map (
            O => \N__34290\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__6554\ : Odrv4
    port map (
            O => \N__34287\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__6553\ : IoInMux
    port map (
            O => \N__34278\,
            I => \N__34275\
        );

    \I__6552\ : LocalMux
    port map (
            O => \N__34275\,
            I => \N__34272\
        );

    \I__6551\ : Span4Mux_s0_v
    port map (
            O => \N__34272\,
            I => \N__34269\
        );

    \I__6550\ : Span4Mux_v
    port map (
            O => \N__34269\,
            I => \N__34266\
        );

    \I__6549\ : Sp12to4
    port map (
            O => \N__34266\,
            I => \N__34262\
        );

    \I__6548\ : InMux
    port map (
            O => \N__34265\,
            I => \N__34259\
        );

    \I__6547\ : Odrv12
    port map (
            O => \N__34262\,
            I => \T01_c\
        );

    \I__6546\ : LocalMux
    port map (
            O => \N__34259\,
            I => \T01_c\
        );

    \I__6545\ : CascadeMux
    port map (
            O => \N__34254\,
            I => \N__34250\
        );

    \I__6544\ : InMux
    port map (
            O => \N__34253\,
            I => \N__34247\
        );

    \I__6543\ : InMux
    port map (
            O => \N__34250\,
            I => \N__34243\
        );

    \I__6542\ : LocalMux
    port map (
            O => \N__34247\,
            I => \N__34240\
        );

    \I__6541\ : InMux
    port map (
            O => \N__34246\,
            I => \N__34237\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__34243\,
            I => \N__34232\
        );

    \I__6539\ : Span4Mux_h
    port map (
            O => \N__34240\,
            I => \N__34232\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__34237\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__6537\ : Odrv4
    port map (
            O => \N__34232\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__6536\ : InMux
    port map (
            O => \N__34227\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__6535\ : CascadeMux
    port map (
            O => \N__34224\,
            I => \N__34221\
        );

    \I__6534\ : InMux
    port map (
            O => \N__34221\,
            I => \N__34218\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__34218\,
            I => \N__34213\
        );

    \I__6532\ : InMux
    port map (
            O => \N__34217\,
            I => \N__34210\
        );

    \I__6531\ : InMux
    port map (
            O => \N__34216\,
            I => \N__34207\
        );

    \I__6530\ : Span4Mux_v
    port map (
            O => \N__34213\,
            I => \N__34204\
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__34210\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__34207\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__6527\ : Odrv4
    port map (
            O => \N__34204\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__6526\ : InMux
    port map (
            O => \N__34197\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__6525\ : InMux
    port map (
            O => \N__34194\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\
        );

    \I__6524\ : InMux
    port map (
            O => \N__34191\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__6523\ : InMux
    port map (
            O => \N__34188\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\
        );

    \I__6522\ : InMux
    port map (
            O => \N__34185\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\
        );

    \I__6521\ : InMux
    port map (
            O => \N__34182\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\
        );

    \I__6520\ : InMux
    port map (
            O => \N__34179\,
            I => \bfn_12_20_0_\
        );

    \I__6519\ : InMux
    port map (
            O => \N__34176\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\
        );

    \I__6518\ : InMux
    port map (
            O => \N__34173\,
            I => \N__34169\
        );

    \I__6517\ : InMux
    port map (
            O => \N__34172\,
            I => \N__34166\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__34169\,
            I => \N__34163\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__34166\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__6514\ : Odrv4
    port map (
            O => \N__34163\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__6513\ : InMux
    port map (
            O => \N__34158\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__6512\ : InMux
    port map (
            O => \N__34155\,
            I => \N__34151\
        );

    \I__6511\ : InMux
    port map (
            O => \N__34154\,
            I => \N__34148\
        );

    \I__6510\ : LocalMux
    port map (
            O => \N__34151\,
            I => \N__34145\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__34148\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__6508\ : Odrv4
    port map (
            O => \N__34145\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__6507\ : InMux
    port map (
            O => \N__34140\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__6506\ : InMux
    port map (
            O => \N__34137\,
            I => \N__34133\
        );

    \I__6505\ : InMux
    port map (
            O => \N__34136\,
            I => \N__34130\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__34133\,
            I => \N__34127\
        );

    \I__6503\ : LocalMux
    port map (
            O => \N__34130\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__6502\ : Odrv4
    port map (
            O => \N__34127\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__6501\ : InMux
    port map (
            O => \N__34122\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__6500\ : InMux
    port map (
            O => \N__34119\,
            I => \N__34115\
        );

    \I__6499\ : InMux
    port map (
            O => \N__34118\,
            I => \N__34112\
        );

    \I__6498\ : LocalMux
    port map (
            O => \N__34115\,
            I => \N__34109\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__34112\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__6496\ : Odrv4
    port map (
            O => \N__34109\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__6495\ : InMux
    port map (
            O => \N__34104\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__6494\ : InMux
    port map (
            O => \N__34101\,
            I => \N__34097\
        );

    \I__6493\ : InMux
    port map (
            O => \N__34100\,
            I => \N__34094\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__34097\,
            I => \N__34091\
        );

    \I__6491\ : LocalMux
    port map (
            O => \N__34094\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__6490\ : Odrv4
    port map (
            O => \N__34091\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__6489\ : InMux
    port map (
            O => \N__34086\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__6488\ : InMux
    port map (
            O => \N__34083\,
            I => \N__34079\
        );

    \I__6487\ : InMux
    port map (
            O => \N__34082\,
            I => \N__34076\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__34079\,
            I => \N__34073\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__34076\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__6484\ : Odrv12
    port map (
            O => \N__34073\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__6483\ : InMux
    port map (
            O => \N__34068\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__6482\ : CascadeMux
    port map (
            O => \N__34065\,
            I => \N__34061\
        );

    \I__6481\ : InMux
    port map (
            O => \N__34064\,
            I => \N__34056\
        );

    \I__6480\ : InMux
    port map (
            O => \N__34061\,
            I => \N__34056\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__34056\,
            I => \N__34052\
        );

    \I__6478\ : InMux
    port map (
            O => \N__34055\,
            I => \N__34049\
        );

    \I__6477\ : Span4Mux_h
    port map (
            O => \N__34052\,
            I => \N__34046\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__34049\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__6475\ : Odrv4
    port map (
            O => \N__34046\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__6474\ : InMux
    port map (
            O => \N__34041\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__6473\ : CascadeMux
    port map (
            O => \N__34038\,
            I => \N__34034\
        );

    \I__6472\ : InMux
    port map (
            O => \N__34037\,
            I => \N__34029\
        );

    \I__6471\ : InMux
    port map (
            O => \N__34034\,
            I => \N__34029\
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__34029\,
            I => \N__34025\
        );

    \I__6469\ : InMux
    port map (
            O => \N__34028\,
            I => \N__34022\
        );

    \I__6468\ : Span4Mux_h
    port map (
            O => \N__34025\,
            I => \N__34019\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__34022\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__6466\ : Odrv4
    port map (
            O => \N__34019\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__6465\ : InMux
    port map (
            O => \N__34014\,
            I => \bfn_12_19_0_\
        );

    \I__6464\ : CascadeMux
    port map (
            O => \N__34011\,
            I => \N__34008\
        );

    \I__6463\ : InMux
    port map (
            O => \N__34008\,
            I => \N__34005\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__34005\,
            I => \N__34002\
        );

    \I__6461\ : Odrv4
    port map (
            O => \N__34002\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\
        );

    \I__6460\ : InMux
    port map (
            O => \N__33999\,
            I => \N__33995\
        );

    \I__6459\ : InMux
    port map (
            O => \N__33998\,
            I => \N__33992\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__33995\,
            I => \N__33989\
        );

    \I__6457\ : LocalMux
    port map (
            O => \N__33992\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__6456\ : Odrv4
    port map (
            O => \N__33989\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__6455\ : InMux
    port map (
            O => \N__33984\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__6454\ : InMux
    port map (
            O => \N__33981\,
            I => \N__33978\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__33978\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNITOIN1Z0Z_28\
        );

    \I__6452\ : CascadeMux
    port map (
            O => \N__33975\,
            I => \N__33971\
        );

    \I__6451\ : InMux
    port map (
            O => \N__33974\,
            I => \N__33968\
        );

    \I__6450\ : InMux
    port map (
            O => \N__33971\,
            I => \N__33965\
        );

    \I__6449\ : LocalMux
    port map (
            O => \N__33968\,
            I => \N__33962\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__33965\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__6447\ : Odrv4
    port map (
            O => \N__33962\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__6446\ : InMux
    port map (
            O => \N__33957\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__6445\ : InMux
    port map (
            O => \N__33954\,
            I => \N__33950\
        );

    \I__6444\ : InMux
    port map (
            O => \N__33953\,
            I => \N__33947\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__33950\,
            I => \N__33944\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__33947\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__6441\ : Odrv4
    port map (
            O => \N__33944\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__6440\ : InMux
    port map (
            O => \N__33939\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__6439\ : InMux
    port map (
            O => \N__33936\,
            I => \N__33932\
        );

    \I__6438\ : InMux
    port map (
            O => \N__33935\,
            I => \N__33929\
        );

    \I__6437\ : LocalMux
    port map (
            O => \N__33932\,
            I => \N__33926\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__33929\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__6435\ : Odrv4
    port map (
            O => \N__33926\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__6434\ : InMux
    port map (
            O => \N__33921\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__6433\ : InMux
    port map (
            O => \N__33918\,
            I => \N__33914\
        );

    \I__6432\ : InMux
    port map (
            O => \N__33917\,
            I => \N__33911\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__33914\,
            I => \N__33908\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__33911\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__6429\ : Odrv4
    port map (
            O => \N__33908\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__6428\ : InMux
    port map (
            O => \N__33903\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__6427\ : InMux
    port map (
            O => \N__33900\,
            I => \N__33896\
        );

    \I__6426\ : InMux
    port map (
            O => \N__33899\,
            I => \N__33893\
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__33896\,
            I => \N__33890\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__33893\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__6423\ : Odrv12
    port map (
            O => \N__33890\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__6422\ : InMux
    port map (
            O => \N__33885\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__6421\ : InMux
    port map (
            O => \N__33882\,
            I => \N__33879\
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__33879\,
            I => \N__33875\
        );

    \I__6419\ : InMux
    port map (
            O => \N__33878\,
            I => \N__33872\
        );

    \I__6418\ : Span4Mux_v
    port map (
            O => \N__33875\,
            I => \N__33869\
        );

    \I__6417\ : LocalMux
    port map (
            O => \N__33872\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__6416\ : Odrv4
    port map (
            O => \N__33869\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__6415\ : InMux
    port map (
            O => \N__33864\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__6414\ : InMux
    port map (
            O => \N__33861\,
            I => \N__33858\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__33858\,
            I => \N__33854\
        );

    \I__6412\ : InMux
    port map (
            O => \N__33857\,
            I => \N__33851\
        );

    \I__6411\ : Span4Mux_v
    port map (
            O => \N__33854\,
            I => \N__33848\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__33851\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__6409\ : Odrv4
    port map (
            O => \N__33848\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__6408\ : InMux
    port map (
            O => \N__33843\,
            I => \bfn_12_18_0_\
        );

    \I__6407\ : InMux
    port map (
            O => \N__33840\,
            I => \N__33837\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__33837\,
            I => \N__33834\
        );

    \I__6405\ : Odrv4
    port map (
            O => \N__33834\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt18\
        );

    \I__6404\ : CascadeMux
    port map (
            O => \N__33831\,
            I => \N__33828\
        );

    \I__6403\ : InMux
    port map (
            O => \N__33828\,
            I => \N__33825\
        );

    \I__6402\ : LocalMux
    port map (
            O => \N__33825\,
            I => \N__33822\
        );

    \I__6401\ : Odrv12
    port map (
            O => \N__33822\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\
        );

    \I__6400\ : CascadeMux
    port map (
            O => \N__33819\,
            I => \N__33816\
        );

    \I__6399\ : InMux
    port map (
            O => \N__33816\,
            I => \N__33813\
        );

    \I__6398\ : LocalMux
    port map (
            O => \N__33813\,
            I => \N__33810\
        );

    \I__6397\ : Odrv12
    port map (
            O => \N__33810\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO\
        );

    \I__6396\ : InMux
    port map (
            O => \N__33807\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_28\
        );

    \I__6395\ : InMux
    port map (
            O => \N__33804\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30\
        );

    \I__6394\ : InMux
    port map (
            O => \N__33801\,
            I => \N__33795\
        );

    \I__6393\ : InMux
    port map (
            O => \N__33800\,
            I => \N__33795\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__33795\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__6391\ : CascadeMux
    port map (
            O => \N__33792\,
            I => \N__33788\
        );

    \I__6390\ : InMux
    port map (
            O => \N__33791\,
            I => \N__33785\
        );

    \I__6389\ : InMux
    port map (
            O => \N__33788\,
            I => \N__33781\
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__33785\,
            I => \N__33778\
        );

    \I__6387\ : InMux
    port map (
            O => \N__33784\,
            I => \N__33775\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__33781\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__6385\ : Odrv4
    port map (
            O => \N__33778\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__6384\ : LocalMux
    port map (
            O => \N__33775\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__6383\ : InMux
    port map (
            O => \N__33768\,
            I => \N__33765\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__33765\,
            I => \N__33762\
        );

    \I__6381\ : Span4Mux_h
    port map (
            O => \N__33762\,
            I => \N__33759\
        );

    \I__6380\ : Odrv4
    port map (
            O => \N__33759\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\
        );

    \I__6379\ : CascadeMux
    port map (
            O => \N__33756\,
            I => \N__33753\
        );

    \I__6378\ : InMux
    port map (
            O => \N__33753\,
            I => \N__33750\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__33750\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\
        );

    \I__6376\ : InMux
    port map (
            O => \N__33747\,
            I => \N__33744\
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__33744\,
            I => \N__33741\
        );

    \I__6374\ : Odrv4
    port map (
            O => \N__33741\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\
        );

    \I__6373\ : CascadeMux
    port map (
            O => \N__33738\,
            I => \N__33735\
        );

    \I__6372\ : InMux
    port map (
            O => \N__33735\,
            I => \N__33732\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__33732\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\
        );

    \I__6370\ : CascadeMux
    port map (
            O => \N__33729\,
            I => \N__33726\
        );

    \I__6369\ : InMux
    port map (
            O => \N__33726\,
            I => \N__33723\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__33723\,
            I => \N__33720\
        );

    \I__6367\ : Odrv4
    port map (
            O => \N__33720\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\
        );

    \I__6366\ : InMux
    port map (
            O => \N__33717\,
            I => \N__33714\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__33714\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\
        );

    \I__6364\ : InMux
    port map (
            O => \N__33711\,
            I => \N__33708\
        );

    \I__6363\ : LocalMux
    port map (
            O => \N__33708\,
            I => \N__33705\
        );

    \I__6362\ : Odrv4
    port map (
            O => \N__33705\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\
        );

    \I__6361\ : CascadeMux
    port map (
            O => \N__33702\,
            I => \N__33699\
        );

    \I__6360\ : InMux
    port map (
            O => \N__33699\,
            I => \N__33696\
        );

    \I__6359\ : LocalMux
    port map (
            O => \N__33696\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\
        );

    \I__6358\ : CascadeMux
    port map (
            O => \N__33693\,
            I => \N__33690\
        );

    \I__6357\ : InMux
    port map (
            O => \N__33690\,
            I => \N__33687\
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__33687\,
            I => \N__33684\
        );

    \I__6355\ : Odrv4
    port map (
            O => \N__33684\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\
        );

    \I__6354\ : InMux
    port map (
            O => \N__33681\,
            I => \N__33678\
        );

    \I__6353\ : LocalMux
    port map (
            O => \N__33678\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\
        );

    \I__6352\ : InMux
    port map (
            O => \N__33675\,
            I => \N__33672\
        );

    \I__6351\ : LocalMux
    port map (
            O => \N__33672\,
            I => \N__33669\
        );

    \I__6350\ : Span4Mux_h
    port map (
            O => \N__33669\,
            I => \N__33666\
        );

    \I__6349\ : Span4Mux_v
    port map (
            O => \N__33666\,
            I => \N__33663\
        );

    \I__6348\ : Odrv4
    port map (
            O => \N__33663\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\
        );

    \I__6347\ : CascadeMux
    port map (
            O => \N__33660\,
            I => \N__33657\
        );

    \I__6346\ : InMux
    port map (
            O => \N__33657\,
            I => \N__33654\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__33654\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\
        );

    \I__6344\ : InMux
    port map (
            O => \N__33651\,
            I => \N__33648\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__33648\,
            I => \N__33645\
        );

    \I__6342\ : Span4Mux_h
    port map (
            O => \N__33645\,
            I => \N__33642\
        );

    \I__6341\ : Odrv4
    port map (
            O => \N__33642\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\
        );

    \I__6340\ : CascadeMux
    port map (
            O => \N__33639\,
            I => \N__33636\
        );

    \I__6339\ : InMux
    port map (
            O => \N__33636\,
            I => \N__33633\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__33633\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\
        );

    \I__6337\ : InMux
    port map (
            O => \N__33630\,
            I => \N__33627\
        );

    \I__6336\ : LocalMux
    port map (
            O => \N__33627\,
            I => \N__33624\
        );

    \I__6335\ : Span4Mux_v
    port map (
            O => \N__33624\,
            I => \N__33621\
        );

    \I__6334\ : Odrv4
    port map (
            O => \N__33621\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt16\
        );

    \I__6333\ : CascadeMux
    port map (
            O => \N__33618\,
            I => \N__33615\
        );

    \I__6332\ : InMux
    port map (
            O => \N__33615\,
            I => \N__33612\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__33612\,
            I => \N__33609\
        );

    \I__6330\ : Span4Mux_v
    port map (
            O => \N__33609\,
            I => \N__33606\
        );

    \I__6329\ : Odrv4
    port map (
            O => \N__33606\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\
        );

    \I__6328\ : InMux
    port map (
            O => \N__33603\,
            I => \N__33600\
        );

    \I__6327\ : LocalMux
    port map (
            O => \N__33600\,
            I => \N__33597\
        );

    \I__6326\ : Odrv4
    port map (
            O => \N__33597\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\
        );

    \I__6325\ : CascadeMux
    port map (
            O => \N__33594\,
            I => \N__33591\
        );

    \I__6324\ : InMux
    port map (
            O => \N__33591\,
            I => \N__33588\
        );

    \I__6323\ : LocalMux
    port map (
            O => \N__33588\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\
        );

    \I__6322\ : InMux
    port map (
            O => \N__33585\,
            I => \N__33582\
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__33582\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\
        );

    \I__6320\ : CascadeMux
    port map (
            O => \N__33579\,
            I => \N__33576\
        );

    \I__6319\ : InMux
    port map (
            O => \N__33576\,
            I => \N__33573\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__33573\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\
        );

    \I__6317\ : InMux
    port map (
            O => \N__33570\,
            I => \N__33567\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__33567\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\
        );

    \I__6315\ : CascadeMux
    port map (
            O => \N__33564\,
            I => \N__33561\
        );

    \I__6314\ : InMux
    port map (
            O => \N__33561\,
            I => \N__33558\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__33558\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\
        );

    \I__6312\ : InMux
    port map (
            O => \N__33555\,
            I => \N__33552\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__33552\,
            I => \N__33549\
        );

    \I__6310\ : Odrv4
    port map (
            O => \N__33549\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\
        );

    \I__6309\ : CascadeMux
    port map (
            O => \N__33546\,
            I => \N__33543\
        );

    \I__6308\ : InMux
    port map (
            O => \N__33543\,
            I => \N__33540\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__33540\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\
        );

    \I__6306\ : InMux
    port map (
            O => \N__33537\,
            I => \N__33534\
        );

    \I__6305\ : LocalMux
    port map (
            O => \N__33534\,
            I => \N__33531\
        );

    \I__6304\ : Span4Mux_h
    port map (
            O => \N__33531\,
            I => \N__33528\
        );

    \I__6303\ : Span4Mux_h
    port map (
            O => \N__33528\,
            I => \N__33525\
        );

    \I__6302\ : Odrv4
    port map (
            O => \N__33525\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\
        );

    \I__6301\ : CascadeMux
    port map (
            O => \N__33522\,
            I => \N__33519\
        );

    \I__6300\ : InMux
    port map (
            O => \N__33519\,
            I => \N__33516\
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__33516\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\
        );

    \I__6298\ : CascadeMux
    port map (
            O => \N__33513\,
            I => \N__33510\
        );

    \I__6297\ : InMux
    port map (
            O => \N__33510\,
            I => \N__33507\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__33507\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\
        );

    \I__6295\ : InMux
    port map (
            O => \N__33504\,
            I => \N__33501\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__33501\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\
        );

    \I__6293\ : InMux
    port map (
            O => \N__33498\,
            I => \N__33495\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__33495\,
            I => \N__33492\
        );

    \I__6291\ : Span4Mux_h
    port map (
            O => \N__33492\,
            I => \N__33489\
        );

    \I__6290\ : Span4Mux_v
    port map (
            O => \N__33489\,
            I => \N__33486\
        );

    \I__6289\ : Odrv4
    port map (
            O => \N__33486\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\
        );

    \I__6288\ : CascadeMux
    port map (
            O => \N__33483\,
            I => \N__33480\
        );

    \I__6287\ : InMux
    port map (
            O => \N__33480\,
            I => \N__33477\
        );

    \I__6286\ : LocalMux
    port map (
            O => \N__33477\,
            I => \N__33474\
        );

    \I__6285\ : Odrv4
    port map (
            O => \N__33474\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\
        );

    \I__6284\ : InMux
    port map (
            O => \N__33471\,
            I => \N__33468\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__33468\,
            I => \N__33465\
        );

    \I__6282\ : Span4Mux_v
    port map (
            O => \N__33465\,
            I => \N__33462\
        );

    \I__6281\ : Odrv4
    port map (
            O => \N__33462\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\
        );

    \I__6280\ : CascadeMux
    port map (
            O => \N__33459\,
            I => \N__33456\
        );

    \I__6279\ : InMux
    port map (
            O => \N__33456\,
            I => \N__33453\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__33453\,
            I => \N__33450\
        );

    \I__6277\ : Odrv4
    port map (
            O => \N__33450\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\
        );

    \I__6276\ : InMux
    port map (
            O => \N__33447\,
            I => \N__33444\
        );

    \I__6275\ : LocalMux
    port map (
            O => \N__33444\,
            I => \N__33440\
        );

    \I__6274\ : InMux
    port map (
            O => \N__33443\,
            I => \N__33437\
        );

    \I__6273\ : Span4Mux_v
    port map (
            O => \N__33440\,
            I => \N__33432\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__33437\,
            I => \N__33432\
        );

    \I__6271\ : Span4Mux_h
    port map (
            O => \N__33432\,
            I => \N__33428\
        );

    \I__6270\ : InMux
    port map (
            O => \N__33431\,
            I => \N__33425\
        );

    \I__6269\ : Odrv4
    port map (
            O => \N__33428\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__33425\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__6267\ : InMux
    port map (
            O => \N__33420\,
            I => \N__33417\
        );

    \I__6266\ : LocalMux
    port map (
            O => \N__33417\,
            I => \N__33414\
        );

    \I__6265\ : Span4Mux_v
    port map (
            O => \N__33414\,
            I => \N__33411\
        );

    \I__6264\ : Odrv4
    port map (
            O => \N__33411\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\
        );

    \I__6263\ : InMux
    port map (
            O => \N__33408\,
            I => \N__33405\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__33405\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\
        );

    \I__6261\ : CascadeMux
    port map (
            O => \N__33402\,
            I => \N__33399\
        );

    \I__6260\ : InMux
    port map (
            O => \N__33399\,
            I => \N__33396\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__33396\,
            I => \N__33393\
        );

    \I__6258\ : Odrv4
    port map (
            O => \N__33393\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\
        );

    \I__6257\ : CascadeMux
    port map (
            O => \N__33390\,
            I => \N__33387\
        );

    \I__6256\ : InMux
    port map (
            O => \N__33387\,
            I => \N__33384\
        );

    \I__6255\ : LocalMux
    port map (
            O => \N__33384\,
            I => \N__33381\
        );

    \I__6254\ : Span4Mux_h
    port map (
            O => \N__33381\,
            I => \N__33376\
        );

    \I__6253\ : InMux
    port map (
            O => \N__33380\,
            I => \N__33371\
        );

    \I__6252\ : InMux
    port map (
            O => \N__33379\,
            I => \N__33371\
        );

    \I__6251\ : Odrv4
    port map (
            O => \N__33376\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__33371\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__6249\ : InMux
    port map (
            O => \N__33366\,
            I => \N__33363\
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__33363\,
            I => \N__33360\
        );

    \I__6247\ : Span4Mux_h
    port map (
            O => \N__33360\,
            I => \N__33357\
        );

    \I__6246\ : Span4Mux_h
    port map (
            O => \N__33357\,
            I => \N__33354\
        );

    \I__6245\ : Odrv4
    port map (
            O => \N__33354\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__6244\ : InMux
    port map (
            O => \N__33351\,
            I => \N__33348\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__33348\,
            I => \N__33344\
        );

    \I__6242\ : InMux
    port map (
            O => \N__33347\,
            I => \N__33341\
        );

    \I__6241\ : Span12Mux_s10_v
    port map (
            O => \N__33344\,
            I => \N__33335\
        );

    \I__6240\ : LocalMux
    port map (
            O => \N__33341\,
            I => \N__33335\
        );

    \I__6239\ : InMux
    port map (
            O => \N__33340\,
            I => \N__33332\
        );

    \I__6238\ : Odrv12
    port map (
            O => \N__33335\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__33332\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__6236\ : InMux
    port map (
            O => \N__33327\,
            I => \N__33324\
        );

    \I__6235\ : LocalMux
    port map (
            O => \N__33324\,
            I => \N__33321\
        );

    \I__6234\ : Span4Mux_h
    port map (
            O => \N__33321\,
            I => \N__33318\
        );

    \I__6233\ : Odrv4
    port map (
            O => \N__33318\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\
        );

    \I__6232\ : CascadeMux
    port map (
            O => \N__33315\,
            I => \N__33311\
        );

    \I__6231\ : InMux
    port map (
            O => \N__33314\,
            I => \N__33301\
        );

    \I__6230\ : InMux
    port map (
            O => \N__33311\,
            I => \N__33301\
        );

    \I__6229\ : InMux
    port map (
            O => \N__33310\,
            I => \N__33298\
        );

    \I__6228\ : CascadeMux
    port map (
            O => \N__33309\,
            I => \N__33295\
        );

    \I__6227\ : InMux
    port map (
            O => \N__33308\,
            I => \N__33288\
        );

    \I__6226\ : InMux
    port map (
            O => \N__33307\,
            I => \N__33283\
        );

    \I__6225\ : InMux
    port map (
            O => \N__33306\,
            I => \N__33283\
        );

    \I__6224\ : LocalMux
    port map (
            O => \N__33301\,
            I => \N__33278\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__33298\,
            I => \N__33278\
        );

    \I__6222\ : InMux
    port map (
            O => \N__33295\,
            I => \N__33275\
        );

    \I__6221\ : InMux
    port map (
            O => \N__33294\,
            I => \N__33270\
        );

    \I__6220\ : InMux
    port map (
            O => \N__33293\,
            I => \N__33270\
        );

    \I__6219\ : InMux
    port map (
            O => \N__33292\,
            I => \N__33267\
        );

    \I__6218\ : InMux
    port map (
            O => \N__33291\,
            I => \N__33264\
        );

    \I__6217\ : LocalMux
    port map (
            O => \N__33288\,
            I => \N__33257\
        );

    \I__6216\ : LocalMux
    port map (
            O => \N__33283\,
            I => \N__33257\
        );

    \I__6215\ : Span4Mux_v
    port map (
            O => \N__33278\,
            I => \N__33257\
        );

    \I__6214\ : LocalMux
    port map (
            O => \N__33275\,
            I => \N__33252\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__33270\,
            I => \N__33252\
        );

    \I__6212\ : LocalMux
    port map (
            O => \N__33267\,
            I => \phase_controller_inst1.stoper_hc.N_328\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__33264\,
            I => \phase_controller_inst1.stoper_hc.N_328\
        );

    \I__6210\ : Odrv4
    port map (
            O => \N__33257\,
            I => \phase_controller_inst1.stoper_hc.N_328\
        );

    \I__6209\ : Odrv4
    port map (
            O => \N__33252\,
            I => \phase_controller_inst1.stoper_hc.N_328\
        );

    \I__6208\ : InMux
    port map (
            O => \N__33243\,
            I => \N__33231\
        );

    \I__6207\ : InMux
    port map (
            O => \N__33242\,
            I => \N__33216\
        );

    \I__6206\ : InMux
    port map (
            O => \N__33241\,
            I => \N__33216\
        );

    \I__6205\ : InMux
    port map (
            O => \N__33240\,
            I => \N__33216\
        );

    \I__6204\ : InMux
    port map (
            O => \N__33239\,
            I => \N__33213\
        );

    \I__6203\ : InMux
    port map (
            O => \N__33238\,
            I => \N__33204\
        );

    \I__6202\ : InMux
    port map (
            O => \N__33237\,
            I => \N__33204\
        );

    \I__6201\ : InMux
    port map (
            O => \N__33236\,
            I => \N__33204\
        );

    \I__6200\ : InMux
    port map (
            O => \N__33235\,
            I => \N__33204\
        );

    \I__6199\ : InMux
    port map (
            O => \N__33234\,
            I => \N__33199\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__33231\,
            I => \N__33196\
        );

    \I__6197\ : InMux
    port map (
            O => \N__33230\,
            I => \N__33191\
        );

    \I__6196\ : InMux
    port map (
            O => \N__33229\,
            I => \N__33191\
        );

    \I__6195\ : InMux
    port map (
            O => \N__33228\,
            I => \N__33167\
        );

    \I__6194\ : InMux
    port map (
            O => \N__33227\,
            I => \N__33167\
        );

    \I__6193\ : InMux
    port map (
            O => \N__33226\,
            I => \N__33167\
        );

    \I__6192\ : InMux
    port map (
            O => \N__33225\,
            I => \N__33167\
        );

    \I__6191\ : InMux
    port map (
            O => \N__33224\,
            I => \N__33167\
        );

    \I__6190\ : InMux
    port map (
            O => \N__33223\,
            I => \N__33167\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__33216\,
            I => \N__33164\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__33213\,
            I => \N__33159\
        );

    \I__6187\ : LocalMux
    port map (
            O => \N__33204\,
            I => \N__33159\
        );

    \I__6186\ : InMux
    port map (
            O => \N__33203\,
            I => \N__33154\
        );

    \I__6185\ : InMux
    port map (
            O => \N__33202\,
            I => \N__33154\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__33199\,
            I => \N__33151\
        );

    \I__6183\ : Span4Mux_v
    port map (
            O => \N__33196\,
            I => \N__33146\
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__33191\,
            I => \N__33146\
        );

    \I__6181\ : InMux
    port map (
            O => \N__33190\,
            I => \N__33135\
        );

    \I__6180\ : InMux
    port map (
            O => \N__33189\,
            I => \N__33135\
        );

    \I__6179\ : InMux
    port map (
            O => \N__33188\,
            I => \N__33135\
        );

    \I__6178\ : InMux
    port map (
            O => \N__33187\,
            I => \N__33135\
        );

    \I__6177\ : InMux
    port map (
            O => \N__33186\,
            I => \N__33135\
        );

    \I__6176\ : InMux
    port map (
            O => \N__33185\,
            I => \N__33132\
        );

    \I__6175\ : InMux
    port map (
            O => \N__33184\,
            I => \N__33127\
        );

    \I__6174\ : InMux
    port map (
            O => \N__33183\,
            I => \N__33127\
        );

    \I__6173\ : InMux
    port map (
            O => \N__33182\,
            I => \N__33122\
        );

    \I__6172\ : InMux
    port map (
            O => \N__33181\,
            I => \N__33122\
        );

    \I__6171\ : CascadeMux
    port map (
            O => \N__33180\,
            I => \N__33114\
        );

    \I__6170\ : LocalMux
    port map (
            O => \N__33167\,
            I => \N__33107\
        );

    \I__6169\ : Span4Mux_v
    port map (
            O => \N__33164\,
            I => \N__33107\
        );

    \I__6168\ : Span4Mux_v
    port map (
            O => \N__33159\,
            I => \N__33107\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__33154\,
            I => \N__33104\
        );

    \I__6166\ : Span4Mux_v
    port map (
            O => \N__33151\,
            I => \N__33101\
        );

    \I__6165\ : Span4Mux_h
    port map (
            O => \N__33146\,
            I => \N__33098\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__33135\,
            I => \N__33095\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__33132\,
            I => \N__33088\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__33127\,
            I => \N__33088\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__33122\,
            I => \N__33088\
        );

    \I__6160\ : InMux
    port map (
            O => \N__33121\,
            I => \N__33085\
        );

    \I__6159\ : InMux
    port map (
            O => \N__33120\,
            I => \N__33078\
        );

    \I__6158\ : InMux
    port map (
            O => \N__33119\,
            I => \N__33078\
        );

    \I__6157\ : InMux
    port map (
            O => \N__33118\,
            I => \N__33078\
        );

    \I__6156\ : InMux
    port map (
            O => \N__33117\,
            I => \N__33073\
        );

    \I__6155\ : InMux
    port map (
            O => \N__33114\,
            I => \N__33073\
        );

    \I__6154\ : Sp12to4
    port map (
            O => \N__33107\,
            I => \N__33070\
        );

    \I__6153\ : Span4Mux_h
    port map (
            O => \N__33104\,
            I => \N__33067\
        );

    \I__6152\ : Span4Mux_h
    port map (
            O => \N__33101\,
            I => \N__33062\
        );

    \I__6151\ : Span4Mux_v
    port map (
            O => \N__33098\,
            I => \N__33062\
        );

    \I__6150\ : Span4Mux_v
    port map (
            O => \N__33095\,
            I => \N__33057\
        );

    \I__6149\ : Span4Mux_v
    port map (
            O => \N__33088\,
            I => \N__33057\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__33085\,
            I => \elapsed_time_ns_1_RNI5IV8E1_0_31\
        );

    \I__6147\ : LocalMux
    port map (
            O => \N__33078\,
            I => \elapsed_time_ns_1_RNI5IV8E1_0_31\
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__33073\,
            I => \elapsed_time_ns_1_RNI5IV8E1_0_31\
        );

    \I__6145\ : Odrv12
    port map (
            O => \N__33070\,
            I => \elapsed_time_ns_1_RNI5IV8E1_0_31\
        );

    \I__6144\ : Odrv4
    port map (
            O => \N__33067\,
            I => \elapsed_time_ns_1_RNI5IV8E1_0_31\
        );

    \I__6143\ : Odrv4
    port map (
            O => \N__33062\,
            I => \elapsed_time_ns_1_RNI5IV8E1_0_31\
        );

    \I__6142\ : Odrv4
    port map (
            O => \N__33057\,
            I => \elapsed_time_ns_1_RNI5IV8E1_0_31\
        );

    \I__6141\ : CascadeMux
    port map (
            O => \N__33042\,
            I => \N__33037\
        );

    \I__6140\ : CascadeMux
    port map (
            O => \N__33041\,
            I => \N__33031\
        );

    \I__6139\ : InMux
    port map (
            O => \N__33040\,
            I => \N__33026\
        );

    \I__6138\ : InMux
    port map (
            O => \N__33037\,
            I => \N__33026\
        );

    \I__6137\ : InMux
    port map (
            O => \N__33036\,
            I => \N__33023\
        );

    \I__6136\ : InMux
    port map (
            O => \N__33035\,
            I => \N__33020\
        );

    \I__6135\ : CascadeMux
    port map (
            O => \N__33034\,
            I => \N__33015\
        );

    \I__6134\ : InMux
    port map (
            O => \N__33031\,
            I => \N__33012\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__33026\,
            I => \N__33007\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__33023\,
            I => \N__33007\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__33020\,
            I => \N__33004\
        );

    \I__6130\ : CascadeMux
    port map (
            O => \N__33019\,
            I => \N__33000\
        );

    \I__6129\ : InMux
    port map (
            O => \N__33018\,
            I => \N__32992\
        );

    \I__6128\ : InMux
    port map (
            O => \N__33015\,
            I => \N__32989\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__33012\,
            I => \N__32986\
        );

    \I__6126\ : Span4Mux_h
    port map (
            O => \N__33007\,
            I => \N__32983\
        );

    \I__6125\ : Span4Mux_v
    port map (
            O => \N__33004\,
            I => \N__32980\
        );

    \I__6124\ : InMux
    port map (
            O => \N__33003\,
            I => \N__32977\
        );

    \I__6123\ : InMux
    port map (
            O => \N__33000\,
            I => \N__32974\
        );

    \I__6122\ : InMux
    port map (
            O => \N__32999\,
            I => \N__32971\
        );

    \I__6121\ : InMux
    port map (
            O => \N__32998\,
            I => \N__32968\
        );

    \I__6120\ : InMux
    port map (
            O => \N__32997\,
            I => \N__32961\
        );

    \I__6119\ : InMux
    port map (
            O => \N__32996\,
            I => \N__32961\
        );

    \I__6118\ : InMux
    port map (
            O => \N__32995\,
            I => \N__32961\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__32992\,
            I => \N__32958\
        );

    \I__6116\ : LocalMux
    port map (
            O => \N__32989\,
            I => \N__32949\
        );

    \I__6115\ : Span4Mux_v
    port map (
            O => \N__32986\,
            I => \N__32949\
        );

    \I__6114\ : Span4Mux_v
    port map (
            O => \N__32983\,
            I => \N__32949\
        );

    \I__6113\ : Span4Mux_h
    port map (
            O => \N__32980\,
            I => \N__32949\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__32977\,
            I => \phase_controller_inst1.stoper_hc.N_326\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__32974\,
            I => \phase_controller_inst1.stoper_hc.N_326\
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__32971\,
            I => \phase_controller_inst1.stoper_hc.N_326\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__32968\,
            I => \phase_controller_inst1.stoper_hc.N_326\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__32961\,
            I => \phase_controller_inst1.stoper_hc.N_326\
        );

    \I__6107\ : Odrv12
    port map (
            O => \N__32958\,
            I => \phase_controller_inst1.stoper_hc.N_326\
        );

    \I__6106\ : Odrv4
    port map (
            O => \N__32949\,
            I => \phase_controller_inst1.stoper_hc.N_326\
        );

    \I__6105\ : InMux
    port map (
            O => \N__32934\,
            I => \N__32931\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__32931\,
            I => \N__32927\
        );

    \I__6103\ : InMux
    port map (
            O => \N__32930\,
            I => \N__32924\
        );

    \I__6102\ : Odrv4
    port map (
            O => \N__32927\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2\
        );

    \I__6101\ : LocalMux
    port map (
            O => \N__32924\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2\
        );

    \I__6100\ : InMux
    port map (
            O => \N__32919\,
            I => \N__32916\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__32916\,
            I => \N__32913\
        );

    \I__6098\ : Span4Mux_v
    port map (
            O => \N__32913\,
            I => \N__32910\
        );

    \I__6097\ : Span4Mux_h
    port map (
            O => \N__32910\,
            I => \N__32907\
        );

    \I__6096\ : Span4Mux_v
    port map (
            O => \N__32907\,
            I => \N__32904\
        );

    \I__6095\ : Odrv4
    port map (
            O => \N__32904\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\
        );

    \I__6094\ : CEMux
    port map (
            O => \N__32901\,
            I => \N__32893\
        );

    \I__6093\ : CEMux
    port map (
            O => \N__32900\,
            I => \N__32890\
        );

    \I__6092\ : CEMux
    port map (
            O => \N__32899\,
            I => \N__32886\
        );

    \I__6091\ : CEMux
    port map (
            O => \N__32898\,
            I => \N__32883\
        );

    \I__6090\ : CEMux
    port map (
            O => \N__32897\,
            I => \N__32880\
        );

    \I__6089\ : CEMux
    port map (
            O => \N__32896\,
            I => \N__32876\
        );

    \I__6088\ : LocalMux
    port map (
            O => \N__32893\,
            I => \N__32873\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__32890\,
            I => \N__32870\
        );

    \I__6086\ : CEMux
    port map (
            O => \N__32889\,
            I => \N__32867\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__32886\,
            I => \N__32841\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__32883\,
            I => \N__32838\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__32880\,
            I => \N__32835\
        );

    \I__6082\ : CEMux
    port map (
            O => \N__32879\,
            I => \N__32832\
        );

    \I__6081\ : LocalMux
    port map (
            O => \N__32876\,
            I => \N__32827\
        );

    \I__6080\ : Span4Mux_v
    port map (
            O => \N__32873\,
            I => \N__32827\
        );

    \I__6079\ : Span4Mux_h
    port map (
            O => \N__32870\,
            I => \N__32824\
        );

    \I__6078\ : LocalMux
    port map (
            O => \N__32867\,
            I => \N__32821\
        );

    \I__6077\ : InMux
    port map (
            O => \N__32866\,
            I => \N__32812\
        );

    \I__6076\ : InMux
    port map (
            O => \N__32865\,
            I => \N__32812\
        );

    \I__6075\ : InMux
    port map (
            O => \N__32864\,
            I => \N__32812\
        );

    \I__6074\ : InMux
    port map (
            O => \N__32863\,
            I => \N__32812\
        );

    \I__6073\ : InMux
    port map (
            O => \N__32862\,
            I => \N__32803\
        );

    \I__6072\ : InMux
    port map (
            O => \N__32861\,
            I => \N__32803\
        );

    \I__6071\ : InMux
    port map (
            O => \N__32860\,
            I => \N__32803\
        );

    \I__6070\ : InMux
    port map (
            O => \N__32859\,
            I => \N__32803\
        );

    \I__6069\ : InMux
    port map (
            O => \N__32858\,
            I => \N__32794\
        );

    \I__6068\ : InMux
    port map (
            O => \N__32857\,
            I => \N__32794\
        );

    \I__6067\ : InMux
    port map (
            O => \N__32856\,
            I => \N__32794\
        );

    \I__6066\ : InMux
    port map (
            O => \N__32855\,
            I => \N__32794\
        );

    \I__6065\ : InMux
    port map (
            O => \N__32854\,
            I => \N__32785\
        );

    \I__6064\ : InMux
    port map (
            O => \N__32853\,
            I => \N__32785\
        );

    \I__6063\ : InMux
    port map (
            O => \N__32852\,
            I => \N__32785\
        );

    \I__6062\ : InMux
    port map (
            O => \N__32851\,
            I => \N__32785\
        );

    \I__6061\ : InMux
    port map (
            O => \N__32850\,
            I => \N__32778\
        );

    \I__6060\ : InMux
    port map (
            O => \N__32849\,
            I => \N__32778\
        );

    \I__6059\ : InMux
    port map (
            O => \N__32848\,
            I => \N__32778\
        );

    \I__6058\ : InMux
    port map (
            O => \N__32847\,
            I => \N__32769\
        );

    \I__6057\ : InMux
    port map (
            O => \N__32846\,
            I => \N__32769\
        );

    \I__6056\ : InMux
    port map (
            O => \N__32845\,
            I => \N__32769\
        );

    \I__6055\ : InMux
    port map (
            O => \N__32844\,
            I => \N__32769\
        );

    \I__6054\ : Span4Mux_v
    port map (
            O => \N__32841\,
            I => \N__32766\
        );

    \I__6053\ : Span4Mux_v
    port map (
            O => \N__32838\,
            I => \N__32751\
        );

    \I__6052\ : Span4Mux_v
    port map (
            O => \N__32835\,
            I => \N__32751\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__32832\,
            I => \N__32751\
        );

    \I__6050\ : Span4Mux_h
    port map (
            O => \N__32827\,
            I => \N__32746\
        );

    \I__6049\ : Span4Mux_v
    port map (
            O => \N__32824\,
            I => \N__32746\
        );

    \I__6048\ : Span4Mux_v
    port map (
            O => \N__32821\,
            I => \N__32743\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__32812\,
            I => \N__32730\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__32803\,
            I => \N__32730\
        );

    \I__6045\ : LocalMux
    port map (
            O => \N__32794\,
            I => \N__32730\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__32785\,
            I => \N__32730\
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__32778\,
            I => \N__32730\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__32769\,
            I => \N__32730\
        );

    \I__6041\ : Span4Mux_v
    port map (
            O => \N__32766\,
            I => \N__32727\
        );

    \I__6040\ : InMux
    port map (
            O => \N__32765\,
            I => \N__32724\
        );

    \I__6039\ : InMux
    port map (
            O => \N__32764\,
            I => \N__32717\
        );

    \I__6038\ : InMux
    port map (
            O => \N__32763\,
            I => \N__32717\
        );

    \I__6037\ : InMux
    port map (
            O => \N__32762\,
            I => \N__32717\
        );

    \I__6036\ : InMux
    port map (
            O => \N__32761\,
            I => \N__32708\
        );

    \I__6035\ : InMux
    port map (
            O => \N__32760\,
            I => \N__32708\
        );

    \I__6034\ : InMux
    port map (
            O => \N__32759\,
            I => \N__32708\
        );

    \I__6033\ : InMux
    port map (
            O => \N__32758\,
            I => \N__32708\
        );

    \I__6032\ : Span4Mux_v
    port map (
            O => \N__32751\,
            I => \N__32703\
        );

    \I__6031\ : Span4Mux_v
    port map (
            O => \N__32746\,
            I => \N__32703\
        );

    \I__6030\ : Span4Mux_h
    port map (
            O => \N__32743\,
            I => \N__32696\
        );

    \I__6029\ : Span4Mux_v
    port map (
            O => \N__32730\,
            I => \N__32696\
        );

    \I__6028\ : Span4Mux_h
    port map (
            O => \N__32727\,
            I => \N__32696\
        );

    \I__6027\ : LocalMux
    port map (
            O => \N__32724\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__32717\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__32708\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__6024\ : Odrv4
    port map (
            O => \N__32703\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__6023\ : Odrv4
    port map (
            O => \N__32696\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__6022\ : InMux
    port map (
            O => \N__32685\,
            I => \N__32682\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__32682\,
            I => \N__32678\
        );

    \I__6020\ : InMux
    port map (
            O => \N__32681\,
            I => \N__32675\
        );

    \I__6019\ : Span4Mux_h
    port map (
            O => \N__32678\,
            I => \N__32670\
        );

    \I__6018\ : LocalMux
    port map (
            O => \N__32675\,
            I => \N__32670\
        );

    \I__6017\ : Span4Mux_h
    port map (
            O => \N__32670\,
            I => \N__32666\
        );

    \I__6016\ : InMux
    port map (
            O => \N__32669\,
            I => \N__32663\
        );

    \I__6015\ : Odrv4
    port map (
            O => \N__32666\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__6014\ : LocalMux
    port map (
            O => \N__32663\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__6013\ : InMux
    port map (
            O => \N__32658\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_5\
        );

    \I__6012\ : InMux
    port map (
            O => \N__32655\,
            I => \N__32651\
        );

    \I__6011\ : InMux
    port map (
            O => \N__32654\,
            I => \N__32647\
        );

    \I__6010\ : LocalMux
    port map (
            O => \N__32651\,
            I => \N__32644\
        );

    \I__6009\ : InMux
    port map (
            O => \N__32650\,
            I => \N__32641\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__32647\,
            I => \N__32638\
        );

    \I__6007\ : Span4Mux_h
    port map (
            O => \N__32644\,
            I => \N__32635\
        );

    \I__6006\ : LocalMux
    port map (
            O => \N__32641\,
            I => \N__32632\
        );

    \I__6005\ : Odrv12
    port map (
            O => \N__32638\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__6004\ : Odrv4
    port map (
            O => \N__32635\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__6003\ : Odrv4
    port map (
            O => \N__32632\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__6002\ : InMux
    port map (
            O => \N__32625\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_6\
        );

    \I__6001\ : InMux
    port map (
            O => \N__32622\,
            I => \bfn_12_11_0_\
        );

    \I__6000\ : InMux
    port map (
            O => \N__32619\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_8\
        );

    \I__5999\ : InMux
    port map (
            O => \N__32616\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_9\
        );

    \I__5998\ : CascadeMux
    port map (
            O => \N__32613\,
            I => \N__32609\
        );

    \I__5997\ : InMux
    port map (
            O => \N__32612\,
            I => \N__32606\
        );

    \I__5996\ : InMux
    port map (
            O => \N__32609\,
            I => \N__32603\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__32606\,
            I => \N__32600\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__32603\,
            I => \N__32596\
        );

    \I__5993\ : Span4Mux_v
    port map (
            O => \N__32600\,
            I => \N__32593\
        );

    \I__5992\ : InMux
    port map (
            O => \N__32599\,
            I => \N__32590\
        );

    \I__5991\ : Span4Mux_v
    port map (
            O => \N__32596\,
            I => \N__32587\
        );

    \I__5990\ : Span4Mux_h
    port map (
            O => \N__32593\,
            I => \N__32582\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__32590\,
            I => \N__32582\
        );

    \I__5988\ : Odrv4
    port map (
            O => \N__32587\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__5987\ : Odrv4
    port map (
            O => \N__32582\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__5986\ : InMux
    port map (
            O => \N__32577\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_10\
        );

    \I__5985\ : InMux
    port map (
            O => \N__32574\,
            I => \N__32570\
        );

    \I__5984\ : InMux
    port map (
            O => \N__32573\,
            I => \N__32567\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__32570\,
            I => \N__32563\
        );

    \I__5982\ : LocalMux
    port map (
            O => \N__32567\,
            I => \N__32560\
        );

    \I__5981\ : InMux
    port map (
            O => \N__32566\,
            I => \N__32557\
        );

    \I__5980\ : Span4Mux_h
    port map (
            O => \N__32563\,
            I => \N__32554\
        );

    \I__5979\ : Span4Mux_h
    port map (
            O => \N__32560\,
            I => \N__32549\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__32557\,
            I => \N__32549\
        );

    \I__5977\ : Odrv4
    port map (
            O => \N__32554\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__5976\ : Odrv4
    port map (
            O => \N__32549\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__5975\ : InMux
    port map (
            O => \N__32544\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_11\
        );

    \I__5974\ : InMux
    port map (
            O => \N__32541\,
            I => \N__32536\
        );

    \I__5973\ : InMux
    port map (
            O => \N__32540\,
            I => \N__32531\
        );

    \I__5972\ : InMux
    port map (
            O => \N__32539\,
            I => \N__32531\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__32536\,
            I => \N__32526\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__32531\,
            I => \N__32526\
        );

    \I__5969\ : Span4Mux_h
    port map (
            O => \N__32526\,
            I => \N__32523\
        );

    \I__5968\ : Odrv4
    port map (
            O => \N__32523\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__5967\ : InMux
    port map (
            O => \N__32520\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_12\
        );

    \I__5966\ : InMux
    port map (
            O => \N__32517\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_13\
        );

    \I__5965\ : InMux
    port map (
            O => \N__32514\,
            I => \N__32511\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__32511\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\
        );

    \I__5963\ : InMux
    port map (
            O => \N__32508\,
            I => \N__32504\
        );

    \I__5962\ : InMux
    port map (
            O => \N__32507\,
            I => \N__32500\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__32504\,
            I => \N__32497\
        );

    \I__5960\ : InMux
    port map (
            O => \N__32503\,
            I => \N__32494\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__32500\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\
        );

    \I__5958\ : Odrv12
    port map (
            O => \N__32497\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__32494\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\
        );

    \I__5956\ : InMux
    port map (
            O => \N__32487\,
            I => \N__32483\
        );

    \I__5955\ : InMux
    port map (
            O => \N__32486\,
            I => \N__32480\
        );

    \I__5954\ : LocalMux
    port map (
            O => \N__32483\,
            I => \N__32474\
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__32480\,
            I => \N__32474\
        );

    \I__5952\ : InMux
    port map (
            O => \N__32479\,
            I => \N__32471\
        );

    \I__5951\ : Odrv4
    port map (
            O => \N__32474\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__32471\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\
        );

    \I__5949\ : InMux
    port map (
            O => \N__32466\,
            I => \N__32463\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__32463\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axb_0\
        );

    \I__5947\ : InMux
    port map (
            O => \N__32460\,
            I => \N__32457\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__32457\,
            I => \N__32454\
        );

    \I__5945\ : Span4Mux_h
    port map (
            O => \N__32454\,
            I => \N__32450\
        );

    \I__5944\ : InMux
    port map (
            O => \N__32453\,
            I => \N__32447\
        );

    \I__5943\ : Span4Mux_h
    port map (
            O => \N__32450\,
            I => \N__32442\
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__32447\,
            I => \N__32442\
        );

    \I__5941\ : Odrv4
    port map (
            O => \N__32442\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__5940\ : InMux
    port map (
            O => \N__32439\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_0\
        );

    \I__5939\ : InMux
    port map (
            O => \N__32436\,
            I => \N__32433\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__32433\,
            I => \N__32430\
        );

    \I__5937\ : Span4Mux_v
    port map (
            O => \N__32430\,
            I => \N__32426\
        );

    \I__5936\ : InMux
    port map (
            O => \N__32429\,
            I => \N__32423\
        );

    \I__5935\ : Span4Mux_h
    port map (
            O => \N__32426\,
            I => \N__32418\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__32423\,
            I => \N__32418\
        );

    \I__5933\ : Odrv4
    port map (
            O => \N__32418\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__5932\ : InMux
    port map (
            O => \N__32415\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_1\
        );

    \I__5931\ : InMux
    port map (
            O => \N__32412\,
            I => \N__32409\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__32409\,
            I => \N__32405\
        );

    \I__5929\ : InMux
    port map (
            O => \N__32408\,
            I => \N__32402\
        );

    \I__5928\ : Span12Mux_h
    port map (
            O => \N__32405\,
            I => \N__32399\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__32402\,
            I => \N__32396\
        );

    \I__5926\ : Odrv12
    port map (
            O => \N__32399\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__5925\ : Odrv4
    port map (
            O => \N__32396\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__5924\ : InMux
    port map (
            O => \N__32391\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_2\
        );

    \I__5923\ : InMux
    port map (
            O => \N__32388\,
            I => \N__32385\
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__32385\,
            I => \N__32380\
        );

    \I__5921\ : InMux
    port map (
            O => \N__32384\,
            I => \N__32377\
        );

    \I__5920\ : InMux
    port map (
            O => \N__32383\,
            I => \N__32374\
        );

    \I__5919\ : Span4Mux_v
    port map (
            O => \N__32380\,
            I => \N__32367\
        );

    \I__5918\ : LocalMux
    port map (
            O => \N__32377\,
            I => \N__32367\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__32374\,
            I => \N__32367\
        );

    \I__5916\ : Span4Mux_h
    port map (
            O => \N__32367\,
            I => \N__32364\
        );

    \I__5915\ : Odrv4
    port map (
            O => \N__32364\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__5914\ : InMux
    port map (
            O => \N__32361\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_3\
        );

    \I__5913\ : InMux
    port map (
            O => \N__32358\,
            I => \N__32355\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__32355\,
            I => \N__32352\
        );

    \I__5911\ : Span4Mux_h
    port map (
            O => \N__32352\,
            I => \N__32348\
        );

    \I__5910\ : CascadeMux
    port map (
            O => \N__32351\,
            I => \N__32345\
        );

    \I__5909\ : Span4Mux_h
    port map (
            O => \N__32348\,
            I => \N__32341\
        );

    \I__5908\ : InMux
    port map (
            O => \N__32345\,
            I => \N__32336\
        );

    \I__5907\ : InMux
    port map (
            O => \N__32344\,
            I => \N__32336\
        );

    \I__5906\ : Odrv4
    port map (
            O => \N__32341\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__32336\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__5904\ : InMux
    port map (
            O => \N__32331\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_4\
        );

    \I__5903\ : InMux
    port map (
            O => \N__32328\,
            I => \N__32323\
        );

    \I__5902\ : InMux
    port map (
            O => \N__32327\,
            I => \N__32319\
        );

    \I__5901\ : InMux
    port map (
            O => \N__32326\,
            I => \N__32316\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__32323\,
            I => \N__32313\
        );

    \I__5899\ : CascadeMux
    port map (
            O => \N__32322\,
            I => \N__32309\
        );

    \I__5898\ : LocalMux
    port map (
            O => \N__32319\,
            I => \N__32306\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__32316\,
            I => \N__32303\
        );

    \I__5896\ : Span4Mux_v
    port map (
            O => \N__32313\,
            I => \N__32300\
        );

    \I__5895\ : InMux
    port map (
            O => \N__32312\,
            I => \N__32295\
        );

    \I__5894\ : InMux
    port map (
            O => \N__32309\,
            I => \N__32295\
        );

    \I__5893\ : Span4Mux_v
    port map (
            O => \N__32306\,
            I => \N__32292\
        );

    \I__5892\ : Odrv4
    port map (
            O => \N__32303\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__5891\ : Odrv4
    port map (
            O => \N__32300\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__32295\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__5889\ : Odrv4
    port map (
            O => \N__32292\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__5888\ : InMux
    port map (
            O => \N__32283\,
            I => \N__32280\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__32280\,
            I => \N__32277\
        );

    \I__5886\ : Span4Mux_h
    port map (
            O => \N__32277\,
            I => \N__32274\
        );

    \I__5885\ : Odrv4
    port map (
            O => \N__32274\,
            I => \current_shift_inst.PI_CTRL.integrator_i_17\
        );

    \I__5884\ : CascadeMux
    port map (
            O => \N__32271\,
            I => \N__32267\
        );

    \I__5883\ : InMux
    port map (
            O => \N__32270\,
            I => \N__32262\
        );

    \I__5882\ : InMux
    port map (
            O => \N__32267\,
            I => \N__32259\
        );

    \I__5881\ : CascadeMux
    port map (
            O => \N__32266\,
            I => \N__32255\
        );

    \I__5880\ : InMux
    port map (
            O => \N__32265\,
            I => \N__32252\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__32262\,
            I => \N__32249\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__32259\,
            I => \N__32246\
        );

    \I__5877\ : InMux
    port map (
            O => \N__32258\,
            I => \N__32241\
        );

    \I__5876\ : InMux
    port map (
            O => \N__32255\,
            I => \N__32241\
        );

    \I__5875\ : LocalMux
    port map (
            O => \N__32252\,
            I => \N__32238\
        );

    \I__5874\ : Span4Mux_h
    port map (
            O => \N__32249\,
            I => \N__32233\
        );

    \I__5873\ : Span4Mux_h
    port map (
            O => \N__32246\,
            I => \N__32233\
        );

    \I__5872\ : LocalMux
    port map (
            O => \N__32241\,
            I => \N__32230\
        );

    \I__5871\ : Span4Mux_h
    port map (
            O => \N__32238\,
            I => \N__32227\
        );

    \I__5870\ : Odrv4
    port map (
            O => \N__32233\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__5869\ : Odrv12
    port map (
            O => \N__32230\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__5868\ : Odrv4
    port map (
            O => \N__32227\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__5867\ : InMux
    port map (
            O => \N__32220\,
            I => \N__32217\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__32217\,
            I => \N__32214\
        );

    \I__5865\ : Span4Mux_h
    port map (
            O => \N__32214\,
            I => \N__32211\
        );

    \I__5864\ : Odrv4
    port map (
            O => \N__32211\,
            I => \current_shift_inst.PI_CTRL.integrator_i_18\
        );

    \I__5863\ : CascadeMux
    port map (
            O => \N__32208\,
            I => \N__32205\
        );

    \I__5862\ : InMux
    port map (
            O => \N__32205\,
            I => \N__32201\
        );

    \I__5861\ : CascadeMux
    port map (
            O => \N__32204\,
            I => \N__32198\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__32201\,
            I => \N__32194\
        );

    \I__5859\ : InMux
    port map (
            O => \N__32198\,
            I => \N__32191\
        );

    \I__5858\ : InMux
    port map (
            O => \N__32197\,
            I => \N__32188\
        );

    \I__5857\ : Span4Mux_h
    port map (
            O => \N__32194\,
            I => \N__32185\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__32191\,
            I => \N__32182\
        );

    \I__5855\ : LocalMux
    port map (
            O => \N__32188\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\
        );

    \I__5854\ : Odrv4
    port map (
            O => \N__32185\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\
        );

    \I__5853\ : Odrv4
    port map (
            O => \N__32182\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\
        );

    \I__5852\ : CascadeMux
    port map (
            O => \N__32175\,
            I => \N__32172\
        );

    \I__5851\ : InMux
    port map (
            O => \N__32172\,
            I => \N__32169\
        );

    \I__5850\ : LocalMux
    port map (
            O => \N__32169\,
            I => \N__32164\
        );

    \I__5849\ : InMux
    port map (
            O => \N__32168\,
            I => \N__32160\
        );

    \I__5848\ : CascadeMux
    port map (
            O => \N__32167\,
            I => \N__32157\
        );

    \I__5847\ : Span4Mux_h
    port map (
            O => \N__32164\,
            I => \N__32154\
        );

    \I__5846\ : InMux
    port map (
            O => \N__32163\,
            I => \N__32150\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__32160\,
            I => \N__32147\
        );

    \I__5844\ : InMux
    port map (
            O => \N__32157\,
            I => \N__32144\
        );

    \I__5843\ : Span4Mux_h
    port map (
            O => \N__32154\,
            I => \N__32141\
        );

    \I__5842\ : InMux
    port map (
            O => \N__32153\,
            I => \N__32138\
        );

    \I__5841\ : LocalMux
    port map (
            O => \N__32150\,
            I => \N__32135\
        );

    \I__5840\ : Odrv4
    port map (
            O => \N__32147\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__32144\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__5838\ : Odrv4
    port map (
            O => \N__32141\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__32138\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__5836\ : Odrv4
    port map (
            O => \N__32135\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__5835\ : InMux
    port map (
            O => \N__32124\,
            I => \N__32121\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__32121\,
            I => \N__32118\
        );

    \I__5833\ : Span4Mux_v
    port map (
            O => \N__32118\,
            I => \N__32115\
        );

    \I__5832\ : Odrv4
    port map (
            O => \N__32115\,
            I => \current_shift_inst.PI_CTRL.integrator_i_12\
        );

    \I__5831\ : CascadeMux
    port map (
            O => \N__32112\,
            I => \N__32109\
        );

    \I__5830\ : InMux
    port map (
            O => \N__32109\,
            I => \N__32105\
        );

    \I__5829\ : InMux
    port map (
            O => \N__32108\,
            I => \N__32102\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__32105\,
            I => \N__32099\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__32102\,
            I => \N__32096\
        );

    \I__5826\ : Span4Mux_v
    port map (
            O => \N__32099\,
            I => \N__32093\
        );

    \I__5825\ : Span4Mux_v
    port map (
            O => \N__32096\,
            I => \N__32088\
        );

    \I__5824\ : Span4Mux_h
    port map (
            O => \N__32093\,
            I => \N__32085\
        );

    \I__5823\ : InMux
    port map (
            O => \N__32092\,
            I => \N__32080\
        );

    \I__5822\ : InMux
    port map (
            O => \N__32091\,
            I => \N__32080\
        );

    \I__5821\ : Odrv4
    port map (
            O => \N__32088\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__5820\ : Odrv4
    port map (
            O => \N__32085\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__32080\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__5818\ : InMux
    port map (
            O => \N__32073\,
            I => \N__32070\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__32070\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_5\
        );

    \I__5816\ : CascadeMux
    port map (
            O => \N__32067\,
            I => \N__32064\
        );

    \I__5815\ : InMux
    port map (
            O => \N__32064\,
            I => \N__32061\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__32061\,
            I => \N__32058\
        );

    \I__5813\ : Span4Mux_h
    port map (
            O => \N__32058\,
            I => \N__32055\
        );

    \I__5812\ : Odrv4
    port map (
            O => \N__32055\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI5R3UZ0Z_5\
        );

    \I__5811\ : InMux
    port map (
            O => \N__32052\,
            I => \N__32049\
        );

    \I__5810\ : LocalMux
    port map (
            O => \N__32049\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\
        );

    \I__5809\ : InMux
    port map (
            O => \N__32046\,
            I => \N__32043\
        );

    \I__5808\ : LocalMux
    port map (
            O => \N__32043\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\
        );

    \I__5807\ : InMux
    port map (
            O => \N__32040\,
            I => \N__32037\
        );

    \I__5806\ : LocalMux
    port map (
            O => \N__32037\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\
        );

    \I__5805\ : InMux
    port map (
            O => \N__32034\,
            I => \N__32031\
        );

    \I__5804\ : LocalMux
    port map (
            O => \N__32031\,
            I => \N__32028\
        );

    \I__5803\ : Glb2LocalMux
    port map (
            O => \N__32028\,
            I => \N__32025\
        );

    \I__5802\ : GlobalMux
    port map (
            O => \N__32025\,
            I => clk_12mhz
        );

    \I__5801\ : IoInMux
    port map (
            O => \N__32022\,
            I => \N__32019\
        );

    \I__5800\ : LocalMux
    port map (
            O => \N__32019\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__5799\ : IoInMux
    port map (
            O => \N__32016\,
            I => \N__32013\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__32013\,
            I => \N__32010\
        );

    \I__5797\ : Span4Mux_s1_v
    port map (
            O => \N__32010\,
            I => \N__32007\
        );

    \I__5796\ : Odrv4
    port map (
            O => \N__32007\,
            I => \delay_measurement_inst.delay_tr_timer.N_395_i\
        );

    \I__5795\ : ClkMux
    port map (
            O => \N__32004\,
            I => \N__32001\
        );

    \I__5794\ : GlobalMux
    port map (
            O => \N__32001\,
            I => \N__31998\
        );

    \I__5793\ : gio2CtrlBuf
    port map (
            O => \N__31998\,
            I => delay_tr_input_c_g
        );

    \I__5792\ : InMux
    port map (
            O => \N__31995\,
            I => \N__31991\
        );

    \I__5791\ : InMux
    port map (
            O => \N__31994\,
            I => \N__31988\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__31991\,
            I => \N__31982\
        );

    \I__5789\ : LocalMux
    port map (
            O => \N__31988\,
            I => \N__31982\
        );

    \I__5788\ : InMux
    port map (
            O => \N__31987\,
            I => \N__31979\
        );

    \I__5787\ : Span4Mux_v
    port map (
            O => \N__31982\,
            I => \N__31976\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__31979\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\
        );

    \I__5785\ : Odrv4
    port map (
            O => \N__31976\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\
        );

    \I__5784\ : InMux
    port map (
            O => \N__31971\,
            I => \N__31965\
        );

    \I__5783\ : InMux
    port map (
            O => \N__31970\,
            I => \N__31962\
        );

    \I__5782\ : InMux
    port map (
            O => \N__31969\,
            I => \N__31958\
        );

    \I__5781\ : InMux
    port map (
            O => \N__31968\,
            I => \N__31955\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__31965\,
            I => \N__31952\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__31962\,
            I => \N__31949\
        );

    \I__5778\ : InMux
    port map (
            O => \N__31961\,
            I => \N__31946\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__31958\,
            I => \N__31941\
        );

    \I__5776\ : LocalMux
    port map (
            O => \N__31955\,
            I => \N__31941\
        );

    \I__5775\ : Span4Mux_h
    port map (
            O => \N__31952\,
            I => \N__31936\
        );

    \I__5774\ : Span4Mux_v
    port map (
            O => \N__31949\,
            I => \N__31936\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__31946\,
            I => \N__31933\
        );

    \I__5772\ : Span4Mux_h
    port map (
            O => \N__31941\,
            I => \N__31930\
        );

    \I__5771\ : Odrv4
    port map (
            O => \N__31936\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__5770\ : Odrv12
    port map (
            O => \N__31933\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__5769\ : Odrv4
    port map (
            O => \N__31930\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__5768\ : InMux
    port map (
            O => \N__31923\,
            I => \N__31920\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__31920\,
            I => \N__31917\
        );

    \I__5766\ : Span4Mux_v
    port map (
            O => \N__31917\,
            I => \N__31914\
        );

    \I__5765\ : Span4Mux_h
    port map (
            O => \N__31914\,
            I => \N__31911\
        );

    \I__5764\ : Odrv4
    port map (
            O => \N__31911\,
            I => \current_shift_inst.PI_CTRL.integrator_i_27\
        );

    \I__5763\ : InMux
    port map (
            O => \N__31908\,
            I => \N__31904\
        );

    \I__5762\ : CascadeMux
    port map (
            O => \N__31907\,
            I => \N__31901\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__31904\,
            I => \N__31896\
        );

    \I__5760\ : InMux
    port map (
            O => \N__31901\,
            I => \N__31893\
        );

    \I__5759\ : InMux
    port map (
            O => \N__31900\,
            I => \N__31890\
        );

    \I__5758\ : InMux
    port map (
            O => \N__31899\,
            I => \N__31887\
        );

    \I__5757\ : Span4Mux_v
    port map (
            O => \N__31896\,
            I => \N__31881\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__31893\,
            I => \N__31881\
        );

    \I__5755\ : LocalMux
    port map (
            O => \N__31890\,
            I => \N__31878\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__31887\,
            I => \N__31875\
        );

    \I__5753\ : InMux
    port map (
            O => \N__31886\,
            I => \N__31872\
        );

    \I__5752\ : Span4Mux_h
    port map (
            O => \N__31881\,
            I => \N__31867\
        );

    \I__5751\ : Span4Mux_h
    port map (
            O => \N__31878\,
            I => \N__31867\
        );

    \I__5750\ : Odrv4
    port map (
            O => \N__31875\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__31872\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__5748\ : Odrv4
    port map (
            O => \N__31867\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__5747\ : InMux
    port map (
            O => \N__31860\,
            I => \N__31857\
        );

    \I__5746\ : LocalMux
    port map (
            O => \N__31857\,
            I => \N__31854\
        );

    \I__5745\ : Span4Mux_h
    port map (
            O => \N__31854\,
            I => \N__31851\
        );

    \I__5744\ : Odrv4
    port map (
            O => \N__31851\,
            I => \current_shift_inst.PI_CTRL.integrator_i_13\
        );

    \I__5743\ : CascadeMux
    port map (
            O => \N__31848\,
            I => \N__31844\
        );

    \I__5742\ : InMux
    port map (
            O => \N__31847\,
            I => \N__31840\
        );

    \I__5741\ : InMux
    port map (
            O => \N__31844\,
            I => \N__31837\
        );

    \I__5740\ : InMux
    port map (
            O => \N__31843\,
            I => \N__31832\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__31840\,
            I => \N__31829\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__31837\,
            I => \N__31826\
        );

    \I__5737\ : InMux
    port map (
            O => \N__31836\,
            I => \N__31821\
        );

    \I__5736\ : InMux
    port map (
            O => \N__31835\,
            I => \N__31821\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__31832\,
            I => \N__31818\
        );

    \I__5734\ : Span12Mux_h
    port map (
            O => \N__31829\,
            I => \N__31813\
        );

    \I__5733\ : Span12Mux_s8_h
    port map (
            O => \N__31826\,
            I => \N__31813\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__31821\,
            I => \N__31810\
        );

    \I__5731\ : Span4Mux_h
    port map (
            O => \N__31818\,
            I => \N__31807\
        );

    \I__5730\ : Odrv12
    port map (
            O => \N__31813\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__5729\ : Odrv12
    port map (
            O => \N__31810\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__5728\ : Odrv4
    port map (
            O => \N__31807\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__5727\ : InMux
    port map (
            O => \N__31800\,
            I => \N__31797\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__31797\,
            I => \N__31794\
        );

    \I__5725\ : Span4Mux_v
    port map (
            O => \N__31794\,
            I => \N__31791\
        );

    \I__5724\ : Odrv4
    port map (
            O => \N__31791\,
            I => \current_shift_inst.PI_CTRL.integrator_i_22\
        );

    \I__5723\ : InMux
    port map (
            O => \N__31788\,
            I => \N__31785\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__31785\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\
        );

    \I__5721\ : CascadeMux
    port map (
            O => \N__31782\,
            I => \N__31779\
        );

    \I__5720\ : InMux
    port map (
            O => \N__31779\,
            I => \N__31776\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__31776\,
            I => \N__31773\
        );

    \I__5718\ : Span4Mux_h
    port map (
            O => \N__31773\,
            I => \N__31769\
        );

    \I__5717\ : InMux
    port map (
            O => \N__31772\,
            I => \N__31766\
        );

    \I__5716\ : Odrv4
    port map (
            O => \N__31769\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__31766\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__5714\ : CascadeMux
    port map (
            O => \N__31761\,
            I => \N__31757\
        );

    \I__5713\ : InMux
    port map (
            O => \N__31760\,
            I => \N__31752\
        );

    \I__5712\ : InMux
    port map (
            O => \N__31757\,
            I => \N__31752\
        );

    \I__5711\ : LocalMux
    port map (
            O => \N__31752\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__5710\ : CascadeMux
    port map (
            O => \N__31749\,
            I => \N__31746\
        );

    \I__5709\ : InMux
    port map (
            O => \N__31746\,
            I => \N__31743\
        );

    \I__5708\ : LocalMux
    port map (
            O => \N__31743\,
            I => \N__31739\
        );

    \I__5707\ : InMux
    port map (
            O => \N__31742\,
            I => \N__31736\
        );

    \I__5706\ : Odrv12
    port map (
            O => \N__31739\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__31736\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__5704\ : InMux
    port map (
            O => \N__31731\,
            I => \N__31728\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__31728\,
            I => \N__31725\
        );

    \I__5702\ : Odrv12
    port map (
            O => \N__31725\,
            I => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_19\
        );

    \I__5701\ : CascadeMux
    port map (
            O => \N__31722\,
            I => \N__31719\
        );

    \I__5700\ : InMux
    port map (
            O => \N__31719\,
            I => \N__31714\
        );

    \I__5699\ : InMux
    port map (
            O => \N__31718\,
            I => \N__31711\
        );

    \I__5698\ : InMux
    port map (
            O => \N__31717\,
            I => \N__31708\
        );

    \I__5697\ : LocalMux
    port map (
            O => \N__31714\,
            I => \N__31701\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__31711\,
            I => \N__31701\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__31708\,
            I => \N__31698\
        );

    \I__5694\ : InMux
    port map (
            O => \N__31707\,
            I => \N__31693\
        );

    \I__5693\ : InMux
    port map (
            O => \N__31706\,
            I => \N__31693\
        );

    \I__5692\ : Span4Mux_v
    port map (
            O => \N__31701\,
            I => \N__31686\
        );

    \I__5691\ : Span4Mux_h
    port map (
            O => \N__31698\,
            I => \N__31686\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__31693\,
            I => \N__31686\
        );

    \I__5689\ : Odrv4
    port map (
            O => \N__31686\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__5688\ : InMux
    port map (
            O => \N__31683\,
            I => \N__31679\
        );

    \I__5687\ : InMux
    port map (
            O => \N__31682\,
            I => \N__31676\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__31679\,
            I => \N__31673\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__31676\,
            I => \N__31670\
        );

    \I__5684\ : Span12Mux_v
    port map (
            O => \N__31673\,
            I => \N__31667\
        );

    \I__5683\ : Odrv12
    port map (
            O => \N__31670\,
            I => state_ns_i_a2_1
        );

    \I__5682\ : Odrv12
    port map (
            O => \N__31667\,
            I => state_ns_i_a2_1
        );

    \I__5681\ : InMux
    port map (
            O => \N__31662\,
            I => \N__31659\
        );

    \I__5680\ : LocalMux
    port map (
            O => \N__31659\,
            I => \phase_controller_inst1.start_timer_hc_RNOZ0Z_0\
        );

    \I__5679\ : InMux
    port map (
            O => \N__31656\,
            I => \N__31653\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__31653\,
            I => \phase_controller_inst1.start_timer_hc_0_sqmuxa\
        );

    \I__5677\ : CascadeMux
    port map (
            O => \N__31650\,
            I => \N__31645\
        );

    \I__5676\ : InMux
    port map (
            O => \N__31649\,
            I => \N__31641\
        );

    \I__5675\ : InMux
    port map (
            O => \N__31648\,
            I => \N__31638\
        );

    \I__5674\ : InMux
    port map (
            O => \N__31645\,
            I => \N__31633\
        );

    \I__5673\ : InMux
    port map (
            O => \N__31644\,
            I => \N__31633\
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__31641\,
            I => \N__31630\
        );

    \I__5671\ : LocalMux
    port map (
            O => \N__31638\,
            I => \N__31627\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__31633\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__5669\ : Odrv12
    port map (
            O => \N__31630\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__5668\ : Odrv4
    port map (
            O => \N__31627\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__5667\ : CascadeMux
    port map (
            O => \N__31620\,
            I => \N__31617\
        );

    \I__5666\ : InMux
    port map (
            O => \N__31617\,
            I => \N__31614\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__31614\,
            I => \N__31609\
        );

    \I__5664\ : InMux
    port map (
            O => \N__31613\,
            I => \N__31606\
        );

    \I__5663\ : InMux
    port map (
            O => \N__31612\,
            I => \N__31603\
        );

    \I__5662\ : Span4Mux_v
    port map (
            O => \N__31609\,
            I => \N__31600\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__31606\,
            I => \N__31597\
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__31603\,
            I => \N__31594\
        );

    \I__5659\ : Span4Mux_h
    port map (
            O => \N__31600\,
            I => \N__31589\
        );

    \I__5658\ : Span4Mux_h
    port map (
            O => \N__31597\,
            I => \N__31589\
        );

    \I__5657\ : Span12Mux_h
    port map (
            O => \N__31594\,
            I => \N__31584\
        );

    \I__5656\ : Sp12to4
    port map (
            O => \N__31589\,
            I => \N__31584\
        );

    \I__5655\ : Span12Mux_v
    port map (
            O => \N__31584\,
            I => \N__31581\
        );

    \I__5654\ : Odrv12
    port map (
            O => \N__31581\,
            I => \il_max_comp1_D2\
        );

    \I__5653\ : CascadeMux
    port map (
            O => \N__31578\,
            I => \N__31574\
        );

    \I__5652\ : InMux
    port map (
            O => \N__31577\,
            I => \N__31571\
        );

    \I__5651\ : InMux
    port map (
            O => \N__31574\,
            I => \N__31568\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__31571\,
            I => \N__31562\
        );

    \I__5649\ : LocalMux
    port map (
            O => \N__31568\,
            I => \N__31562\
        );

    \I__5648\ : InMux
    port map (
            O => \N__31567\,
            I => \N__31559\
        );

    \I__5647\ : Span4Mux_v
    port map (
            O => \N__31562\,
            I => \N__31553\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__31559\,
            I => \N__31553\
        );

    \I__5645\ : InMux
    port map (
            O => \N__31558\,
            I => \N__31550\
        );

    \I__5644\ : Span4Mux_h
    port map (
            O => \N__31553\,
            I => \N__31547\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__31550\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__5642\ : Odrv4
    port map (
            O => \N__31547\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__5641\ : CascadeMux
    port map (
            O => \N__31542\,
            I => \N__31538\
        );

    \I__5640\ : InMux
    port map (
            O => \N__31541\,
            I => \N__31534\
        );

    \I__5639\ : InMux
    port map (
            O => \N__31538\,
            I => \N__31531\
        );

    \I__5638\ : InMux
    port map (
            O => \N__31537\,
            I => \N__31528\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__31534\,
            I => \N__31525\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__31531\,
            I => \N__31521\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__31528\,
            I => \N__31516\
        );

    \I__5634\ : Span4Mux_v
    port map (
            O => \N__31525\,
            I => \N__31516\
        );

    \I__5633\ : InMux
    port map (
            O => \N__31524\,
            I => \N__31513\
        );

    \I__5632\ : Odrv4
    port map (
            O => \N__31521\,
            I => \elapsed_time_ns_1_RNI5GT8E1_0_13\
        );

    \I__5631\ : Odrv4
    port map (
            O => \N__31516\,
            I => \elapsed_time_ns_1_RNI5GT8E1_0_13\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__31513\,
            I => \elapsed_time_ns_1_RNI5GT8E1_0_13\
        );

    \I__5629\ : CascadeMux
    port map (
            O => \N__31506\,
            I => \N__31499\
        );

    \I__5628\ : CascadeMux
    port map (
            O => \N__31505\,
            I => \N__31496\
        );

    \I__5627\ : CascadeMux
    port map (
            O => \N__31504\,
            I => \N__31490\
        );

    \I__5626\ : InMux
    port map (
            O => \N__31503\,
            I => \N__31480\
        );

    \I__5625\ : InMux
    port map (
            O => \N__31502\,
            I => \N__31480\
        );

    \I__5624\ : InMux
    port map (
            O => \N__31499\,
            I => \N__31480\
        );

    \I__5623\ : InMux
    port map (
            O => \N__31496\,
            I => \N__31480\
        );

    \I__5622\ : InMux
    port map (
            O => \N__31495\,
            I => \N__31470\
        );

    \I__5621\ : InMux
    port map (
            O => \N__31494\,
            I => \N__31470\
        );

    \I__5620\ : InMux
    port map (
            O => \N__31493\,
            I => \N__31470\
        );

    \I__5619\ : InMux
    port map (
            O => \N__31490\,
            I => \N__31470\
        );

    \I__5618\ : InMux
    port map (
            O => \N__31489\,
            I => \N__31467\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__31480\,
            I => \N__31464\
        );

    \I__5616\ : InMux
    port map (
            O => \N__31479\,
            I => \N__31461\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__31470\,
            I => \N__31456\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__31467\,
            I => \N__31456\
        );

    \I__5613\ : Span4Mux_v
    port map (
            O => \N__31464\,
            I => \N__31453\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__31461\,
            I => \N__31448\
        );

    \I__5611\ : Span4Mux_v
    port map (
            O => \N__31456\,
            I => \N__31448\
        );

    \I__5610\ : Odrv4
    port map (
            O => \N__31453\,
            I => \phase_controller_inst1.stoper_hc.N_316\
        );

    \I__5609\ : Odrv4
    port map (
            O => \N__31448\,
            I => \phase_controller_inst1.stoper_hc.N_316\
        );

    \I__5608\ : CascadeMux
    port map (
            O => \N__31443\,
            I => \N__31434\
        );

    \I__5607\ : CascadeMux
    port map (
            O => \N__31442\,
            I => \N__31426\
        );

    \I__5606\ : CascadeMux
    port map (
            O => \N__31441\,
            I => \N__31422\
        );

    \I__5605\ : CascadeMux
    port map (
            O => \N__31440\,
            I => \N__31419\
        );

    \I__5604\ : InMux
    port map (
            O => \N__31439\,
            I => \N__31410\
        );

    \I__5603\ : InMux
    port map (
            O => \N__31438\,
            I => \N__31410\
        );

    \I__5602\ : InMux
    port map (
            O => \N__31437\,
            I => \N__31410\
        );

    \I__5601\ : InMux
    port map (
            O => \N__31434\,
            I => \N__31410\
        );

    \I__5600\ : InMux
    port map (
            O => \N__31433\,
            I => \N__31401\
        );

    \I__5599\ : InMux
    port map (
            O => \N__31432\,
            I => \N__31401\
        );

    \I__5598\ : InMux
    port map (
            O => \N__31431\,
            I => \N__31401\
        );

    \I__5597\ : InMux
    port map (
            O => \N__31430\,
            I => \N__31401\
        );

    \I__5596\ : InMux
    port map (
            O => \N__31429\,
            I => \N__31392\
        );

    \I__5595\ : InMux
    port map (
            O => \N__31426\,
            I => \N__31389\
        );

    \I__5594\ : InMux
    port map (
            O => \N__31425\,
            I => \N__31382\
        );

    \I__5593\ : InMux
    port map (
            O => \N__31422\,
            I => \N__31382\
        );

    \I__5592\ : InMux
    port map (
            O => \N__31419\,
            I => \N__31382\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__31410\,
            I => \N__31377\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__31401\,
            I => \N__31377\
        );

    \I__5589\ : CascadeMux
    port map (
            O => \N__31400\,
            I => \N__31373\
        );

    \I__5588\ : InMux
    port map (
            O => \N__31399\,
            I => \N__31359\
        );

    \I__5587\ : InMux
    port map (
            O => \N__31398\,
            I => \N__31359\
        );

    \I__5586\ : InMux
    port map (
            O => \N__31397\,
            I => \N__31359\
        );

    \I__5585\ : InMux
    port map (
            O => \N__31396\,
            I => \N__31359\
        );

    \I__5584\ : InMux
    port map (
            O => \N__31395\,
            I => \N__31359\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__31392\,
            I => \N__31350\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__31389\,
            I => \N__31350\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__31382\,
            I => \N__31350\
        );

    \I__5580\ : Span4Mux_v
    port map (
            O => \N__31377\,
            I => \N__31350\
        );

    \I__5579\ : InMux
    port map (
            O => \N__31376\,
            I => \N__31347\
        );

    \I__5578\ : InMux
    port map (
            O => \N__31373\,
            I => \N__31341\
        );

    \I__5577\ : InMux
    port map (
            O => \N__31372\,
            I => \N__31334\
        );

    \I__5576\ : InMux
    port map (
            O => \N__31371\,
            I => \N__31334\
        );

    \I__5575\ : InMux
    port map (
            O => \N__31370\,
            I => \N__31334\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__31359\,
            I => \N__31331\
        );

    \I__5573\ : Span4Mux_v
    port map (
            O => \N__31350\,
            I => \N__31326\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__31347\,
            I => \N__31326\
        );

    \I__5571\ : InMux
    port map (
            O => \N__31346\,
            I => \N__31323\
        );

    \I__5570\ : InMux
    port map (
            O => \N__31345\,
            I => \N__31318\
        );

    \I__5569\ : InMux
    port map (
            O => \N__31344\,
            I => \N__31318\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__31341\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__31334\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\
        );

    \I__5566\ : Odrv4
    port map (
            O => \N__31331\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\
        );

    \I__5565\ : Odrv4
    port map (
            O => \N__31326\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\
        );

    \I__5564\ : LocalMux
    port map (
            O => \N__31323\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__31318\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\
        );

    \I__5562\ : InMux
    port map (
            O => \N__31305\,
            I => \N__31301\
        );

    \I__5561\ : InMux
    port map (
            O => \N__31304\,
            I => \N__31298\
        );

    \I__5560\ : LocalMux
    port map (
            O => \N__31301\,
            I => \N__31295\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__31298\,
            I => \N__31292\
        );

    \I__5558\ : Span4Mux_v
    port map (
            O => \N__31295\,
            I => \N__31287\
        );

    \I__5557\ : Span4Mux_h
    port map (
            O => \N__31292\,
            I => \N__31284\
        );

    \I__5556\ : InMux
    port map (
            O => \N__31291\,
            I => \N__31279\
        );

    \I__5555\ : InMux
    port map (
            O => \N__31290\,
            I => \N__31279\
        );

    \I__5554\ : Odrv4
    port map (
            O => \N__31287\,
            I => \elapsed_time_ns_1_RNIHHC6P1_0_18\
        );

    \I__5553\ : Odrv4
    port map (
            O => \N__31284\,
            I => \elapsed_time_ns_1_RNIHHC6P1_0_18\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__31279\,
            I => \elapsed_time_ns_1_RNIHHC6P1_0_18\
        );

    \I__5551\ : InMux
    port map (
            O => \N__31272\,
            I => \N__31269\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__31269\,
            I => \N__31265\
        );

    \I__5549\ : InMux
    port map (
            O => \N__31268\,
            I => \N__31262\
        );

    \I__5548\ : Span4Mux_h
    port map (
            O => \N__31265\,
            I => \N__31259\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__31262\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\
        );

    \I__5546\ : Odrv4
    port map (
            O => \N__31259\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\
        );

    \I__5545\ : InMux
    port map (
            O => \N__31254\,
            I => \N__31251\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__31251\,
            I => \N__31248\
        );

    \I__5543\ : Span4Mux_v
    port map (
            O => \N__31248\,
            I => \N__31244\
        );

    \I__5542\ : InMux
    port map (
            O => \N__31247\,
            I => \N__31241\
        );

    \I__5541\ : Odrv4
    port map (
            O => \N__31244\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__31241\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\
        );

    \I__5539\ : InMux
    port map (
            O => \N__31236\,
            I => \N__31232\
        );

    \I__5538\ : InMux
    port map (
            O => \N__31235\,
            I => \N__31227\
        );

    \I__5537\ : LocalMux
    port map (
            O => \N__31232\,
            I => \N__31224\
        );

    \I__5536\ : InMux
    port map (
            O => \N__31231\,
            I => \N__31221\
        );

    \I__5535\ : InMux
    port map (
            O => \N__31230\,
            I => \N__31218\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__31227\,
            I => \N__31213\
        );

    \I__5533\ : Span4Mux_v
    port map (
            O => \N__31224\,
            I => \N__31213\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__31221\,
            I => \N__31210\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__31218\,
            I => \elapsed_time_ns_1_RNIPKKEE1_0_8\
        );

    \I__5530\ : Odrv4
    port map (
            O => \N__31213\,
            I => \elapsed_time_ns_1_RNIPKKEE1_0_8\
        );

    \I__5529\ : Odrv12
    port map (
            O => \N__31210\,
            I => \elapsed_time_ns_1_RNIPKKEE1_0_8\
        );

    \I__5528\ : InMux
    port map (
            O => \N__31203\,
            I => \N__31200\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__31200\,
            I => \N__31196\
        );

    \I__5526\ : InMux
    port map (
            O => \N__31199\,
            I => \N__31193\
        );

    \I__5525\ : Odrv4
    port map (
            O => \N__31196\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__31193\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__5523\ : InMux
    port map (
            O => \N__31188\,
            I => \N__31185\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__31185\,
            I => \N__31181\
        );

    \I__5521\ : InMux
    port map (
            O => \N__31184\,
            I => \N__31178\
        );

    \I__5520\ : Odrv4
    port map (
            O => \N__31181\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__31178\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__5518\ : InMux
    port map (
            O => \N__31173\,
            I => \N__31169\
        );

    \I__5517\ : CascadeMux
    port map (
            O => \N__31172\,
            I => \N__31166\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__31169\,
            I => \N__31163\
        );

    \I__5515\ : InMux
    port map (
            O => \N__31166\,
            I => \N__31160\
        );

    \I__5514\ : Odrv4
    port map (
            O => \N__31163\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__31160\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__5512\ : InMux
    port map (
            O => \N__31155\,
            I => \N__31152\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__31152\,
            I => \N__31148\
        );

    \I__5510\ : InMux
    port map (
            O => \N__31151\,
            I => \N__31145\
        );

    \I__5509\ : Odrv4
    port map (
            O => \N__31148\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__31145\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__5507\ : InMux
    port map (
            O => \N__31140\,
            I => \N__31137\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__31137\,
            I => \N__31134\
        );

    \I__5505\ : Sp12to4
    port map (
            O => \N__31134\,
            I => \N__31131\
        );

    \I__5504\ : Odrv12
    port map (
            O => \N__31131\,
            I => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_17\
        );

    \I__5503\ : InMux
    port map (
            O => \N__31128\,
            I => \N__31125\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__31125\,
            I => \N__31119\
        );

    \I__5501\ : InMux
    port map (
            O => \N__31124\,
            I => \N__31116\
        );

    \I__5500\ : InMux
    port map (
            O => \N__31123\,
            I => \N__31113\
        );

    \I__5499\ : CascadeMux
    port map (
            O => \N__31122\,
            I => \N__31100\
        );

    \I__5498\ : Span4Mux_v
    port map (
            O => \N__31119\,
            I => \N__31094\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__31116\,
            I => \N__31094\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__31113\,
            I => \N__31089\
        );

    \I__5495\ : InMux
    port map (
            O => \N__31112\,
            I => \N__31086\
        );

    \I__5494\ : CascadeMux
    port map (
            O => \N__31111\,
            I => \N__31082\
        );

    \I__5493\ : CascadeMux
    port map (
            O => \N__31110\,
            I => \N__31077\
        );

    \I__5492\ : CascadeMux
    port map (
            O => \N__31109\,
            I => \N__31074\
        );

    \I__5491\ : CascadeMux
    port map (
            O => \N__31108\,
            I => \N__31069\
        );

    \I__5490\ : CascadeMux
    port map (
            O => \N__31107\,
            I => \N__31063\
        );

    \I__5489\ : InMux
    port map (
            O => \N__31106\,
            I => \N__31058\
        );

    \I__5488\ : InMux
    port map (
            O => \N__31105\,
            I => \N__31058\
        );

    \I__5487\ : CascadeMux
    port map (
            O => \N__31104\,
            I => \N__31052\
        );

    \I__5486\ : InMux
    port map (
            O => \N__31103\,
            I => \N__31049\
        );

    \I__5485\ : InMux
    port map (
            O => \N__31100\,
            I => \N__31044\
        );

    \I__5484\ : InMux
    port map (
            O => \N__31099\,
            I => \N__31044\
        );

    \I__5483\ : Span4Mux_v
    port map (
            O => \N__31094\,
            I => \N__31039\
        );

    \I__5482\ : InMux
    port map (
            O => \N__31093\,
            I => \N__31036\
        );

    \I__5481\ : InMux
    port map (
            O => \N__31092\,
            I => \N__31033\
        );

    \I__5480\ : Span12Mux_h
    port map (
            O => \N__31089\,
            I => \N__31028\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__31086\,
            I => \N__31028\
        );

    \I__5478\ : InMux
    port map (
            O => \N__31085\,
            I => \N__31019\
        );

    \I__5477\ : InMux
    port map (
            O => \N__31082\,
            I => \N__31019\
        );

    \I__5476\ : InMux
    port map (
            O => \N__31081\,
            I => \N__31019\
        );

    \I__5475\ : InMux
    port map (
            O => \N__31080\,
            I => \N__31019\
        );

    \I__5474\ : InMux
    port map (
            O => \N__31077\,
            I => \N__31010\
        );

    \I__5473\ : InMux
    port map (
            O => \N__31074\,
            I => \N__31010\
        );

    \I__5472\ : InMux
    port map (
            O => \N__31073\,
            I => \N__31010\
        );

    \I__5471\ : InMux
    port map (
            O => \N__31072\,
            I => \N__31010\
        );

    \I__5470\ : InMux
    port map (
            O => \N__31069\,
            I => \N__30999\
        );

    \I__5469\ : InMux
    port map (
            O => \N__31068\,
            I => \N__30999\
        );

    \I__5468\ : InMux
    port map (
            O => \N__31067\,
            I => \N__30999\
        );

    \I__5467\ : InMux
    port map (
            O => \N__31066\,
            I => \N__30999\
        );

    \I__5466\ : InMux
    port map (
            O => \N__31063\,
            I => \N__30999\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__31058\,
            I => \N__30996\
        );

    \I__5464\ : InMux
    port map (
            O => \N__31057\,
            I => \N__30987\
        );

    \I__5463\ : InMux
    port map (
            O => \N__31056\,
            I => \N__30987\
        );

    \I__5462\ : InMux
    port map (
            O => \N__31055\,
            I => \N__30987\
        );

    \I__5461\ : InMux
    port map (
            O => \N__31052\,
            I => \N__30987\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__31049\,
            I => \N__30982\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__31044\,
            I => \N__30982\
        );

    \I__5458\ : InMux
    port map (
            O => \N__31043\,
            I => \N__30977\
        );

    \I__5457\ : InMux
    port map (
            O => \N__31042\,
            I => \N__30977\
        );

    \I__5456\ : Odrv4
    port map (
            O => \N__31039\,
            I => \delay_measurement_inst.delay_hc_timer.N_365_clk\
        );

    \I__5455\ : LocalMux
    port map (
            O => \N__31036\,
            I => \delay_measurement_inst.delay_hc_timer.N_365_clk\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__31033\,
            I => \delay_measurement_inst.delay_hc_timer.N_365_clk\
        );

    \I__5453\ : Odrv12
    port map (
            O => \N__31028\,
            I => \delay_measurement_inst.delay_hc_timer.N_365_clk\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__31019\,
            I => \delay_measurement_inst.delay_hc_timer.N_365_clk\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__31010\,
            I => \delay_measurement_inst.delay_hc_timer.N_365_clk\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__30999\,
            I => \delay_measurement_inst.delay_hc_timer.N_365_clk\
        );

    \I__5449\ : Odrv4
    port map (
            O => \N__30996\,
            I => \delay_measurement_inst.delay_hc_timer.N_365_clk\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__30987\,
            I => \delay_measurement_inst.delay_hc_timer.N_365_clk\
        );

    \I__5447\ : Odrv4
    port map (
            O => \N__30982\,
            I => \delay_measurement_inst.delay_hc_timer.N_365_clk\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__30977\,
            I => \delay_measurement_inst.delay_hc_timer.N_365_clk\
        );

    \I__5445\ : CascadeMux
    port map (
            O => \N__30954\,
            I => \N__30951\
        );

    \I__5444\ : InMux
    port map (
            O => \N__30951\,
            I => \N__30946\
        );

    \I__5443\ : InMux
    port map (
            O => \N__30950\,
            I => \N__30942\
        );

    \I__5442\ : CascadeMux
    port map (
            O => \N__30949\,
            I => \N__30939\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__30946\,
            I => \N__30935\
        );

    \I__5440\ : InMux
    port map (
            O => \N__30945\,
            I => \N__30932\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__30942\,
            I => \N__30929\
        );

    \I__5438\ : InMux
    port map (
            O => \N__30939\,
            I => \N__30924\
        );

    \I__5437\ : InMux
    port map (
            O => \N__30938\,
            I => \N__30924\
        );

    \I__5436\ : Odrv4
    port map (
            O => \N__30935\,
            I => \elapsed_time_ns_1_RNIIIC6P1_0_19\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__30932\,
            I => \elapsed_time_ns_1_RNIIIC6P1_0_19\
        );

    \I__5434\ : Odrv12
    port map (
            O => \N__30929\,
            I => \elapsed_time_ns_1_RNIIIC6P1_0_19\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__30924\,
            I => \elapsed_time_ns_1_RNIIIC6P1_0_19\
        );

    \I__5432\ : InMux
    port map (
            O => \N__30915\,
            I => \N__30912\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__30912\,
            I => \N__30909\
        );

    \I__5430\ : Odrv4
    port map (
            O => \N__30909\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19\
        );

    \I__5429\ : InMux
    port map (
            O => \N__30906\,
            I => \N__30903\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__30903\,
            I => \N__30900\
        );

    \I__5427\ : Span4Mux_v
    port map (
            O => \N__30900\,
            I => \N__30896\
        );

    \I__5426\ : InMux
    port map (
            O => \N__30899\,
            I => \N__30893\
        );

    \I__5425\ : Odrv4
    port map (
            O => \N__30896\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__30893\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__5423\ : CascadeMux
    port map (
            O => \N__30888\,
            I => \N__30885\
        );

    \I__5422\ : InMux
    port map (
            O => \N__30885\,
            I => \N__30882\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__30882\,
            I => \N__30878\
        );

    \I__5420\ : InMux
    port map (
            O => \N__30881\,
            I => \N__30875\
        );

    \I__5419\ : Odrv12
    port map (
            O => \N__30878\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__30875\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__5417\ : InMux
    port map (
            O => \N__30870\,
            I => \N__30866\
        );

    \I__5416\ : CascadeMux
    port map (
            O => \N__30869\,
            I => \N__30863\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__30866\,
            I => \N__30860\
        );

    \I__5414\ : InMux
    port map (
            O => \N__30863\,
            I => \N__30857\
        );

    \I__5413\ : Odrv12
    port map (
            O => \N__30860\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__30857\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__5411\ : InMux
    port map (
            O => \N__30852\,
            I => \N__30849\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__30849\,
            I => \N__30846\
        );

    \I__5409\ : Span4Mux_v
    port map (
            O => \N__30846\,
            I => \N__30842\
        );

    \I__5408\ : InMux
    port map (
            O => \N__30845\,
            I => \N__30839\
        );

    \I__5407\ : Odrv4
    port map (
            O => \N__30842\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__30839\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__5405\ : InMux
    port map (
            O => \N__30834\,
            I => \N__30831\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__30831\,
            I => \N__30828\
        );

    \I__5403\ : Odrv4
    port map (
            O => \N__30828\,
            I => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_18\
        );

    \I__5402\ : InMux
    port map (
            O => \N__30825\,
            I => \N__30822\
        );

    \I__5401\ : LocalMux
    port map (
            O => \N__30822\,
            I => \N__30818\
        );

    \I__5400\ : InMux
    port map (
            O => \N__30821\,
            I => \N__30815\
        );

    \I__5399\ : Odrv12
    port map (
            O => \N__30818\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__30815\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__5397\ : CascadeMux
    port map (
            O => \N__30810\,
            I => \N__30807\
        );

    \I__5396\ : InMux
    port map (
            O => \N__30807\,
            I => \N__30803\
        );

    \I__5395\ : InMux
    port map (
            O => \N__30806\,
            I => \N__30800\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__30803\,
            I => \N__30797\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__30800\,
            I => \N__30794\
        );

    \I__5392\ : Span4Mux_v
    port map (
            O => \N__30797\,
            I => \N__30791\
        );

    \I__5391\ : Odrv4
    port map (
            O => \N__30794\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__5390\ : Odrv4
    port map (
            O => \N__30791\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__5389\ : InMux
    port map (
            O => \N__30786\,
            I => \N__30782\
        );

    \I__5388\ : InMux
    port map (
            O => \N__30785\,
            I => \N__30779\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__30782\,
            I => \N__30776\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__30779\,
            I => \N__30773\
        );

    \I__5385\ : Span12Mux_v
    port map (
            O => \N__30776\,
            I => \N__30770\
        );

    \I__5384\ : Span4Mux_h
    port map (
            O => \N__30773\,
            I => \N__30767\
        );

    \I__5383\ : Odrv12
    port map (
            O => \N__30770\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__5382\ : Odrv4
    port map (
            O => \N__30767\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__5381\ : InMux
    port map (
            O => \N__30762\,
            I => \N__30759\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__30759\,
            I => \N__30755\
        );

    \I__5379\ : InMux
    port map (
            O => \N__30758\,
            I => \N__30752\
        );

    \I__5378\ : Span4Mux_h
    port map (
            O => \N__30755\,
            I => \N__30747\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__30752\,
            I => \N__30747\
        );

    \I__5376\ : Odrv4
    port map (
            O => \N__30747\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__5375\ : CascadeMux
    port map (
            O => \N__30744\,
            I => \N__30740\
        );

    \I__5374\ : InMux
    port map (
            O => \N__30743\,
            I => \N__30737\
        );

    \I__5373\ : InMux
    port map (
            O => \N__30740\,
            I => \N__30734\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__30737\,
            I => \N__30731\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__30734\,
            I => \N__30728\
        );

    \I__5370\ : Span4Mux_h
    port map (
            O => \N__30731\,
            I => \N__30723\
        );

    \I__5369\ : Span4Mux_h
    port map (
            O => \N__30728\,
            I => \N__30723\
        );

    \I__5368\ : Odrv4
    port map (
            O => \N__30723\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__5367\ : InMux
    port map (
            O => \N__30720\,
            I => \N__30717\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__30717\,
            I => \N__30713\
        );

    \I__5365\ : InMux
    port map (
            O => \N__30716\,
            I => \N__30710\
        );

    \I__5364\ : Span4Mux_v
    port map (
            O => \N__30713\,
            I => \N__30707\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__30710\,
            I => \N__30704\
        );

    \I__5362\ : Odrv4
    port map (
            O => \N__30707\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__5361\ : Odrv4
    port map (
            O => \N__30704\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__5360\ : CascadeMux
    port map (
            O => \N__30699\,
            I => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_16_cascade_\
        );

    \I__5359\ : InMux
    port map (
            O => \N__30696\,
            I => \N__30693\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__30693\,
            I => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_25\
        );

    \I__5357\ : CascadeMux
    port map (
            O => \N__30690\,
            I => \N__30687\
        );

    \I__5356\ : InMux
    port map (
            O => \N__30687\,
            I => \N__30681\
        );

    \I__5355\ : CascadeMux
    port map (
            O => \N__30686\,
            I => \N__30678\
        );

    \I__5354\ : CascadeMux
    port map (
            O => \N__30685\,
            I => \N__30674\
        );

    \I__5353\ : CascadeMux
    port map (
            O => \N__30684\,
            I => \N__30658\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__30681\,
            I => \N__30652\
        );

    \I__5351\ : InMux
    port map (
            O => \N__30678\,
            I => \N__30649\
        );

    \I__5350\ : InMux
    port map (
            O => \N__30677\,
            I => \N__30644\
        );

    \I__5349\ : InMux
    port map (
            O => \N__30674\,
            I => \N__30644\
        );

    \I__5348\ : InMux
    port map (
            O => \N__30673\,
            I => \N__30641\
        );

    \I__5347\ : InMux
    port map (
            O => \N__30672\,
            I => \N__30634\
        );

    \I__5346\ : InMux
    port map (
            O => \N__30671\,
            I => \N__30634\
        );

    \I__5345\ : InMux
    port map (
            O => \N__30670\,
            I => \N__30634\
        );

    \I__5344\ : InMux
    port map (
            O => \N__30669\,
            I => \N__30627\
        );

    \I__5343\ : InMux
    port map (
            O => \N__30668\,
            I => \N__30627\
        );

    \I__5342\ : InMux
    port map (
            O => \N__30667\,
            I => \N__30627\
        );

    \I__5341\ : InMux
    port map (
            O => \N__30666\,
            I => \N__30616\
        );

    \I__5340\ : InMux
    port map (
            O => \N__30665\,
            I => \N__30616\
        );

    \I__5339\ : InMux
    port map (
            O => \N__30664\,
            I => \N__30616\
        );

    \I__5338\ : InMux
    port map (
            O => \N__30663\,
            I => \N__30616\
        );

    \I__5337\ : InMux
    port map (
            O => \N__30662\,
            I => \N__30616\
        );

    \I__5336\ : InMux
    port map (
            O => \N__30661\,
            I => \N__30607\
        );

    \I__5335\ : InMux
    port map (
            O => \N__30658\,
            I => \N__30607\
        );

    \I__5334\ : InMux
    port map (
            O => \N__30657\,
            I => \N__30607\
        );

    \I__5333\ : InMux
    port map (
            O => \N__30656\,
            I => \N__30607\
        );

    \I__5332\ : InMux
    port map (
            O => \N__30655\,
            I => \N__30604\
        );

    \I__5331\ : Span4Mux_h
    port map (
            O => \N__30652\,
            I => \N__30597\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__30649\,
            I => \N__30597\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__30644\,
            I => \N__30597\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__30641\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__30634\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__30627\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__30616\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__30607\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__30604\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31\
        );

    \I__5322\ : Odrv4
    port map (
            O => \N__30597\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31\
        );

    \I__5321\ : InMux
    port map (
            O => \N__30582\,
            I => \N__30578\
        );

    \I__5320\ : InMux
    port map (
            O => \N__30581\,
            I => \N__30575\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__30578\,
            I => \elapsed_time_ns_1_RNI3FU8E1_0_20\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__30575\,
            I => \elapsed_time_ns_1_RNI3FU8E1_0_20\
        );

    \I__5317\ : CascadeMux
    port map (
            O => \N__30570\,
            I => \N__30567\
        );

    \I__5316\ : InMux
    port map (
            O => \N__30567\,
            I => \N__30563\
        );

    \I__5315\ : InMux
    port map (
            O => \N__30566\,
            I => \N__30559\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__30563\,
            I => \N__30556\
        );

    \I__5313\ : CascadeMux
    port map (
            O => \N__30562\,
            I => \N__30553\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__30559\,
            I => \N__30548\
        );

    \I__5311\ : Span4Mux_v
    port map (
            O => \N__30556\,
            I => \N__30548\
        );

    \I__5310\ : InMux
    port map (
            O => \N__30553\,
            I => \N__30545\
        );

    \I__5309\ : Odrv4
    port map (
            O => \N__30548\,
            I => \elapsed_time_ns_1_RNI2DT8E1_0_10\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__30545\,
            I => \elapsed_time_ns_1_RNI2DT8E1_0_10\
        );

    \I__5307\ : CascadeMux
    port map (
            O => \N__30540\,
            I => \N__30535\
        );

    \I__5306\ : InMux
    port map (
            O => \N__30539\,
            I => \N__30532\
        );

    \I__5305\ : CascadeMux
    port map (
            O => \N__30538\,
            I => \N__30529\
        );

    \I__5304\ : InMux
    port map (
            O => \N__30535\,
            I => \N__30526\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__30532\,
            I => \N__30523\
        );

    \I__5302\ : InMux
    port map (
            O => \N__30529\,
            I => \N__30519\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__30526\,
            I => \N__30516\
        );

    \I__5300\ : Span4Mux_v
    port map (
            O => \N__30523\,
            I => \N__30513\
        );

    \I__5299\ : InMux
    port map (
            O => \N__30522\,
            I => \N__30510\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__30519\,
            I => \elapsed_time_ns_1_RNI3ET8E1_0_11\
        );

    \I__5297\ : Odrv12
    port map (
            O => \N__30516\,
            I => \elapsed_time_ns_1_RNI3ET8E1_0_11\
        );

    \I__5296\ : Odrv4
    port map (
            O => \N__30513\,
            I => \elapsed_time_ns_1_RNI3ET8E1_0_11\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__30510\,
            I => \elapsed_time_ns_1_RNI3ET8E1_0_11\
        );

    \I__5294\ : CascadeMux
    port map (
            O => \N__30501\,
            I => \N__30498\
        );

    \I__5293\ : InMux
    port map (
            O => \N__30498\,
            I => \N__30495\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__30495\,
            I => \N__30490\
        );

    \I__5291\ : InMux
    port map (
            O => \N__30494\,
            I => \N__30486\
        );

    \I__5290\ : InMux
    port map (
            O => \N__30493\,
            I => \N__30483\
        );

    \I__5289\ : Span4Mux_v
    port map (
            O => \N__30490\,
            I => \N__30480\
        );

    \I__5288\ : InMux
    port map (
            O => \N__30489\,
            I => \N__30477\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__30486\,
            I => \elapsed_time_ns_1_RNI4FT8E1_0_12\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__30483\,
            I => \elapsed_time_ns_1_RNI4FT8E1_0_12\
        );

    \I__5285\ : Odrv4
    port map (
            O => \N__30480\,
            I => \elapsed_time_ns_1_RNI4FT8E1_0_12\
        );

    \I__5284\ : LocalMux
    port map (
            O => \N__30477\,
            I => \elapsed_time_ns_1_RNI4FT8E1_0_12\
        );

    \I__5283\ : InMux
    port map (
            O => \N__30468\,
            I => \N__30464\
        );

    \I__5282\ : InMux
    port map (
            O => \N__30467\,
            I => \N__30461\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__30464\,
            I => \elapsed_time_ns_1_RNI4GU8E1_0_21\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__30461\,
            I => \elapsed_time_ns_1_RNI4GU8E1_0_21\
        );

    \I__5279\ : CascadeMux
    port map (
            O => \N__30456\,
            I => \elapsed_time_ns_1_RNICOU8E1_0_29_cascade_\
        );

    \I__5278\ : InMux
    port map (
            O => \N__30453\,
            I => \N__30450\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__30450\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15\
        );

    \I__5276\ : CascadeMux
    port map (
            O => \N__30447\,
            I => \N__30444\
        );

    \I__5275\ : InMux
    port map (
            O => \N__30444\,
            I => \N__30437\
        );

    \I__5274\ : InMux
    port map (
            O => \N__30443\,
            I => \N__30437\
        );

    \I__5273\ : InMux
    port map (
            O => \N__30442\,
            I => \N__30434\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__30437\,
            I => \N__30429\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__30434\,
            I => \N__30426\
        );

    \I__5270\ : InMux
    port map (
            O => \N__30433\,
            I => \N__30423\
        );

    \I__5269\ : InMux
    port map (
            O => \N__30432\,
            I => \N__30420\
        );

    \I__5268\ : Span4Mux_v
    port map (
            O => \N__30429\,
            I => \N__30415\
        );

    \I__5267\ : Span4Mux_h
    port map (
            O => \N__30426\,
            I => \N__30415\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__30423\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__30420\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__5264\ : Odrv4
    port map (
            O => \N__30415\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__5263\ : InMux
    port map (
            O => \N__30408\,
            I => \N__30402\
        );

    \I__5262\ : InMux
    port map (
            O => \N__30407\,
            I => \N__30402\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__30402\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\
        );

    \I__5260\ : CascadeMux
    port map (
            O => \N__30399\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\
        );

    \I__5259\ : InMux
    port map (
            O => \N__30396\,
            I => \N__30393\
        );

    \I__5258\ : LocalMux
    port map (
            O => \N__30393\,
            I => \N__30386\
        );

    \I__5257\ : InMux
    port map (
            O => \N__30392\,
            I => \N__30377\
        );

    \I__5256\ : InMux
    port map (
            O => \N__30391\,
            I => \N__30377\
        );

    \I__5255\ : InMux
    port map (
            O => \N__30390\,
            I => \N__30377\
        );

    \I__5254\ : InMux
    port map (
            O => \N__30389\,
            I => \N__30377\
        );

    \I__5253\ : Span4Mux_h
    port map (
            O => \N__30386\,
            I => \N__30374\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__30377\,
            I => \N__30371\
        );

    \I__5251\ : Odrv4
    port map (
            O => \N__30374\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__5250\ : Odrv12
    port map (
            O => \N__30371\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__5249\ : CascadeMux
    port map (
            O => \N__30366\,
            I => \N__30363\
        );

    \I__5248\ : InMux
    port map (
            O => \N__30363\,
            I => \N__30359\
        );

    \I__5247\ : InMux
    port map (
            O => \N__30362\,
            I => \N__30356\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__30359\,
            I => \elapsed_time_ns_1_RNI8KU8E1_0_25\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__30356\,
            I => \elapsed_time_ns_1_RNI8KU8E1_0_25\
        );

    \I__5244\ : InMux
    port map (
            O => \N__30351\,
            I => \N__30347\
        );

    \I__5243\ : InMux
    port map (
            O => \N__30350\,
            I => \N__30344\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__30347\,
            I => \N__30339\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__30344\,
            I => \N__30339\
        );

    \I__5240\ : Span4Mux_v
    port map (
            O => \N__30339\,
            I => \N__30336\
        );

    \I__5239\ : Odrv4
    port map (
            O => \N__30336\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__5238\ : CascadeMux
    port map (
            O => \N__30333\,
            I => \elapsed_time_ns_1_RNI2DT8E1_0_10_cascade_\
        );

    \I__5237\ : CascadeMux
    port map (
            O => \N__30330\,
            I => \N__30327\
        );

    \I__5236\ : InMux
    port map (
            O => \N__30327\,
            I => \N__30324\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__30324\,
            I => \N__30319\
        );

    \I__5234\ : InMux
    port map (
            O => \N__30323\,
            I => \N__30316\
        );

    \I__5233\ : InMux
    port map (
            O => \N__30322\,
            I => \N__30313\
        );

    \I__5232\ : Span4Mux_h
    port map (
            O => \N__30319\,
            I => \N__30310\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__30316\,
            I => \N__30305\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__30313\,
            I => \N__30305\
        );

    \I__5229\ : Odrv4
    port map (
            O => \N__30310\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2\
        );

    \I__5228\ : Odrv4
    port map (
            O => \N__30305\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2\
        );

    \I__5227\ : InMux
    port map (
            O => \N__30300\,
            I => \N__30297\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__30297\,
            I => \N__30293\
        );

    \I__5225\ : InMux
    port map (
            O => \N__30296\,
            I => \N__30290\
        );

    \I__5224\ : Span4Mux_v
    port map (
            O => \N__30293\,
            I => \N__30287\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__30290\,
            I => \N__30284\
        );

    \I__5222\ : Odrv4
    port map (
            O => \N__30287\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__5221\ : Odrv12
    port map (
            O => \N__30284\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__5220\ : InMux
    port map (
            O => \N__30279\,
            I => \N__30273\
        );

    \I__5219\ : InMux
    port map (
            O => \N__30278\,
            I => \N__30273\
        );

    \I__5218\ : LocalMux
    port map (
            O => \N__30273\,
            I => \elapsed_time_ns_1_RNI4HV8E1_0_30\
        );

    \I__5217\ : InMux
    port map (
            O => \N__30270\,
            I => \N__30267\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__30267\,
            I => \N__30264\
        );

    \I__5215\ : Span4Mux_v
    port map (
            O => \N__30264\,
            I => \N__30261\
        );

    \I__5214\ : Odrv4
    port map (
            O => \N__30261\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__5213\ : CascadeMux
    port map (
            O => \N__30258\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_\
        );

    \I__5212\ : CascadeMux
    port map (
            O => \N__30255\,
            I => \N__30248\
        );

    \I__5211\ : InMux
    port map (
            O => \N__30254\,
            I => \N__30245\
        );

    \I__5210\ : InMux
    port map (
            O => \N__30253\,
            I => \N__30242\
        );

    \I__5209\ : InMux
    port map (
            O => \N__30252\,
            I => \N__30239\
        );

    \I__5208\ : InMux
    port map (
            O => \N__30251\,
            I => \N__30233\
        );

    \I__5207\ : InMux
    port map (
            O => \N__30248\,
            I => \N__30233\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__30245\,
            I => \N__30228\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__30242\,
            I => \N__30225\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__30239\,
            I => \N__30222\
        );

    \I__5203\ : InMux
    port map (
            O => \N__30238\,
            I => \N__30219\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__30233\,
            I => \N__30216\
        );

    \I__5201\ : InMux
    port map (
            O => \N__30232\,
            I => \N__30213\
        );

    \I__5200\ : InMux
    port map (
            O => \N__30231\,
            I => \N__30210\
        );

    \I__5199\ : Odrv4
    port map (
            O => \N__30228\,
            I => \delay_measurement_inst.delay_hc_timer.N_342_i\
        );

    \I__5198\ : Odrv4
    port map (
            O => \N__30225\,
            I => \delay_measurement_inst.delay_hc_timer.N_342_i\
        );

    \I__5197\ : Odrv4
    port map (
            O => \N__30222\,
            I => \delay_measurement_inst.delay_hc_timer.N_342_i\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__30219\,
            I => \delay_measurement_inst.delay_hc_timer.N_342_i\
        );

    \I__5195\ : Odrv4
    port map (
            O => \N__30216\,
            I => \delay_measurement_inst.delay_hc_timer.N_342_i\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__30213\,
            I => \delay_measurement_inst.delay_hc_timer.N_342_i\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__30210\,
            I => \delay_measurement_inst.delay_hc_timer.N_342_i\
        );

    \I__5192\ : InMux
    port map (
            O => \N__30195\,
            I => \N__30191\
        );

    \I__5191\ : CascadeMux
    port map (
            O => \N__30194\,
            I => \N__30186\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__30191\,
            I => \N__30183\
        );

    \I__5189\ : InMux
    port map (
            O => \N__30190\,
            I => \N__30178\
        );

    \I__5188\ : InMux
    port map (
            O => \N__30189\,
            I => \N__30178\
        );

    \I__5187\ : InMux
    port map (
            O => \N__30186\,
            I => \N__30175\
        );

    \I__5186\ : Span4Mux_h
    port map (
            O => \N__30183\,
            I => \N__30172\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__30178\,
            I => \N__30169\
        );

    \I__5184\ : LocalMux
    port map (
            O => \N__30175\,
            I => \elapsed_time_ns_1_RNIP93CP1_0_1\
        );

    \I__5183\ : Odrv4
    port map (
            O => \N__30172\,
            I => \elapsed_time_ns_1_RNIP93CP1_0_1\
        );

    \I__5182\ : Odrv4
    port map (
            O => \N__30169\,
            I => \elapsed_time_ns_1_RNIP93CP1_0_1\
        );

    \I__5181\ : InMux
    port map (
            O => \N__30162\,
            I => \N__30159\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__30159\,
            I => \N__30156\
        );

    \I__5179\ : Span4Mux_v
    port map (
            O => \N__30156\,
            I => \N__30151\
        );

    \I__5178\ : InMux
    port map (
            O => \N__30155\,
            I => \N__30144\
        );

    \I__5177\ : InMux
    port map (
            O => \N__30154\,
            I => \N__30144\
        );

    \I__5176\ : Span4Mux_h
    port map (
            O => \N__30151\,
            I => \N__30141\
        );

    \I__5175\ : InMux
    port map (
            O => \N__30150\,
            I => \N__30136\
        );

    \I__5174\ : InMux
    port map (
            O => \N__30149\,
            I => \N__30136\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__30144\,
            I => \elapsed_time_ns_1_RNIRB3CP1_0_3\
        );

    \I__5172\ : Odrv4
    port map (
            O => \N__30141\,
            I => \elapsed_time_ns_1_RNIRB3CP1_0_3\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__30136\,
            I => \elapsed_time_ns_1_RNIRB3CP1_0_3\
        );

    \I__5170\ : CascadeMux
    port map (
            O => \N__30129\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3_cascade_\
        );

    \I__5169\ : InMux
    port map (
            O => \N__30126\,
            I => \N__30123\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__30123\,
            I => \N__30119\
        );

    \I__5167\ : InMux
    port map (
            O => \N__30122\,
            I => \N__30115\
        );

    \I__5166\ : Span4Mux_v
    port map (
            O => \N__30119\,
            I => \N__30111\
        );

    \I__5165\ : InMux
    port map (
            O => \N__30118\,
            I => \N__30108\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__30115\,
            I => \N__30105\
        );

    \I__5163\ : InMux
    port map (
            O => \N__30114\,
            I => \N__30102\
        );

    \I__5162\ : Span4Mux_h
    port map (
            O => \N__30111\,
            I => \N__30099\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__30108\,
            I => \N__30094\
        );

    \I__5160\ : Span4Mux_h
    port map (
            O => \N__30105\,
            I => \N__30094\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__30102\,
            I => \elapsed_time_ns_1_RNIOJKEE1_0_7\
        );

    \I__5158\ : Odrv4
    port map (
            O => \N__30099\,
            I => \elapsed_time_ns_1_RNIOJKEE1_0_7\
        );

    \I__5157\ : Odrv4
    port map (
            O => \N__30094\,
            I => \elapsed_time_ns_1_RNIOJKEE1_0_7\
        );

    \I__5156\ : CascadeMux
    port map (
            O => \N__30087\,
            I => \N__30084\
        );

    \I__5155\ : InMux
    port map (
            O => \N__30084\,
            I => \N__30079\
        );

    \I__5154\ : InMux
    port map (
            O => \N__30083\,
            I => \N__30076\
        );

    \I__5153\ : InMux
    port map (
            O => \N__30082\,
            I => \N__30073\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__30079\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2\
        );

    \I__5151\ : LocalMux
    port map (
            O => \N__30076\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__30073\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2\
        );

    \I__5149\ : CascadeMux
    port map (
            O => \N__30066\,
            I => \N__30059\
        );

    \I__5148\ : InMux
    port map (
            O => \N__30065\,
            I => \N__30052\
        );

    \I__5147\ : InMux
    port map (
            O => \N__30064\,
            I => \N__30052\
        );

    \I__5146\ : InMux
    port map (
            O => \N__30063\,
            I => \N__30048\
        );

    \I__5145\ : InMux
    port map (
            O => \N__30062\,
            I => \N__30045\
        );

    \I__5144\ : InMux
    port map (
            O => \N__30059\,
            I => \N__30042\
        );

    \I__5143\ : InMux
    port map (
            O => \N__30058\,
            I => \N__30039\
        );

    \I__5142\ : InMux
    port map (
            O => \N__30057\,
            I => \N__30036\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__30052\,
            I => \N__30033\
        );

    \I__5140\ : InMux
    port map (
            O => \N__30051\,
            I => \N__30030\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__30048\,
            I => \N__30027\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__30045\,
            I => \N__30022\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__30042\,
            I => \N__30022\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__30039\,
            I => \elapsed_time_ns_1_RNI7IT8E1_0_15\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__30036\,
            I => \elapsed_time_ns_1_RNI7IT8E1_0_15\
        );

    \I__5134\ : Odrv4
    port map (
            O => \N__30033\,
            I => \elapsed_time_ns_1_RNI7IT8E1_0_15\
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__30030\,
            I => \elapsed_time_ns_1_RNI7IT8E1_0_15\
        );

    \I__5132\ : Odrv4
    port map (
            O => \N__30027\,
            I => \elapsed_time_ns_1_RNI7IT8E1_0_15\
        );

    \I__5131\ : Odrv4
    port map (
            O => \N__30022\,
            I => \elapsed_time_ns_1_RNI7IT8E1_0_15\
        );

    \I__5130\ : CascadeMux
    port map (
            O => \N__30009\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_\
        );

    \I__5129\ : CascadeMux
    port map (
            O => \N__30006\,
            I => \N__30002\
        );

    \I__5128\ : InMux
    port map (
            O => \N__30005\,
            I => \N__29996\
        );

    \I__5127\ : InMux
    port map (
            O => \N__30002\,
            I => \N__29996\
        );

    \I__5126\ : InMux
    port map (
            O => \N__30001\,
            I => \N__29993\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__29996\,
            I => \N__29990\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__29993\,
            I => \elapsed_time_ns_1_RNIUE3CP1_0_6\
        );

    \I__5123\ : Odrv4
    port map (
            O => \N__29990\,
            I => \elapsed_time_ns_1_RNIUE3CP1_0_6\
        );

    \I__5122\ : CascadeMux
    port map (
            O => \N__29985\,
            I => \phase_controller_inst1.stoper_hc.N_328_cascade_\
        );

    \I__5121\ : InMux
    port map (
            O => \N__29982\,
            I => \N__29978\
        );

    \I__5120\ : CascadeMux
    port map (
            O => \N__29981\,
            I => \N__29975\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__29978\,
            I => \N__29972\
        );

    \I__5118\ : InMux
    port map (
            O => \N__29975\,
            I => \N__29969\
        );

    \I__5117\ : Span4Mux_h
    port map (
            O => \N__29972\,
            I => \N__29966\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__29969\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__5115\ : Odrv4
    port map (
            O => \N__29966\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__5114\ : CascadeMux
    port map (
            O => \N__29961\,
            I => \N__29957\
        );

    \I__5113\ : InMux
    port map (
            O => \N__29960\,
            I => \N__29952\
        );

    \I__5112\ : InMux
    port map (
            O => \N__29957\,
            I => \N__29952\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__29952\,
            I => \N__29947\
        );

    \I__5110\ : InMux
    port map (
            O => \N__29951\,
            I => \N__29944\
        );

    \I__5109\ : InMux
    port map (
            O => \N__29950\,
            I => \N__29941\
        );

    \I__5108\ : Span4Mux_h
    port map (
            O => \N__29947\,
            I => \N__29938\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__29944\,
            I => \N__29935\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__29941\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__5105\ : Odrv4
    port map (
            O => \N__29938\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__5104\ : Odrv12
    port map (
            O => \N__29935\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__5103\ : InMux
    port map (
            O => \N__29928\,
            I => \N__29925\
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__29925\,
            I => \N__29921\
        );

    \I__5101\ : InMux
    port map (
            O => \N__29924\,
            I => \N__29918\
        );

    \I__5100\ : Span4Mux_v
    port map (
            O => \N__29921\,
            I => \N__29915\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__29918\,
            I => \N__29912\
        );

    \I__5098\ : Odrv4
    port map (
            O => \N__29915\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__5097\ : Odrv12
    port map (
            O => \N__29912\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__5096\ : InMux
    port map (
            O => \N__29907\,
            I => \N__29904\
        );

    \I__5095\ : LocalMux
    port map (
            O => \N__29904\,
            I => \elapsed_time_ns_1_RNICOU8E1_0_29\
        );

    \I__5094\ : InMux
    port map (
            O => \N__29901\,
            I => \N__29898\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__29898\,
            I => \N__29895\
        );

    \I__5092\ : Span4Mux_v
    port map (
            O => \N__29895\,
            I => \N__29892\
        );

    \I__5091\ : Span4Mux_v
    port map (
            O => \N__29892\,
            I => \N__29889\
        );

    \I__5090\ : Odrv4
    port map (
            O => \N__29889\,
            I => \il_min_comp1_D1\
        );

    \I__5089\ : InMux
    port map (
            O => \N__29886\,
            I => \N__29881\
        );

    \I__5088\ : InMux
    port map (
            O => \N__29885\,
            I => \N__29876\
        );

    \I__5087\ : InMux
    port map (
            O => \N__29884\,
            I => \N__29876\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__29881\,
            I => \N__29871\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__29876\,
            I => \N__29871\
        );

    \I__5084\ : Odrv4
    port map (
            O => \N__29871\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_i_0_14\
        );

    \I__5083\ : InMux
    port map (
            O => \N__29868\,
            I => \N__29863\
        );

    \I__5082\ : InMux
    port map (
            O => \N__29867\,
            I => \N__29860\
        );

    \I__5081\ : InMux
    port map (
            O => \N__29866\,
            I => \N__29857\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__29863\,
            I => \N__29854\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__29860\,
            I => \N__29851\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__29857\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\
        );

    \I__5077\ : Odrv4
    port map (
            O => \N__29854\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\
        );

    \I__5076\ : Odrv4
    port map (
            O => \N__29851\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\
        );

    \I__5075\ : InMux
    port map (
            O => \N__29844\,
            I => \N__29841\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__29841\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\
        );

    \I__5073\ : CascadeMux
    port map (
            O => \N__29838\,
            I => \N__29835\
        );

    \I__5072\ : InMux
    port map (
            O => \N__29835\,
            I => \N__29832\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__29832\,
            I => \N__29829\
        );

    \I__5070\ : Odrv4
    port map (
            O => \N__29829\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9JZ0\
        );

    \I__5069\ : InMux
    port map (
            O => \N__29826\,
            I => \N__29822\
        );

    \I__5068\ : InMux
    port map (
            O => \N__29825\,
            I => \N__29819\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__29822\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__29819\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\
        );

    \I__5065\ : InMux
    port map (
            O => \N__29814\,
            I => \N__29810\
        );

    \I__5064\ : InMux
    port map (
            O => \N__29813\,
            I => \N__29807\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__29810\,
            I => \N__29801\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__29807\,
            I => \N__29798\
        );

    \I__5061\ : InMux
    port map (
            O => \N__29806\,
            I => \N__29795\
        );

    \I__5060\ : InMux
    port map (
            O => \N__29805\,
            I => \N__29792\
        );

    \I__5059\ : InMux
    port map (
            O => \N__29804\,
            I => \N__29789\
        );

    \I__5058\ : Span4Mux_v
    port map (
            O => \N__29801\,
            I => \N__29784\
        );

    \I__5057\ : Span4Mux_v
    port map (
            O => \N__29798\,
            I => \N__29784\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__29795\,
            I => \N__29779\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__29792\,
            I => \N__29779\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__29789\,
            I => \N__29776\
        );

    \I__5053\ : Span4Mux_h
    port map (
            O => \N__29784\,
            I => \N__29773\
        );

    \I__5052\ : Span4Mux_v
    port map (
            O => \N__29779\,
            I => \N__29770\
        );

    \I__5051\ : Odrv12
    port map (
            O => \N__29776\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__5050\ : Odrv4
    port map (
            O => \N__29773\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__5049\ : Odrv4
    port map (
            O => \N__29770\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__5048\ : CascadeMux
    port map (
            O => \N__29763\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27_cascade_\
        );

    \I__5047\ : InMux
    port map (
            O => \N__29760\,
            I => \N__29757\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__29757\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\
        );

    \I__5045\ : CascadeMux
    port map (
            O => \N__29754\,
            I => \N__29751\
        );

    \I__5044\ : InMux
    port map (
            O => \N__29751\,
            I => \N__29748\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__29748\,
            I => \N__29745\
        );

    \I__5042\ : Odrv12
    port map (
            O => \N__29745\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7JZ0\
        );

    \I__5041\ : InMux
    port map (
            O => \N__29742\,
            I => \N__29738\
        );

    \I__5040\ : CascadeMux
    port map (
            O => \N__29741\,
            I => \N__29735\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__29738\,
            I => \N__29732\
        );

    \I__5038\ : InMux
    port map (
            O => \N__29735\,
            I => \N__29729\
        );

    \I__5037\ : Span4Mux_v
    port map (
            O => \N__29732\,
            I => \N__29726\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__29729\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__5035\ : Odrv4
    port map (
            O => \N__29726\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__5034\ : InMux
    port map (
            O => \N__29721\,
            I => \N__29717\
        );

    \I__5033\ : InMux
    port map (
            O => \N__29720\,
            I => \N__29714\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__29717\,
            I => \N__29711\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__29714\,
            I => \N__29708\
        );

    \I__5030\ : Span4Mux_v
    port map (
            O => \N__29711\,
            I => \N__29703\
        );

    \I__5029\ : Span4Mux_v
    port map (
            O => \N__29708\,
            I => \N__29703\
        );

    \I__5028\ : Odrv4
    port map (
            O => \N__29703\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__5027\ : InMux
    port map (
            O => \N__29700\,
            I => \N__29697\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__29697\,
            I => \N__29694\
        );

    \I__5025\ : Span4Mux_h
    port map (
            O => \N__29694\,
            I => \N__29691\
        );

    \I__5024\ : Odrv4
    port map (
            O => \N__29691\,
            I => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_15\
        );

    \I__5023\ : InMux
    port map (
            O => \N__29688\,
            I => \N__29684\
        );

    \I__5022\ : InMux
    port map (
            O => \N__29687\,
            I => \N__29681\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__29684\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__29681\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2\
        );

    \I__5019\ : CascadeMux
    port map (
            O => \N__29676\,
            I => \N__29673\
        );

    \I__5018\ : InMux
    port map (
            O => \N__29673\,
            I => \N__29670\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__29670\,
            I => \N__29667\
        );

    \I__5016\ : Odrv4
    port map (
            O => \N__29667\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3\
        );

    \I__5015\ : InMux
    port map (
            O => \N__29664\,
            I => \N__29660\
        );

    \I__5014\ : InMux
    port map (
            O => \N__29663\,
            I => \N__29657\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__29660\,
            I => \N__29652\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__29657\,
            I => \N__29652\
        );

    \I__5011\ : Span4Mux_h
    port map (
            O => \N__29652\,
            I => \N__29648\
        );

    \I__5010\ : InMux
    port map (
            O => \N__29651\,
            I => \N__29645\
        );

    \I__5009\ : Span4Mux_h
    port map (
            O => \N__29648\,
            I => \N__29642\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__29645\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\
        );

    \I__5007\ : Odrv4
    port map (
            O => \N__29642\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\
        );

    \I__5006\ : CascadeMux
    port map (
            O => \N__29637\,
            I => \N__29634\
        );

    \I__5005\ : InMux
    port map (
            O => \N__29634\,
            I => \N__29631\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__29631\,
            I => \N__29628\
        );

    \I__5003\ : Sp12to4
    port map (
            O => \N__29628\,
            I => \N__29625\
        );

    \I__5002\ : Odrv12
    port map (
            O => \N__29625\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO\
        );

    \I__5001\ : InMux
    port map (
            O => \N__29622\,
            I => \bfn_11_11_0_\
        );

    \I__5000\ : InMux
    port map (
            O => \N__29619\,
            I => \N__29616\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__29616\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO\
        );

    \I__4998\ : InMux
    port map (
            O => \N__29613\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\
        );

    \I__4997\ : InMux
    port map (
            O => \N__29610\,
            I => \N__29606\
        );

    \I__4996\ : InMux
    port map (
            O => \N__29609\,
            I => \N__29603\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__29606\,
            I => \N__29598\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__29603\,
            I => \N__29598\
        );

    \I__4993\ : Span4Mux_h
    port map (
            O => \N__29598\,
            I => \N__29594\
        );

    \I__4992\ : InMux
    port map (
            O => \N__29597\,
            I => \N__29591\
        );

    \I__4991\ : Span4Mux_h
    port map (
            O => \N__29594\,
            I => \N__29588\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__29591\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\
        );

    \I__4989\ : Odrv4
    port map (
            O => \N__29588\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\
        );

    \I__4988\ : InMux
    port map (
            O => \N__29583\,
            I => \N__29580\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__29580\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\
        );

    \I__4986\ : InMux
    port map (
            O => \N__29577\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\
        );

    \I__4985\ : InMux
    port map (
            O => \N__29574\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\
        );

    \I__4984\ : InMux
    port map (
            O => \N__29571\,
            I => \N__29568\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__29568\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\
        );

    \I__4982\ : InMux
    port map (
            O => \N__29565\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\
        );

    \I__4981\ : InMux
    port map (
            O => \N__29562\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\
        );

    \I__4980\ : InMux
    port map (
            O => \N__29559\,
            I => \N__29556\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__29556\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\
        );

    \I__4978\ : InMux
    port map (
            O => \N__29553\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\
        );

    \I__4977\ : InMux
    port map (
            O => \N__29550\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_31\
        );

    \I__4976\ : CascadeMux
    port map (
            O => \N__29547\,
            I => \N__29544\
        );

    \I__4975\ : InMux
    port map (
            O => \N__29544\,
            I => \N__29541\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__29541\,
            I => \N__29538\
        );

    \I__4973\ : Span4Mux_h
    port map (
            O => \N__29538\,
            I => \N__29535\
        );

    \I__4972\ : Odrv4
    port map (
            O => \N__29535\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74KZ0\
        );

    \I__4971\ : CascadeMux
    port map (
            O => \N__29532\,
            I => \N__29529\
        );

    \I__4970\ : InMux
    port map (
            O => \N__29529\,
            I => \N__29526\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__29526\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO\
        );

    \I__4968\ : InMux
    port map (
            O => \N__29523\,
            I => \bfn_11_10_0_\
        );

    \I__4967\ : InMux
    port map (
            O => \N__29520\,
            I => \N__29517\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__29517\,
            I => \N__29512\
        );

    \I__4965\ : InMux
    port map (
            O => \N__29516\,
            I => \N__29509\
        );

    \I__4964\ : InMux
    port map (
            O => \N__29515\,
            I => \N__29506\
        );

    \I__4963\ : Sp12to4
    port map (
            O => \N__29512\,
            I => \N__29501\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__29509\,
            I => \N__29501\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__29506\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\
        );

    \I__4960\ : Odrv12
    port map (
            O => \N__29501\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\
        );

    \I__4959\ : CascadeMux
    port map (
            O => \N__29496\,
            I => \N__29493\
        );

    \I__4958\ : InMux
    port map (
            O => \N__29493\,
            I => \N__29490\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__29490\,
            I => \N__29487\
        );

    \I__4956\ : Odrv4
    port map (
            O => \N__29487\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO\
        );

    \I__4955\ : InMux
    port map (
            O => \N__29484\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\
        );

    \I__4954\ : CascadeMux
    port map (
            O => \N__29481\,
            I => \N__29478\
        );

    \I__4953\ : InMux
    port map (
            O => \N__29478\,
            I => \N__29475\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__29475\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO\
        );

    \I__4951\ : InMux
    port map (
            O => \N__29472\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\
        );

    \I__4950\ : InMux
    port map (
            O => \N__29469\,
            I => \N__29466\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__29466\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO\
        );

    \I__4948\ : InMux
    port map (
            O => \N__29463\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\
        );

    \I__4947\ : InMux
    port map (
            O => \N__29460\,
            I => \N__29456\
        );

    \I__4946\ : InMux
    port map (
            O => \N__29459\,
            I => \N__29453\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__29456\,
            I => \N__29450\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__29453\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\
        );

    \I__4943\ : Odrv4
    port map (
            O => \N__29450\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\
        );

    \I__4942\ : InMux
    port map (
            O => \N__29445\,
            I => \N__29442\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__29442\,
            I => \N__29439\
        );

    \I__4940\ : Odrv4
    port map (
            O => \N__29439\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO\
        );

    \I__4939\ : InMux
    port map (
            O => \N__29436\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\
        );

    \I__4938\ : InMux
    port map (
            O => \N__29433\,
            I => \N__29430\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__29430\,
            I => \N__29425\
        );

    \I__4936\ : InMux
    port map (
            O => \N__29429\,
            I => \N__29422\
        );

    \I__4935\ : InMux
    port map (
            O => \N__29428\,
            I => \N__29419\
        );

    \I__4934\ : Span4Mux_v
    port map (
            O => \N__29425\,
            I => \N__29416\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__29422\,
            I => \N__29413\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__29419\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\
        );

    \I__4931\ : Odrv4
    port map (
            O => \N__29416\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\
        );

    \I__4930\ : Odrv12
    port map (
            O => \N__29413\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\
        );

    \I__4929\ : InMux
    port map (
            O => \N__29406\,
            I => \N__29403\
        );

    \I__4928\ : LocalMux
    port map (
            O => \N__29403\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO\
        );

    \I__4927\ : InMux
    port map (
            O => \N__29400\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\
        );

    \I__4926\ : InMux
    port map (
            O => \N__29397\,
            I => \N__29393\
        );

    \I__4925\ : InMux
    port map (
            O => \N__29396\,
            I => \N__29390\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__29393\,
            I => \N__29384\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__29390\,
            I => \N__29384\
        );

    \I__4922\ : InMux
    port map (
            O => \N__29389\,
            I => \N__29381\
        );

    \I__4921\ : Span4Mux_v
    port map (
            O => \N__29384\,
            I => \N__29378\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__29381\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\
        );

    \I__4919\ : Odrv4
    port map (
            O => \N__29378\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\
        );

    \I__4918\ : InMux
    port map (
            O => \N__29373\,
            I => \N__29370\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__29370\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO\
        );

    \I__4916\ : InMux
    port map (
            O => \N__29367\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\
        );

    \I__4915\ : InMux
    port map (
            O => \N__29364\,
            I => \N__29359\
        );

    \I__4914\ : InMux
    port map (
            O => \N__29363\,
            I => \N__29356\
        );

    \I__4913\ : InMux
    port map (
            O => \N__29362\,
            I => \N__29353\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__29359\,
            I => \N__29348\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__29356\,
            I => \N__29348\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__29353\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\
        );

    \I__4909\ : Odrv4
    port map (
            O => \N__29348\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\
        );

    \I__4908\ : CascadeMux
    port map (
            O => \N__29343\,
            I => \N__29340\
        );

    \I__4907\ : InMux
    port map (
            O => \N__29340\,
            I => \N__29337\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__29337\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO\
        );

    \I__4905\ : InMux
    port map (
            O => \N__29334\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\
        );

    \I__4904\ : InMux
    port map (
            O => \N__29331\,
            I => \N__29328\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__29328\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_8\
        );

    \I__4902\ : InMux
    port map (
            O => \N__29325\,
            I => \bfn_11_9_0_\
        );

    \I__4901\ : InMux
    port map (
            O => \N__29322\,
            I => \N__29319\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__29319\,
            I => \N__29316\
        );

    \I__4899\ : Span4Mux_h
    port map (
            O => \N__29316\,
            I => \N__29313\
        );

    \I__4898\ : Odrv4
    port map (
            O => \N__29313\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_9\
        );

    \I__4897\ : InMux
    port map (
            O => \N__29310\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\
        );

    \I__4896\ : CascadeMux
    port map (
            O => \N__29307\,
            I => \N__29304\
        );

    \I__4895\ : InMux
    port map (
            O => \N__29304\,
            I => \N__29301\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__29301\,
            I => \N__29298\
        );

    \I__4893\ : Odrv4
    port map (
            O => \N__29298\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_10\
        );

    \I__4892\ : InMux
    port map (
            O => \N__29295\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\
        );

    \I__4891\ : InMux
    port map (
            O => \N__29292\,
            I => \N__29289\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__29289\,
            I => \N__29286\
        );

    \I__4889\ : Odrv4
    port map (
            O => \N__29286\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_11\
        );

    \I__4888\ : InMux
    port map (
            O => \N__29283\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\
        );

    \I__4887\ : CascadeMux
    port map (
            O => \N__29280\,
            I => \N__29277\
        );

    \I__4886\ : InMux
    port map (
            O => \N__29277\,
            I => \N__29274\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__29274\,
            I => \N__29271\
        );

    \I__4884\ : Odrv4
    port map (
            O => \N__29271\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_12\
        );

    \I__4883\ : InMux
    port map (
            O => \N__29268\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\
        );

    \I__4882\ : InMux
    port map (
            O => \N__29265\,
            I => \N__29262\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__29262\,
            I => \N__29259\
        );

    \I__4880\ : Span4Mux_h
    port map (
            O => \N__29259\,
            I => \N__29256\
        );

    \I__4879\ : Odrv4
    port map (
            O => \N__29256\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\
        );

    \I__4878\ : InMux
    port map (
            O => \N__29253\,
            I => \N__29250\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__29250\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_13\
        );

    \I__4876\ : InMux
    port map (
            O => \N__29247\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\
        );

    \I__4875\ : InMux
    port map (
            O => \N__29244\,
            I => \N__29241\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__29241\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO\
        );

    \I__4873\ : InMux
    port map (
            O => \N__29238\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\
        );

    \I__4872\ : CascadeMux
    port map (
            O => \N__29235\,
            I => \N__29232\
        );

    \I__4871\ : InMux
    port map (
            O => \N__29232\,
            I => \N__29229\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__29229\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO\
        );

    \I__4869\ : InMux
    port map (
            O => \N__29226\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\
        );

    \I__4868\ : CascadeMux
    port map (
            O => \N__29223\,
            I => \N__29218\
        );

    \I__4867\ : InMux
    port map (
            O => \N__29222\,
            I => \N__29215\
        );

    \I__4866\ : CascadeMux
    port map (
            O => \N__29221\,
            I => \N__29211\
        );

    \I__4865\ : InMux
    port map (
            O => \N__29218\,
            I => \N__29208\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__29215\,
            I => \N__29205\
        );

    \I__4863\ : InMux
    port map (
            O => \N__29214\,
            I => \N__29202\
        );

    \I__4862\ : InMux
    port map (
            O => \N__29211\,
            I => \N__29199\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__29208\,
            I => \N__29196\
        );

    \I__4860\ : Span4Mux_h
    port map (
            O => \N__29205\,
            I => \N__29193\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__29202\,
            I => \N__29190\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__29199\,
            I => \N__29187\
        );

    \I__4857\ : Span4Mux_h
    port map (
            O => \N__29196\,
            I => \N__29184\
        );

    \I__4856\ : Span4Mux_v
    port map (
            O => \N__29193\,
            I => \N__29181\
        );

    \I__4855\ : Span4Mux_v
    port map (
            O => \N__29190\,
            I => \N__29176\
        );

    \I__4854\ : Span4Mux_h
    port map (
            O => \N__29187\,
            I => \N__29176\
        );

    \I__4853\ : Odrv4
    port map (
            O => \N__29184\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__4852\ : Odrv4
    port map (
            O => \N__29181\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__4851\ : Odrv4
    port map (
            O => \N__29176\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__4850\ : CascadeMux
    port map (
            O => \N__29169\,
            I => \N__29166\
        );

    \I__4849\ : InMux
    port map (
            O => \N__29166\,
            I => \N__29163\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__29163\,
            I => \N__29160\
        );

    \I__4847\ : Span12Mux_v
    port map (
            O => \N__29160\,
            I => \N__29157\
        );

    \I__4846\ : Odrv12
    port map (
            O => \N__29157\,
            I => \current_shift_inst.PI_CTRL.integrator_i_28\
        );

    \I__4845\ : InMux
    port map (
            O => \N__29154\,
            I => \N__29151\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__29151\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\
        );

    \I__4843\ : InMux
    port map (
            O => \N__29148\,
            I => \N__29145\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__29145\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\
        );

    \I__4841\ : InMux
    port map (
            O => \N__29142\,
            I => \N__29139\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__29139\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\
        );

    \I__4839\ : InMux
    port map (
            O => \N__29136\,
            I => \N__29133\
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__29133\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\
        );

    \I__4837\ : InMux
    port map (
            O => \N__29130\,
            I => \N__29127\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__29127\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\
        );

    \I__4835\ : InMux
    port map (
            O => \N__29124\,
            I => \N__29121\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__29121\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_4\
        );

    \I__4833\ : InMux
    port map (
            O => \N__29118\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\
        );

    \I__4832\ : InMux
    port map (
            O => \N__29115\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\
        );

    \I__4831\ : InMux
    port map (
            O => \N__29112\,
            I => \N__29109\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__29109\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_6\
        );

    \I__4829\ : InMux
    port map (
            O => \N__29106\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\
        );

    \I__4828\ : InMux
    port map (
            O => \N__29103\,
            I => \N__29100\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__29100\,
            I => \N__29097\
        );

    \I__4826\ : Odrv4
    port map (
            O => \N__29097\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_7\
        );

    \I__4825\ : InMux
    port map (
            O => \N__29094\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\
        );

    \I__4824\ : CascadeMux
    port map (
            O => \N__29091\,
            I => \N__29087\
        );

    \I__4823\ : InMux
    port map (
            O => \N__29090\,
            I => \N__29084\
        );

    \I__4822\ : InMux
    port map (
            O => \N__29087\,
            I => \N__29080\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__29084\,
            I => \N__29077\
        );

    \I__4820\ : InMux
    port map (
            O => \N__29083\,
            I => \N__29074\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__29080\,
            I => \N__29071\
        );

    \I__4818\ : Span4Mux_v
    port map (
            O => \N__29077\,
            I => \N__29066\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__29074\,
            I => \N__29066\
        );

    \I__4816\ : Span4Mux_v
    port map (
            O => \N__29071\,
            I => \N__29061\
        );

    \I__4815\ : Span4Mux_v
    port map (
            O => \N__29066\,
            I => \N__29058\
        );

    \I__4814\ : InMux
    port map (
            O => \N__29065\,
            I => \N__29053\
        );

    \I__4813\ : InMux
    port map (
            O => \N__29064\,
            I => \N__29053\
        );

    \I__4812\ : Odrv4
    port map (
            O => \N__29061\,
            I => \elapsed_time_ns_1_RNIGGC6P1_0_17\
        );

    \I__4811\ : Odrv4
    port map (
            O => \N__29058\,
            I => \elapsed_time_ns_1_RNIGGC6P1_0_17\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__29053\,
            I => \elapsed_time_ns_1_RNIGGC6P1_0_17\
        );

    \I__4809\ : CascadeMux
    port map (
            O => \N__29046\,
            I => \N__29042\
        );

    \I__4808\ : InMux
    port map (
            O => \N__29045\,
            I => \N__29037\
        );

    \I__4807\ : InMux
    port map (
            O => \N__29042\,
            I => \N__29037\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__29037\,
            I => \N__29034\
        );

    \I__4805\ : Odrv4
    port map (
            O => \N__29034\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__4804\ : InMux
    port map (
            O => \N__29031\,
            I => \N__29028\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__29028\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\
        );

    \I__4802\ : CascadeMux
    port map (
            O => \N__29025\,
            I => \N__29021\
        );

    \I__4801\ : InMux
    port map (
            O => \N__29024\,
            I => \N__29016\
        );

    \I__4800\ : InMux
    port map (
            O => \N__29021\,
            I => \N__29016\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__29016\,
            I => \N__29013\
        );

    \I__4798\ : Odrv4
    port map (
            O => \N__29013\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__4797\ : InMux
    port map (
            O => \N__29010\,
            I => \N__29007\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__29007\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\
        );

    \I__4795\ : CascadeMux
    port map (
            O => \N__29004\,
            I => \N__29000\
        );

    \I__4794\ : CascadeMux
    port map (
            O => \N__29003\,
            I => \N__28994\
        );

    \I__4793\ : InMux
    port map (
            O => \N__29000\,
            I => \N__28991\
        );

    \I__4792\ : InMux
    port map (
            O => \N__28999\,
            I => \N__28988\
        );

    \I__4791\ : InMux
    port map (
            O => \N__28998\,
            I => \N__28985\
        );

    \I__4790\ : InMux
    port map (
            O => \N__28997\,
            I => \N__28982\
        );

    \I__4789\ : InMux
    port map (
            O => \N__28994\,
            I => \N__28979\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__28991\,
            I => \N__28976\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__28988\,
            I => \N__28973\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__28985\,
            I => \N__28970\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__28982\,
            I => \N__28967\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__28979\,
            I => \N__28962\
        );

    \I__4783\ : Span4Mux_h
    port map (
            O => \N__28976\,
            I => \N__28962\
        );

    \I__4782\ : Span4Mux_h
    port map (
            O => \N__28973\,
            I => \N__28957\
        );

    \I__4781\ : Span4Mux_h
    port map (
            O => \N__28970\,
            I => \N__28957\
        );

    \I__4780\ : Odrv4
    port map (
            O => \N__28967\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__4779\ : Odrv4
    port map (
            O => \N__28962\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__4778\ : Odrv4
    port map (
            O => \N__28957\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__4777\ : InMux
    port map (
            O => \N__28950\,
            I => \N__28947\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__28947\,
            I => \N__28944\
        );

    \I__4775\ : Span4Mux_h
    port map (
            O => \N__28944\,
            I => \N__28941\
        );

    \I__4774\ : Odrv4
    port map (
            O => \N__28941\,
            I => \current_shift_inst.PI_CTRL.integrator_i_14\
        );

    \I__4773\ : InMux
    port map (
            O => \N__28938\,
            I => \N__28934\
        );

    \I__4772\ : InMux
    port map (
            O => \N__28937\,
            I => \N__28930\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__28934\,
            I => \N__28926\
        );

    \I__4770\ : InMux
    port map (
            O => \N__28933\,
            I => \N__28923\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__28930\,
            I => \N__28920\
        );

    \I__4768\ : InMux
    port map (
            O => \N__28929\,
            I => \N__28917\
        );

    \I__4767\ : Span4Mux_h
    port map (
            O => \N__28926\,
            I => \N__28914\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__28923\,
            I => \N__28911\
        );

    \I__4765\ : Odrv4
    port map (
            O => \N__28920\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__28917\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__4763\ : Odrv4
    port map (
            O => \N__28914\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__4762\ : Odrv12
    port map (
            O => \N__28911\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__4761\ : InMux
    port map (
            O => \N__28902\,
            I => \N__28899\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__28899\,
            I => \N__28896\
        );

    \I__4759\ : Span4Mux_h
    port map (
            O => \N__28896\,
            I => \N__28893\
        );

    \I__4758\ : Odrv4
    port map (
            O => \N__28893\,
            I => \current_shift_inst.PI_CTRL.integrator_i_2\
        );

    \I__4757\ : InMux
    port map (
            O => \N__28890\,
            I => \N__28884\
        );

    \I__4756\ : InMux
    port map (
            O => \N__28889\,
            I => \N__28884\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__28884\,
            I => \N__28880\
        );

    \I__4754\ : InMux
    port map (
            O => \N__28883\,
            I => \N__28877\
        );

    \I__4753\ : Span4Mux_v
    port map (
            O => \N__28880\,
            I => \N__28874\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__28877\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__4751\ : Odrv4
    port map (
            O => \N__28874\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__4750\ : InMux
    port map (
            O => \N__28869\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__4749\ : InMux
    port map (
            O => \N__28866\,
            I => \N__28860\
        );

    \I__4748\ : InMux
    port map (
            O => \N__28865\,
            I => \N__28860\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__28860\,
            I => \N__28856\
        );

    \I__4746\ : InMux
    port map (
            O => \N__28859\,
            I => \N__28853\
        );

    \I__4745\ : Span4Mux_v
    port map (
            O => \N__28856\,
            I => \N__28850\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__28853\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__4743\ : Odrv4
    port map (
            O => \N__28850\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__4742\ : InMux
    port map (
            O => \N__28845\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__4741\ : CascadeMux
    port map (
            O => \N__28842\,
            I => \N__28838\
        );

    \I__4740\ : CascadeMux
    port map (
            O => \N__28841\,
            I => \N__28835\
        );

    \I__4739\ : InMux
    port map (
            O => \N__28838\,
            I => \N__28832\
        );

    \I__4738\ : InMux
    port map (
            O => \N__28835\,
            I => \N__28829\
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__28832\,
            I => \N__28823\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__28829\,
            I => \N__28823\
        );

    \I__4735\ : InMux
    port map (
            O => \N__28828\,
            I => \N__28820\
        );

    \I__4734\ : Span4Mux_v
    port map (
            O => \N__28823\,
            I => \N__28817\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__28820\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__4732\ : Odrv4
    port map (
            O => \N__28817\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__4731\ : CascadeMux
    port map (
            O => \N__28812\,
            I => \N__28808\
        );

    \I__4730\ : InMux
    port map (
            O => \N__28811\,
            I => \N__28803\
        );

    \I__4729\ : InMux
    port map (
            O => \N__28808\,
            I => \N__28803\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__28803\,
            I => \N__28800\
        );

    \I__4727\ : Odrv12
    port map (
            O => \N__28800\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__4726\ : InMux
    port map (
            O => \N__28797\,
            I => \bfn_10_22_0_\
        );

    \I__4725\ : CascadeMux
    port map (
            O => \N__28794\,
            I => \N__28790\
        );

    \I__4724\ : CascadeMux
    port map (
            O => \N__28793\,
            I => \N__28787\
        );

    \I__4723\ : InMux
    port map (
            O => \N__28790\,
            I => \N__28784\
        );

    \I__4722\ : InMux
    port map (
            O => \N__28787\,
            I => \N__28781\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__28784\,
            I => \N__28776\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__28781\,
            I => \N__28776\
        );

    \I__4719\ : Span4Mux_v
    port map (
            O => \N__28776\,
            I => \N__28772\
        );

    \I__4718\ : InMux
    port map (
            O => \N__28775\,
            I => \N__28769\
        );

    \I__4717\ : Span4Mux_h
    port map (
            O => \N__28772\,
            I => \N__28766\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__28769\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__4715\ : Odrv4
    port map (
            O => \N__28766\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__4714\ : InMux
    port map (
            O => \N__28761\,
            I => \N__28757\
        );

    \I__4713\ : InMux
    port map (
            O => \N__28760\,
            I => \N__28754\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__28757\,
            I => \N__28751\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__28754\,
            I => \N__28748\
        );

    \I__4710\ : Span4Mux_v
    port map (
            O => \N__28751\,
            I => \N__28743\
        );

    \I__4709\ : Span4Mux_v
    port map (
            O => \N__28748\,
            I => \N__28743\
        );

    \I__4708\ : Odrv4
    port map (
            O => \N__28743\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__4707\ : InMux
    port map (
            O => \N__28740\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__4706\ : InMux
    port map (
            O => \N__28737\,
            I => \N__28730\
        );

    \I__4705\ : InMux
    port map (
            O => \N__28736\,
            I => \N__28730\
        );

    \I__4704\ : InMux
    port map (
            O => \N__28735\,
            I => \N__28727\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__28730\,
            I => \N__28724\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__28727\,
            I => \N__28719\
        );

    \I__4701\ : Span4Mux_v
    port map (
            O => \N__28724\,
            I => \N__28719\
        );

    \I__4700\ : Odrv4
    port map (
            O => \N__28719\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__4699\ : CascadeMux
    port map (
            O => \N__28716\,
            I => \N__28713\
        );

    \I__4698\ : InMux
    port map (
            O => \N__28713\,
            I => \N__28710\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__28710\,
            I => \N__28706\
        );

    \I__4696\ : InMux
    port map (
            O => \N__28709\,
            I => \N__28703\
        );

    \I__4695\ : Span4Mux_v
    port map (
            O => \N__28706\,
            I => \N__28700\
        );

    \I__4694\ : LocalMux
    port map (
            O => \N__28703\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__4693\ : Odrv4
    port map (
            O => \N__28700\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__4692\ : InMux
    port map (
            O => \N__28695\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__4691\ : InMux
    port map (
            O => \N__28692\,
            I => \N__28689\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__28689\,
            I => \N__28685\
        );

    \I__4689\ : InMux
    port map (
            O => \N__28688\,
            I => \N__28682\
        );

    \I__4688\ : Span4Mux_v
    port map (
            O => \N__28685\,
            I => \N__28679\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__28682\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__4686\ : Odrv4
    port map (
            O => \N__28679\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__4685\ : CascadeMux
    port map (
            O => \N__28674\,
            I => \N__28671\
        );

    \I__4684\ : InMux
    port map (
            O => \N__28671\,
            I => \N__28667\
        );

    \I__4683\ : InMux
    port map (
            O => \N__28670\,
            I => \N__28664\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__28667\,
            I => \N__28659\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__28664\,
            I => \N__28659\
        );

    \I__4680\ : Span4Mux_h
    port map (
            O => \N__28659\,
            I => \N__28655\
        );

    \I__4679\ : InMux
    port map (
            O => \N__28658\,
            I => \N__28652\
        );

    \I__4678\ : Span4Mux_v
    port map (
            O => \N__28655\,
            I => \N__28649\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__28652\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__4676\ : Odrv4
    port map (
            O => \N__28649\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__4675\ : InMux
    port map (
            O => \N__28644\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__4674\ : InMux
    port map (
            O => \N__28641\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__4673\ : InMux
    port map (
            O => \N__28638\,
            I => \N__28634\
        );

    \I__4672\ : InMux
    port map (
            O => \N__28637\,
            I => \N__28631\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__28634\,
            I => \N__28626\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__28631\,
            I => \N__28626\
        );

    \I__4669\ : Odrv12
    port map (
            O => \N__28626\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__4668\ : CEMux
    port map (
            O => \N__28623\,
            I => \N__28605\
        );

    \I__4667\ : CEMux
    port map (
            O => \N__28622\,
            I => \N__28605\
        );

    \I__4666\ : CEMux
    port map (
            O => \N__28621\,
            I => \N__28605\
        );

    \I__4665\ : CEMux
    port map (
            O => \N__28620\,
            I => \N__28605\
        );

    \I__4664\ : CEMux
    port map (
            O => \N__28619\,
            I => \N__28605\
        );

    \I__4663\ : CEMux
    port map (
            O => \N__28618\,
            I => \N__28605\
        );

    \I__4662\ : GlobalMux
    port map (
            O => \N__28605\,
            I => \N__28602\
        );

    \I__4661\ : gio2CtrlBuf
    port map (
            O => \N__28602\,
            I => \delay_measurement_inst.delay_hc_timer.N_393_i_g\
        );

    \I__4660\ : InMux
    port map (
            O => \N__28599\,
            I => \N__28593\
        );

    \I__4659\ : InMux
    port map (
            O => \N__28598\,
            I => \N__28593\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__28593\,
            I => \N__28590\
        );

    \I__4657\ : Odrv4
    port map (
            O => \N__28590\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__4656\ : CascadeMux
    port map (
            O => \N__28587\,
            I => \N__28583\
        );

    \I__4655\ : CascadeMux
    port map (
            O => \N__28586\,
            I => \N__28580\
        );

    \I__4654\ : InMux
    port map (
            O => \N__28583\,
            I => \N__28575\
        );

    \I__4653\ : InMux
    port map (
            O => \N__28580\,
            I => \N__28575\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__28575\,
            I => \N__28572\
        );

    \I__4651\ : Span4Mux_v
    port map (
            O => \N__28572\,
            I => \N__28568\
        );

    \I__4650\ : InMux
    port map (
            O => \N__28571\,
            I => \N__28565\
        );

    \I__4649\ : Span4Mux_h
    port map (
            O => \N__28568\,
            I => \N__28562\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__28565\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__4647\ : Odrv4
    port map (
            O => \N__28562\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__4646\ : InMux
    port map (
            O => \N__28557\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__4645\ : CascadeMux
    port map (
            O => \N__28554\,
            I => \N__28551\
        );

    \I__4644\ : InMux
    port map (
            O => \N__28551\,
            I => \N__28547\
        );

    \I__4643\ : InMux
    port map (
            O => \N__28550\,
            I => \N__28544\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__28547\,
            I => \N__28541\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__28544\,
            I => \N__28538\
        );

    \I__4640\ : Span4Mux_h
    port map (
            O => \N__28541\,
            I => \N__28532\
        );

    \I__4639\ : Span4Mux_h
    port map (
            O => \N__28538\,
            I => \N__28532\
        );

    \I__4638\ : InMux
    port map (
            O => \N__28537\,
            I => \N__28529\
        );

    \I__4637\ : Span4Mux_v
    port map (
            O => \N__28532\,
            I => \N__28526\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__28529\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__4635\ : Odrv4
    port map (
            O => \N__28526\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__4634\ : InMux
    port map (
            O => \N__28521\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__4633\ : CascadeMux
    port map (
            O => \N__28518\,
            I => \N__28515\
        );

    \I__4632\ : InMux
    port map (
            O => \N__28515\,
            I => \N__28511\
        );

    \I__4631\ : InMux
    port map (
            O => \N__28514\,
            I => \N__28508\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__28511\,
            I => \N__28502\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__28508\,
            I => \N__28502\
        );

    \I__4628\ : InMux
    port map (
            O => \N__28507\,
            I => \N__28499\
        );

    \I__4627\ : Span4Mux_v
    port map (
            O => \N__28502\,
            I => \N__28496\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__28499\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__4625\ : Odrv4
    port map (
            O => \N__28496\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__4624\ : InMux
    port map (
            O => \N__28491\,
            I => \bfn_10_21_0_\
        );

    \I__4623\ : InMux
    port map (
            O => \N__28488\,
            I => \N__28484\
        );

    \I__4622\ : InMux
    port map (
            O => \N__28487\,
            I => \N__28481\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__28484\,
            I => \N__28475\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__28481\,
            I => \N__28475\
        );

    \I__4619\ : InMux
    port map (
            O => \N__28480\,
            I => \N__28472\
        );

    \I__4618\ : Span4Mux_v
    port map (
            O => \N__28475\,
            I => \N__28469\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__28472\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__4616\ : Odrv4
    port map (
            O => \N__28469\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__4615\ : InMux
    port map (
            O => \N__28464\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__4614\ : InMux
    port map (
            O => \N__28461\,
            I => \N__28454\
        );

    \I__4613\ : InMux
    port map (
            O => \N__28460\,
            I => \N__28454\
        );

    \I__4612\ : InMux
    port map (
            O => \N__28459\,
            I => \N__28451\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__28454\,
            I => \N__28448\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__28451\,
            I => \N__28443\
        );

    \I__4609\ : Span4Mux_v
    port map (
            O => \N__28448\,
            I => \N__28443\
        );

    \I__4608\ : Odrv4
    port map (
            O => \N__28443\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__4607\ : InMux
    port map (
            O => \N__28440\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__4606\ : CascadeMux
    port map (
            O => \N__28437\,
            I => \N__28433\
        );

    \I__4605\ : CascadeMux
    port map (
            O => \N__28436\,
            I => \N__28430\
        );

    \I__4604\ : InMux
    port map (
            O => \N__28433\,
            I => \N__28424\
        );

    \I__4603\ : InMux
    port map (
            O => \N__28430\,
            I => \N__28424\
        );

    \I__4602\ : InMux
    port map (
            O => \N__28429\,
            I => \N__28421\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__28424\,
            I => \N__28418\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__28421\,
            I => \N__28413\
        );

    \I__4599\ : Span4Mux_v
    port map (
            O => \N__28418\,
            I => \N__28413\
        );

    \I__4598\ : Odrv4
    port map (
            O => \N__28413\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__4597\ : InMux
    port map (
            O => \N__28410\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__4596\ : CascadeMux
    port map (
            O => \N__28407\,
            I => \N__28403\
        );

    \I__4595\ : CascadeMux
    port map (
            O => \N__28406\,
            I => \N__28400\
        );

    \I__4594\ : InMux
    port map (
            O => \N__28403\,
            I => \N__28395\
        );

    \I__4593\ : InMux
    port map (
            O => \N__28400\,
            I => \N__28395\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__28395\,
            I => \N__28391\
        );

    \I__4591\ : InMux
    port map (
            O => \N__28394\,
            I => \N__28388\
        );

    \I__4590\ : Span4Mux_v
    port map (
            O => \N__28391\,
            I => \N__28385\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__28388\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__4588\ : Odrv4
    port map (
            O => \N__28385\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__4587\ : InMux
    port map (
            O => \N__28380\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__4586\ : CascadeMux
    port map (
            O => \N__28377\,
            I => \N__28374\
        );

    \I__4585\ : InMux
    port map (
            O => \N__28374\,
            I => \N__28370\
        );

    \I__4584\ : InMux
    port map (
            O => \N__28373\,
            I => \N__28367\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__28370\,
            I => \N__28361\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__28367\,
            I => \N__28361\
        );

    \I__4581\ : InMux
    port map (
            O => \N__28366\,
            I => \N__28358\
        );

    \I__4580\ : Span4Mux_v
    port map (
            O => \N__28361\,
            I => \N__28355\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__28358\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__4578\ : Odrv4
    port map (
            O => \N__28355\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__4577\ : InMux
    port map (
            O => \N__28350\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__4576\ : CascadeMux
    port map (
            O => \N__28347\,
            I => \N__28344\
        );

    \I__4575\ : InMux
    port map (
            O => \N__28344\,
            I => \N__28340\
        );

    \I__4574\ : InMux
    port map (
            O => \N__28343\,
            I => \N__28337\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__28340\,
            I => \N__28331\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__28337\,
            I => \N__28331\
        );

    \I__4571\ : InMux
    port map (
            O => \N__28336\,
            I => \N__28328\
        );

    \I__4570\ : Span4Mux_v
    port map (
            O => \N__28331\,
            I => \N__28325\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__28328\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__4568\ : Odrv4
    port map (
            O => \N__28325\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__4567\ : InMux
    port map (
            O => \N__28320\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__4566\ : InMux
    port map (
            O => \N__28317\,
            I => \N__28311\
        );

    \I__4565\ : InMux
    port map (
            O => \N__28316\,
            I => \N__28311\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__28311\,
            I => \N__28307\
        );

    \I__4563\ : InMux
    port map (
            O => \N__28310\,
            I => \N__28304\
        );

    \I__4562\ : Span4Mux_v
    port map (
            O => \N__28307\,
            I => \N__28301\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__28304\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__4560\ : Odrv4
    port map (
            O => \N__28301\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__4559\ : InMux
    port map (
            O => \N__28296\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__4558\ : InMux
    port map (
            O => \N__28293\,
            I => \N__28286\
        );

    \I__4557\ : InMux
    port map (
            O => \N__28292\,
            I => \N__28286\
        );

    \I__4556\ : InMux
    port map (
            O => \N__28291\,
            I => \N__28283\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__28286\,
            I => \N__28280\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__28283\,
            I => \N__28275\
        );

    \I__4553\ : Span4Mux_v
    port map (
            O => \N__28280\,
            I => \N__28275\
        );

    \I__4552\ : Odrv4
    port map (
            O => \N__28275\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__4551\ : InMux
    port map (
            O => \N__28272\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__4550\ : CascadeMux
    port map (
            O => \N__28269\,
            I => \N__28265\
        );

    \I__4549\ : CascadeMux
    port map (
            O => \N__28268\,
            I => \N__28262\
        );

    \I__4548\ : InMux
    port map (
            O => \N__28265\,
            I => \N__28259\
        );

    \I__4547\ : InMux
    port map (
            O => \N__28262\,
            I => \N__28256\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__28259\,
            I => \N__28250\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__28256\,
            I => \N__28250\
        );

    \I__4544\ : InMux
    port map (
            O => \N__28255\,
            I => \N__28247\
        );

    \I__4543\ : Span4Mux_v
    port map (
            O => \N__28250\,
            I => \N__28244\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__28247\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__4541\ : Odrv4
    port map (
            O => \N__28244\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__4540\ : InMux
    port map (
            O => \N__28239\,
            I => \bfn_10_20_0_\
        );

    \I__4539\ : CascadeMux
    port map (
            O => \N__28236\,
            I => \N__28233\
        );

    \I__4538\ : InMux
    port map (
            O => \N__28233\,
            I => \N__28229\
        );

    \I__4537\ : CascadeMux
    port map (
            O => \N__28232\,
            I => \N__28226\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__28229\,
            I => \N__28222\
        );

    \I__4535\ : InMux
    port map (
            O => \N__28226\,
            I => \N__28219\
        );

    \I__4534\ : InMux
    port map (
            O => \N__28225\,
            I => \N__28216\
        );

    \I__4533\ : Span4Mux_h
    port map (
            O => \N__28222\,
            I => \N__28211\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__28219\,
            I => \N__28211\
        );

    \I__4531\ : LocalMux
    port map (
            O => \N__28216\,
            I => \N__28206\
        );

    \I__4530\ : Span4Mux_v
    port map (
            O => \N__28211\,
            I => \N__28206\
        );

    \I__4529\ : Odrv4
    port map (
            O => \N__28206\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__4528\ : InMux
    port map (
            O => \N__28203\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__4527\ : CascadeMux
    port map (
            O => \N__28200\,
            I => \N__28197\
        );

    \I__4526\ : InMux
    port map (
            O => \N__28197\,
            I => \N__28193\
        );

    \I__4525\ : InMux
    port map (
            O => \N__28196\,
            I => \N__28190\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__28193\,
            I => \N__28186\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__28190\,
            I => \N__28183\
        );

    \I__4522\ : InMux
    port map (
            O => \N__28189\,
            I => \N__28180\
        );

    \I__4521\ : Span4Mux_h
    port map (
            O => \N__28186\,
            I => \N__28175\
        );

    \I__4520\ : Span4Mux_h
    port map (
            O => \N__28183\,
            I => \N__28175\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__28180\,
            I => \N__28170\
        );

    \I__4518\ : Span4Mux_v
    port map (
            O => \N__28175\,
            I => \N__28170\
        );

    \I__4517\ : Odrv4
    port map (
            O => \N__28170\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__4516\ : InMux
    port map (
            O => \N__28167\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__4515\ : InMux
    port map (
            O => \N__28164\,
            I => \N__28158\
        );

    \I__4514\ : InMux
    port map (
            O => \N__28163\,
            I => \N__28158\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__28158\,
            I => \N__28155\
        );

    \I__4512\ : Span4Mux_h
    port map (
            O => \N__28155\,
            I => \N__28151\
        );

    \I__4511\ : InMux
    port map (
            O => \N__28154\,
            I => \N__28148\
        );

    \I__4510\ : Span4Mux_v
    port map (
            O => \N__28151\,
            I => \N__28145\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__28148\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__4508\ : Odrv4
    port map (
            O => \N__28145\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__4507\ : InMux
    port map (
            O => \N__28140\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__4506\ : InMux
    port map (
            O => \N__28137\,
            I => \N__28131\
        );

    \I__4505\ : InMux
    port map (
            O => \N__28136\,
            I => \N__28131\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__28131\,
            I => \N__28127\
        );

    \I__4503\ : InMux
    port map (
            O => \N__28130\,
            I => \N__28124\
        );

    \I__4502\ : Span4Mux_v
    port map (
            O => \N__28127\,
            I => \N__28121\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__28124\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__4500\ : Odrv4
    port map (
            O => \N__28121\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__4499\ : InMux
    port map (
            O => \N__28116\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__4498\ : CascadeMux
    port map (
            O => \N__28113\,
            I => \N__28109\
        );

    \I__4497\ : CascadeMux
    port map (
            O => \N__28112\,
            I => \N__28106\
        );

    \I__4496\ : InMux
    port map (
            O => \N__28109\,
            I => \N__28101\
        );

    \I__4495\ : InMux
    port map (
            O => \N__28106\,
            I => \N__28101\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__28101\,
            I => \N__28097\
        );

    \I__4493\ : InMux
    port map (
            O => \N__28100\,
            I => \N__28094\
        );

    \I__4492\ : Span4Mux_v
    port map (
            O => \N__28097\,
            I => \N__28091\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__28094\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__4490\ : Odrv4
    port map (
            O => \N__28091\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__4489\ : InMux
    port map (
            O => \N__28086\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__4488\ : InMux
    port map (
            O => \N__28083\,
            I => \N__28079\
        );

    \I__4487\ : InMux
    port map (
            O => \N__28082\,
            I => \N__28074\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__28079\,
            I => \N__28071\
        );

    \I__4485\ : InMux
    port map (
            O => \N__28078\,
            I => \N__28068\
        );

    \I__4484\ : InMux
    port map (
            O => \N__28077\,
            I => \N__28065\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__28074\,
            I => \elapsed_time_ns_1_RNIMHKEE1_0_5\
        );

    \I__4482\ : Odrv4
    port map (
            O => \N__28071\,
            I => \elapsed_time_ns_1_RNIMHKEE1_0_5\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__28068\,
            I => \elapsed_time_ns_1_RNIMHKEE1_0_5\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__28065\,
            I => \elapsed_time_ns_1_RNIMHKEE1_0_5\
        );

    \I__4479\ : CascadeMux
    port map (
            O => \N__28056\,
            I => \elapsed_time_ns_1_RNI5IV8E1_0_31_cascade_\
        );

    \I__4478\ : InMux
    port map (
            O => \N__28053\,
            I => \N__28050\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__28050\,
            I => \N__28046\
        );

    \I__4476\ : InMux
    port map (
            O => \N__28049\,
            I => \N__28043\
        );

    \I__4475\ : Span4Mux_h
    port map (
            O => \N__28046\,
            I => \N__28037\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__28043\,
            I => \N__28037\
        );

    \I__4473\ : InMux
    port map (
            O => \N__28042\,
            I => \N__28034\
        );

    \I__4472\ : Span4Mux_v
    port map (
            O => \N__28037\,
            I => \N__28031\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__28034\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__4470\ : Odrv4
    port map (
            O => \N__28031\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__4469\ : InMux
    port map (
            O => \N__28026\,
            I => \N__28022\
        );

    \I__4468\ : InMux
    port map (
            O => \N__28025\,
            I => \N__28019\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__28022\,
            I => \N__28016\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__28019\,
            I => \N__28013\
        );

    \I__4465\ : Span4Mux_v
    port map (
            O => \N__28016\,
            I => \N__28008\
        );

    \I__4464\ : Span4Mux_v
    port map (
            O => \N__28013\,
            I => \N__28008\
        );

    \I__4463\ : Odrv4
    port map (
            O => \N__28008\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__4462\ : InMux
    port map (
            O => \N__28005\,
            I => \N__28002\
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__28002\,
            I => \N__27998\
        );

    \I__4460\ : InMux
    port map (
            O => \N__28001\,
            I => \N__27995\
        );

    \I__4459\ : Span4Mux_v
    port map (
            O => \N__27998\,
            I => \N__27990\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__27995\,
            I => \N__27990\
        );

    \I__4457\ : Span4Mux_v
    port map (
            O => \N__27990\,
            I => \N__27986\
        );

    \I__4456\ : InMux
    port map (
            O => \N__27989\,
            I => \N__27983\
        );

    \I__4455\ : Odrv4
    port map (
            O => \N__27986\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__27983\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__4453\ : CascadeMux
    port map (
            O => \N__27978\,
            I => \N__27974\
        );

    \I__4452\ : InMux
    port map (
            O => \N__27977\,
            I => \N__27971\
        );

    \I__4451\ : InMux
    port map (
            O => \N__27974\,
            I => \N__27968\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__27971\,
            I => \N__27965\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__27968\,
            I => \N__27962\
        );

    \I__4448\ : Span4Mux_v
    port map (
            O => \N__27965\,
            I => \N__27959\
        );

    \I__4447\ : Span4Mux_v
    port map (
            O => \N__27962\,
            I => \N__27956\
        );

    \I__4446\ : Odrv4
    port map (
            O => \N__27959\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__4445\ : Odrv4
    port map (
            O => \N__27956\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__4444\ : InMux
    port map (
            O => \N__27951\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__4443\ : CascadeMux
    port map (
            O => \N__27948\,
            I => \N__27944\
        );

    \I__4442\ : InMux
    port map (
            O => \N__27947\,
            I => \N__27941\
        );

    \I__4441\ : InMux
    port map (
            O => \N__27944\,
            I => \N__27938\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__27941\,
            I => \N__27932\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__27938\,
            I => \N__27932\
        );

    \I__4438\ : InMux
    port map (
            O => \N__27937\,
            I => \N__27929\
        );

    \I__4437\ : Span4Mux_h
    port map (
            O => \N__27932\,
            I => \N__27926\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__27929\,
            I => \N__27921\
        );

    \I__4435\ : Span4Mux_v
    port map (
            O => \N__27926\,
            I => \N__27921\
        );

    \I__4434\ : Odrv4
    port map (
            O => \N__27921\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__4433\ : CascadeMux
    port map (
            O => \N__27918\,
            I => \N__27914\
        );

    \I__4432\ : InMux
    port map (
            O => \N__27917\,
            I => \N__27911\
        );

    \I__4431\ : InMux
    port map (
            O => \N__27914\,
            I => \N__27908\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__27911\,
            I => \N__27905\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__27908\,
            I => \N__27900\
        );

    \I__4428\ : Span4Mux_h
    port map (
            O => \N__27905\,
            I => \N__27900\
        );

    \I__4427\ : Odrv4
    port map (
            O => \N__27900\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__4426\ : InMux
    port map (
            O => \N__27897\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__4425\ : CascadeMux
    port map (
            O => \N__27894\,
            I => \N__27890\
        );

    \I__4424\ : CascadeMux
    port map (
            O => \N__27893\,
            I => \N__27887\
        );

    \I__4423\ : InMux
    port map (
            O => \N__27890\,
            I => \N__27882\
        );

    \I__4422\ : InMux
    port map (
            O => \N__27887\,
            I => \N__27882\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__27882\,
            I => \N__27879\
        );

    \I__4420\ : Span4Mux_h
    port map (
            O => \N__27879\,
            I => \N__27875\
        );

    \I__4419\ : InMux
    port map (
            O => \N__27878\,
            I => \N__27872\
        );

    \I__4418\ : Span4Mux_v
    port map (
            O => \N__27875\,
            I => \N__27869\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__27872\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__4416\ : Odrv4
    port map (
            O => \N__27869\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__4415\ : CascadeMux
    port map (
            O => \N__27864\,
            I => \N__27861\
        );

    \I__4414\ : InMux
    port map (
            O => \N__27861\,
            I => \N__27857\
        );

    \I__4413\ : InMux
    port map (
            O => \N__27860\,
            I => \N__27854\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__27857\,
            I => \N__27849\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__27854\,
            I => \N__27849\
        );

    \I__4410\ : Span4Mux_v
    port map (
            O => \N__27849\,
            I => \N__27846\
        );

    \I__4409\ : Odrv4
    port map (
            O => \N__27846\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__4408\ : InMux
    port map (
            O => \N__27843\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__4407\ : CascadeMux
    port map (
            O => \N__27840\,
            I => \N__27836\
        );

    \I__4406\ : CascadeMux
    port map (
            O => \N__27839\,
            I => \N__27833\
        );

    \I__4405\ : InMux
    port map (
            O => \N__27836\,
            I => \N__27828\
        );

    \I__4404\ : InMux
    port map (
            O => \N__27833\,
            I => \N__27828\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__27828\,
            I => \N__27825\
        );

    \I__4402\ : Span4Mux_h
    port map (
            O => \N__27825\,
            I => \N__27821\
        );

    \I__4401\ : InMux
    port map (
            O => \N__27824\,
            I => \N__27818\
        );

    \I__4400\ : Span4Mux_v
    port map (
            O => \N__27821\,
            I => \N__27815\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__27818\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__4398\ : Odrv4
    port map (
            O => \N__27815\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__4397\ : InMux
    port map (
            O => \N__27810\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__4396\ : InMux
    port map (
            O => \N__27807\,
            I => \N__27803\
        );

    \I__4395\ : InMux
    port map (
            O => \N__27806\,
            I => \N__27800\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__27803\,
            I => \elapsed_time_ns_1_RNI7JU8E1_0_24\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__27800\,
            I => \elapsed_time_ns_1_RNI7JU8E1_0_24\
        );

    \I__4392\ : InMux
    port map (
            O => \N__27795\,
            I => \N__27791\
        );

    \I__4391\ : InMux
    port map (
            O => \N__27794\,
            I => \N__27788\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__27791\,
            I => \elapsed_time_ns_1_RNIBNU8E1_0_28\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__27788\,
            I => \elapsed_time_ns_1_RNIBNU8E1_0_28\
        );

    \I__4388\ : CascadeMux
    port map (
            O => \N__27783\,
            I => \delay_measurement_inst.delay_hc_timer.N_365_clk_cascade_\
        );

    \I__4387\ : InMux
    port map (
            O => \N__27780\,
            I => \N__27773\
        );

    \I__4386\ : InMux
    port map (
            O => \N__27779\,
            I => \N__27773\
        );

    \I__4385\ : InMux
    port map (
            O => \N__27778\,
            I => \N__27770\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__27773\,
            I => \delay_measurement_inst.delay_hc_timer.N_367\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__27770\,
            I => \delay_measurement_inst.delay_hc_timer.N_367\
        );

    \I__4382\ : CascadeMux
    port map (
            O => \N__27765\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31_cascade_\
        );

    \I__4381\ : CascadeMux
    port map (
            O => \N__27762\,
            I => \N__27759\
        );

    \I__4380\ : InMux
    port map (
            O => \N__27759\,
            I => \N__27755\
        );

    \I__4379\ : InMux
    port map (
            O => \N__27758\,
            I => \N__27751\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__27755\,
            I => \N__27748\
        );

    \I__4377\ : InMux
    port map (
            O => \N__27754\,
            I => \N__27745\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__27751\,
            I => \N__27735\
        );

    \I__4375\ : Span4Mux_v
    port map (
            O => \N__27748\,
            I => \N__27735\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__27745\,
            I => \N__27735\
        );

    \I__4373\ : InMux
    port map (
            O => \N__27744\,
            I => \N__27731\
        );

    \I__4372\ : InMux
    port map (
            O => \N__27743\,
            I => \N__27728\
        );

    \I__4371\ : InMux
    port map (
            O => \N__27742\,
            I => \N__27725\
        );

    \I__4370\ : Span4Mux_v
    port map (
            O => \N__27735\,
            I => \N__27722\
        );

    \I__4369\ : InMux
    port map (
            O => \N__27734\,
            I => \N__27719\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__27731\,
            I => \N__27714\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__27728\,
            I => \N__27714\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__27725\,
            I => \elapsed_time_ns_1_RNIDDC6P1_0_14\
        );

    \I__4365\ : Odrv4
    port map (
            O => \N__27722\,
            I => \elapsed_time_ns_1_RNIDDC6P1_0_14\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__27719\,
            I => \elapsed_time_ns_1_RNIDDC6P1_0_14\
        );

    \I__4363\ : Odrv4
    port map (
            O => \N__27714\,
            I => \elapsed_time_ns_1_RNIDDC6P1_0_14\
        );

    \I__4362\ : InMux
    port map (
            O => \N__27705\,
            I => \N__27702\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__27702\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14\
        );

    \I__4360\ : CascadeMux
    port map (
            O => \N__27699\,
            I => \elapsed_time_ns_1_RNI6IU8E1_0_23_cascade_\
        );

    \I__4359\ : CascadeMux
    port map (
            O => \N__27696\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15_cascade_\
        );

    \I__4358\ : InMux
    port map (
            O => \N__27693\,
            I => \N__27690\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__27690\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15\
        );

    \I__4356\ : InMux
    port map (
            O => \N__27687\,
            I => \N__27684\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__27684\,
            I => \N__27681\
        );

    \I__4354\ : Odrv4
    port map (
            O => \N__27681\,
            I => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_1\
        );

    \I__4353\ : CascadeMux
    port map (
            O => \N__27678\,
            I => \N__27675\
        );

    \I__4352\ : InMux
    port map (
            O => \N__27675\,
            I => \N__27671\
        );

    \I__4351\ : InMux
    port map (
            O => \N__27674\,
            I => \N__27668\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__27671\,
            I => \elapsed_time_ns_1_RNI9LU8E1_0_26\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__27668\,
            I => \elapsed_time_ns_1_RNI9LU8E1_0_26\
        );

    \I__4348\ : CascadeMux
    port map (
            O => \N__27663\,
            I => \N__27660\
        );

    \I__4347\ : InMux
    port map (
            O => \N__27660\,
            I => \N__27657\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__27657\,
            I => \N__27654\
        );

    \I__4345\ : Odrv12
    port map (
            O => \N__27654\,
            I => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_14\
        );

    \I__4344\ : InMux
    port map (
            O => \N__27651\,
            I => \N__27648\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__27648\,
            I => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_20\
        );

    \I__4342\ : CascadeMux
    port map (
            O => \N__27645\,
            I => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlt31_0_cascade_\
        );

    \I__4341\ : InMux
    port map (
            O => \N__27642\,
            I => \N__27638\
        );

    \I__4340\ : InMux
    port map (
            O => \N__27641\,
            I => \N__27635\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__27638\,
            I => \elapsed_time_ns_1_RNI5HU8E1_0_22\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__27635\,
            I => \elapsed_time_ns_1_RNI5HU8E1_0_22\
        );

    \I__4337\ : InMux
    port map (
            O => \N__27630\,
            I => \N__27622\
        );

    \I__4336\ : InMux
    port map (
            O => \N__27629\,
            I => \N__27622\
        );

    \I__4335\ : InMux
    port map (
            O => \N__27628\,
            I => \N__27619\
        );

    \I__4334\ : InMux
    port map (
            O => \N__27627\,
            I => \N__27616\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__27622\,
            I => \N__27613\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__27619\,
            I => \N__27608\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__27616\,
            I => \N__27608\
        );

    \I__4330\ : Odrv4
    port map (
            O => \N__27613\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9\
        );

    \I__4329\ : Odrv4
    port map (
            O => \N__27608\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9\
        );

    \I__4328\ : CascadeMux
    port map (
            O => \N__27603\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0Z0Z_6_cascade_\
        );

    \I__4327\ : CascadeMux
    port map (
            O => \N__27600\,
            I => \phase_controller_inst1.stoper_hc.N_326_cascade_\
        );

    \I__4326\ : CascadeMux
    port map (
            O => \N__27597\,
            I => \N__27594\
        );

    \I__4325\ : InMux
    port map (
            O => \N__27594\,
            I => \N__27591\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__27591\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1\
        );

    \I__4323\ : CascadeMux
    port map (
            O => \N__27588\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1_cascade_\
        );

    \I__4322\ : InMux
    port map (
            O => \N__27585\,
            I => \N__27582\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__27582\,
            I => \N__27578\
        );

    \I__4320\ : InMux
    port map (
            O => \N__27581\,
            I => \N__27575\
        );

    \I__4319\ : Odrv4
    port map (
            O => \N__27578\,
            I => \phase_controller_inst1.stoper_hc.N_308\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__27575\,
            I => \phase_controller_inst1.stoper_hc.N_308\
        );

    \I__4317\ : InMux
    port map (
            O => \N__27570\,
            I => \N__27566\
        );

    \I__4316\ : InMux
    port map (
            O => \N__27569\,
            I => \N__27562\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__27566\,
            I => \N__27559\
        );

    \I__4314\ : CascadeMux
    port map (
            O => \N__27565\,
            I => \N__27556\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__27562\,
            I => \N__27553\
        );

    \I__4312\ : Span4Mux_h
    port map (
            O => \N__27559\,
            I => \N__27550\
        );

    \I__4311\ : InMux
    port map (
            O => \N__27556\,
            I => \N__27547\
        );

    \I__4310\ : Odrv4
    port map (
            O => \N__27553\,
            I => \elapsed_time_ns_1_RNILGKEE1_0_4\
        );

    \I__4309\ : Odrv4
    port map (
            O => \N__27550\,
            I => \elapsed_time_ns_1_RNILGKEE1_0_4\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__27547\,
            I => \elapsed_time_ns_1_RNILGKEE1_0_4\
        );

    \I__4307\ : InMux
    port map (
            O => \N__27540\,
            I => \N__27537\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__27537\,
            I => \elapsed_time_ns_1_RNIAMU8E1_0_27\
        );

    \I__4305\ : CascadeMux
    port map (
            O => \N__27534\,
            I => \elapsed_time_ns_1_RNIAMU8E1_0_27_cascade_\
        );

    \I__4304\ : InMux
    port map (
            O => \N__27531\,
            I => \N__27528\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__27528\,
            I => \elapsed_time_ns_1_RNI6IU8E1_0_23\
        );

    \I__4302\ : CascadeMux
    port map (
            O => \N__27525\,
            I => \N__27509\
        );

    \I__4301\ : CascadeMux
    port map (
            O => \N__27524\,
            I => \N__27506\
        );

    \I__4300\ : CascadeMux
    port map (
            O => \N__27523\,
            I => \N__27503\
        );

    \I__4299\ : InMux
    port map (
            O => \N__27522\,
            I => \N__27481\
        );

    \I__4298\ : InMux
    port map (
            O => \N__27521\,
            I => \N__27481\
        );

    \I__4297\ : InMux
    port map (
            O => \N__27520\,
            I => \N__27481\
        );

    \I__4296\ : InMux
    port map (
            O => \N__27519\,
            I => \N__27481\
        );

    \I__4295\ : InMux
    port map (
            O => \N__27518\,
            I => \N__27481\
        );

    \I__4294\ : InMux
    port map (
            O => \N__27517\,
            I => \N__27481\
        );

    \I__4293\ : InMux
    port map (
            O => \N__27516\,
            I => \N__27481\
        );

    \I__4292\ : InMux
    port map (
            O => \N__27515\,
            I => \N__27478\
        );

    \I__4291\ : InMux
    port map (
            O => \N__27514\,
            I => \N__27470\
        );

    \I__4290\ : InMux
    port map (
            O => \N__27513\,
            I => \N__27459\
        );

    \I__4289\ : InMux
    port map (
            O => \N__27512\,
            I => \N__27459\
        );

    \I__4288\ : InMux
    port map (
            O => \N__27509\,
            I => \N__27459\
        );

    \I__4287\ : InMux
    port map (
            O => \N__27506\,
            I => \N__27459\
        );

    \I__4286\ : InMux
    port map (
            O => \N__27503\,
            I => \N__27459\
        );

    \I__4285\ : InMux
    port map (
            O => \N__27502\,
            I => \N__27454\
        );

    \I__4284\ : InMux
    port map (
            O => \N__27501\,
            I => \N__27454\
        );

    \I__4283\ : InMux
    port map (
            O => \N__27500\,
            I => \N__27443\
        );

    \I__4282\ : InMux
    port map (
            O => \N__27499\,
            I => \N__27443\
        );

    \I__4281\ : InMux
    port map (
            O => \N__27498\,
            I => \N__27443\
        );

    \I__4280\ : InMux
    port map (
            O => \N__27497\,
            I => \N__27443\
        );

    \I__4279\ : InMux
    port map (
            O => \N__27496\,
            I => \N__27443\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__27481\,
            I => \N__27440\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__27478\,
            I => \N__27431\
        );

    \I__4276\ : InMux
    port map (
            O => \N__27477\,
            I => \N__27420\
        );

    \I__4275\ : InMux
    port map (
            O => \N__27476\,
            I => \N__27420\
        );

    \I__4274\ : InMux
    port map (
            O => \N__27475\,
            I => \N__27420\
        );

    \I__4273\ : InMux
    port map (
            O => \N__27474\,
            I => \N__27420\
        );

    \I__4272\ : InMux
    port map (
            O => \N__27473\,
            I => \N__27420\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__27470\,
            I => \N__27413\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__27459\,
            I => \N__27413\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__27454\,
            I => \N__27413\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__27443\,
            I => \N__27408\
        );

    \I__4267\ : Span4Mux_h
    port map (
            O => \N__27440\,
            I => \N__27408\
        );

    \I__4266\ : InMux
    port map (
            O => \N__27439\,
            I => \N__27405\
        );

    \I__4265\ : InMux
    port map (
            O => \N__27438\,
            I => \N__27394\
        );

    \I__4264\ : InMux
    port map (
            O => \N__27437\,
            I => \N__27394\
        );

    \I__4263\ : InMux
    port map (
            O => \N__27436\,
            I => \N__27394\
        );

    \I__4262\ : InMux
    port map (
            O => \N__27435\,
            I => \N__27394\
        );

    \I__4261\ : InMux
    port map (
            O => \N__27434\,
            I => \N__27394\
        );

    \I__4260\ : Span4Mux_h
    port map (
            O => \N__27431\,
            I => \N__27391\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__27420\,
            I => \N__27386\
        );

    \I__4258\ : Span4Mux_v
    port map (
            O => \N__27413\,
            I => \N__27386\
        );

    \I__4257\ : Span4Mux_v
    port map (
            O => \N__27408\,
            I => \N__27383\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__27405\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__27394\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__4254\ : Odrv4
    port map (
            O => \N__27391\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__4253\ : Odrv4
    port map (
            O => \N__27386\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__4252\ : Odrv4
    port map (
            O => \N__27383\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__4251\ : InMux
    port map (
            O => \N__27372\,
            I => \N__27362\
        );

    \I__4250\ : InMux
    port map (
            O => \N__27371\,
            I => \N__27362\
        );

    \I__4249\ : InMux
    port map (
            O => \N__27370\,
            I => \N__27362\
        );

    \I__4248\ : InMux
    port map (
            O => \N__27369\,
            I => \N__27340\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__27362\,
            I => \N__27337\
        );

    \I__4246\ : InMux
    port map (
            O => \N__27361\,
            I => \N__27328\
        );

    \I__4245\ : InMux
    port map (
            O => \N__27360\,
            I => \N__27328\
        );

    \I__4244\ : InMux
    port map (
            O => \N__27359\,
            I => \N__27328\
        );

    \I__4243\ : InMux
    port map (
            O => \N__27358\,
            I => \N__27328\
        );

    \I__4242\ : CascadeMux
    port map (
            O => \N__27357\,
            I => \N__27325\
        );

    \I__4241\ : InMux
    port map (
            O => \N__27356\,
            I => \N__27322\
        );

    \I__4240\ : InMux
    port map (
            O => \N__27355\,
            I => \N__27319\
        );

    \I__4239\ : InMux
    port map (
            O => \N__27354\,
            I => \N__27296\
        );

    \I__4238\ : InMux
    port map (
            O => \N__27353\,
            I => \N__27296\
        );

    \I__4237\ : InMux
    port map (
            O => \N__27352\,
            I => \N__27296\
        );

    \I__4236\ : InMux
    port map (
            O => \N__27351\,
            I => \N__27296\
        );

    \I__4235\ : InMux
    port map (
            O => \N__27350\,
            I => \N__27296\
        );

    \I__4234\ : InMux
    port map (
            O => \N__27349\,
            I => \N__27296\
        );

    \I__4233\ : InMux
    port map (
            O => \N__27348\,
            I => \N__27296\
        );

    \I__4232\ : InMux
    port map (
            O => \N__27347\,
            I => \N__27285\
        );

    \I__4231\ : InMux
    port map (
            O => \N__27346\,
            I => \N__27285\
        );

    \I__4230\ : InMux
    port map (
            O => \N__27345\,
            I => \N__27285\
        );

    \I__4229\ : InMux
    port map (
            O => \N__27344\,
            I => \N__27285\
        );

    \I__4228\ : InMux
    port map (
            O => \N__27343\,
            I => \N__27285\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__27340\,
            I => \N__27278\
        );

    \I__4226\ : Span4Mux_v
    port map (
            O => \N__27337\,
            I => \N__27278\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__27328\,
            I => \N__27278\
        );

    \I__4224\ : InMux
    port map (
            O => \N__27325\,
            I => \N__27274\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__27322\,
            I => \N__27271\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__27319\,
            I => \N__27268\
        );

    \I__4221\ : InMux
    port map (
            O => \N__27318\,
            I => \N__27263\
        );

    \I__4220\ : InMux
    port map (
            O => \N__27317\,
            I => \N__27263\
        );

    \I__4219\ : InMux
    port map (
            O => \N__27316\,
            I => \N__27260\
        );

    \I__4218\ : InMux
    port map (
            O => \N__27315\,
            I => \N__27249\
        );

    \I__4217\ : InMux
    port map (
            O => \N__27314\,
            I => \N__27249\
        );

    \I__4216\ : InMux
    port map (
            O => \N__27313\,
            I => \N__27249\
        );

    \I__4215\ : InMux
    port map (
            O => \N__27312\,
            I => \N__27249\
        );

    \I__4214\ : InMux
    port map (
            O => \N__27311\,
            I => \N__27249\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__27296\,
            I => \N__27244\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__27285\,
            I => \N__27244\
        );

    \I__4211\ : Span4Mux_v
    port map (
            O => \N__27278\,
            I => \N__27241\
        );

    \I__4210\ : InMux
    port map (
            O => \N__27277\,
            I => \N__27238\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__27274\,
            I => \N__27233\
        );

    \I__4208\ : Span12Mux_s11_v
    port map (
            O => \N__27271\,
            I => \N__27233\
        );

    \I__4207\ : Sp12to4
    port map (
            O => \N__27268\,
            I => \N__27226\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__27263\,
            I => \N__27226\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__27260\,
            I => \N__27226\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__27249\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4203\ : Odrv4
    port map (
            O => \N__27244\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4202\ : Odrv4
    port map (
            O => \N__27241\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__27238\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4200\ : Odrv12
    port map (
            O => \N__27233\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4199\ : Odrv12
    port map (
            O => \N__27226\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4198\ : CascadeMux
    port map (
            O => \N__27213\,
            I => \N__27210\
        );

    \I__4197\ : InMux
    port map (
            O => \N__27210\,
            I => \N__27207\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__27207\,
            I => \N__27204\
        );

    \I__4195\ : Span4Mux_v
    port map (
            O => \N__27204\,
            I => \N__27201\
        );

    \I__4194\ : Odrv4
    port map (
            O => \N__27201\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__4193\ : CascadeMux
    port map (
            O => \N__27198\,
            I => \N__27192\
        );

    \I__4192\ : CascadeMux
    port map (
            O => \N__27197\,
            I => \N__27184\
        );

    \I__4191\ : CascadeMux
    port map (
            O => \N__27196\,
            I => \N__27181\
        );

    \I__4190\ : CascadeMux
    port map (
            O => \N__27195\,
            I => \N__27178\
        );

    \I__4189\ : InMux
    port map (
            O => \N__27192\,
            I => \N__27171\
        );

    \I__4188\ : CascadeMux
    port map (
            O => \N__27191\,
            I => \N__27157\
        );

    \I__4187\ : CascadeMux
    port map (
            O => \N__27190\,
            I => \N__27154\
        );

    \I__4186\ : CascadeMux
    port map (
            O => \N__27189\,
            I => \N__27151\
        );

    \I__4185\ : InMux
    port map (
            O => \N__27188\,
            I => \N__27140\
        );

    \I__4184\ : InMux
    port map (
            O => \N__27187\,
            I => \N__27140\
        );

    \I__4183\ : InMux
    port map (
            O => \N__27184\,
            I => \N__27140\
        );

    \I__4182\ : InMux
    port map (
            O => \N__27181\,
            I => \N__27140\
        );

    \I__4181\ : InMux
    port map (
            O => \N__27178\,
            I => \N__27140\
        );

    \I__4180\ : CascadeMux
    port map (
            O => \N__27177\,
            I => \N__27134\
        );

    \I__4179\ : CascadeMux
    port map (
            O => \N__27176\,
            I => \N__27129\
        );

    \I__4178\ : CascadeMux
    port map (
            O => \N__27175\,
            I => \N__27123\
        );

    \I__4177\ : CascadeMux
    port map (
            O => \N__27174\,
            I => \N__27120\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__27171\,
            I => \N__27117\
        );

    \I__4175\ : InMux
    port map (
            O => \N__27170\,
            I => \N__27114\
        );

    \I__4174\ : InMux
    port map (
            O => \N__27169\,
            I => \N__27111\
        );

    \I__4173\ : InMux
    port map (
            O => \N__27168\,
            I => \N__27100\
        );

    \I__4172\ : InMux
    port map (
            O => \N__27167\,
            I => \N__27100\
        );

    \I__4171\ : InMux
    port map (
            O => \N__27166\,
            I => \N__27100\
        );

    \I__4170\ : InMux
    port map (
            O => \N__27165\,
            I => \N__27100\
        );

    \I__4169\ : InMux
    port map (
            O => \N__27164\,
            I => \N__27100\
        );

    \I__4168\ : InMux
    port map (
            O => \N__27163\,
            I => \N__27085\
        );

    \I__4167\ : InMux
    port map (
            O => \N__27162\,
            I => \N__27085\
        );

    \I__4166\ : InMux
    port map (
            O => \N__27161\,
            I => \N__27085\
        );

    \I__4165\ : InMux
    port map (
            O => \N__27160\,
            I => \N__27085\
        );

    \I__4164\ : InMux
    port map (
            O => \N__27157\,
            I => \N__27085\
        );

    \I__4163\ : InMux
    port map (
            O => \N__27154\,
            I => \N__27085\
        );

    \I__4162\ : InMux
    port map (
            O => \N__27151\,
            I => \N__27085\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__27140\,
            I => \N__27082\
        );

    \I__4160\ : InMux
    port map (
            O => \N__27139\,
            I => \N__27071\
        );

    \I__4159\ : InMux
    port map (
            O => \N__27138\,
            I => \N__27071\
        );

    \I__4158\ : InMux
    port map (
            O => \N__27137\,
            I => \N__27071\
        );

    \I__4157\ : InMux
    port map (
            O => \N__27134\,
            I => \N__27071\
        );

    \I__4156\ : InMux
    port map (
            O => \N__27133\,
            I => \N__27071\
        );

    \I__4155\ : InMux
    port map (
            O => \N__27132\,
            I => \N__27066\
        );

    \I__4154\ : InMux
    port map (
            O => \N__27129\,
            I => \N__27066\
        );

    \I__4153\ : InMux
    port map (
            O => \N__27128\,
            I => \N__27055\
        );

    \I__4152\ : InMux
    port map (
            O => \N__27127\,
            I => \N__27055\
        );

    \I__4151\ : InMux
    port map (
            O => \N__27126\,
            I => \N__27055\
        );

    \I__4150\ : InMux
    port map (
            O => \N__27123\,
            I => \N__27055\
        );

    \I__4149\ : InMux
    port map (
            O => \N__27120\,
            I => \N__27055\
        );

    \I__4148\ : Span4Mux_v
    port map (
            O => \N__27117\,
            I => \N__27050\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__27114\,
            I => \N__27050\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__27111\,
            I => \N__27043\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__27100\,
            I => \N__27043\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__27085\,
            I => \N__27043\
        );

    \I__4143\ : Span4Mux_v
    port map (
            O => \N__27082\,
            I => \N__27040\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__27071\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__27066\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__27055\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__4139\ : Odrv4
    port map (
            O => \N__27050\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__4138\ : Odrv12
    port map (
            O => \N__27043\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__4137\ : Odrv4
    port map (
            O => \N__27040\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__4136\ : InMux
    port map (
            O => \N__27027\,
            I => \N__27023\
        );

    \I__4135\ : InMux
    port map (
            O => \N__27026\,
            I => \N__27019\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__27023\,
            I => \N__27016\
        );

    \I__4133\ : InMux
    port map (
            O => \N__27022\,
            I => \N__27013\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__27019\,
            I => \N__27010\
        );

    \I__4131\ : Span4Mux_h
    port map (
            O => \N__27016\,
            I => \N__27005\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__27013\,
            I => \N__27002\
        );

    \I__4129\ : Span4Mux_h
    port map (
            O => \N__27010\,
            I => \N__26999\
        );

    \I__4128\ : InMux
    port map (
            O => \N__27009\,
            I => \N__26994\
        );

    \I__4127\ : InMux
    port map (
            O => \N__27008\,
            I => \N__26994\
        );

    \I__4126\ : Span4Mux_h
    port map (
            O => \N__27005\,
            I => \N__26991\
        );

    \I__4125\ : Span12Mux_s11_v
    port map (
            O => \N__27002\,
            I => \N__26988\
        );

    \I__4124\ : Sp12to4
    port map (
            O => \N__26999\,
            I => \N__26983\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__26994\,
            I => \N__26983\
        );

    \I__4122\ : Odrv4
    port map (
            O => \N__26991\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__4121\ : Odrv12
    port map (
            O => \N__26988\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__4120\ : Odrv12
    port map (
            O => \N__26983\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__4119\ : InMux
    port map (
            O => \N__26976\,
            I => \N__26973\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__26973\,
            I => \N__26970\
        );

    \I__4117\ : Span4Mux_h
    port map (
            O => \N__26970\,
            I => \N__26967\
        );

    \I__4116\ : Odrv4
    port map (
            O => \N__26967\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4Z0Z_2\
        );

    \I__4115\ : CascadeMux
    port map (
            O => \N__26964\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2_cascade_\
        );

    \I__4114\ : CascadeMux
    port map (
            O => \N__26961\,
            I => \elapsed_time_ns_1_RNIJEKEE1_0_2_cascade_\
        );

    \I__4113\ : InMux
    port map (
            O => \N__26958\,
            I => \N__26955\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__26955\,
            I => \phase_controller_inst1.stoper_hc.N_284\
        );

    \I__4111\ : CascadeMux
    port map (
            O => \N__26952\,
            I => \N__26949\
        );

    \I__4110\ : InMux
    port map (
            O => \N__26949\,
            I => \N__26943\
        );

    \I__4109\ : InMux
    port map (
            O => \N__26948\,
            I => \N__26943\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__26943\,
            I => \elapsed_time_ns_1_RNIJEKEE1_0_2\
        );

    \I__4107\ : InMux
    port map (
            O => \N__26940\,
            I => \N__26934\
        );

    \I__4106\ : InMux
    port map (
            O => \N__26939\,
            I => \N__26934\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__26934\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__4104\ : InMux
    port map (
            O => \N__26931\,
            I => \N__26927\
        );

    \I__4103\ : InMux
    port map (
            O => \N__26930\,
            I => \N__26924\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__26927\,
            I => \N__26916\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__26924\,
            I => \N__26916\
        );

    \I__4100\ : InMux
    port map (
            O => \N__26923\,
            I => \N__26911\
        );

    \I__4099\ : InMux
    port map (
            O => \N__26922\,
            I => \N__26911\
        );

    \I__4098\ : InMux
    port map (
            O => \N__26921\,
            I => \N__26908\
        );

    \I__4097\ : Span4Mux_v
    port map (
            O => \N__26916\,
            I => \N__26905\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__26911\,
            I => \elapsed_time_ns_1_RNI1I3CP1_0_9\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__26908\,
            I => \elapsed_time_ns_1_RNI1I3CP1_0_9\
        );

    \I__4094\ : Odrv4
    port map (
            O => \N__26905\,
            I => \elapsed_time_ns_1_RNI1I3CP1_0_9\
        );

    \I__4093\ : InMux
    port map (
            O => \N__26898\,
            I => \N__26893\
        );

    \I__4092\ : InMux
    port map (
            O => \N__26897\,
            I => \N__26886\
        );

    \I__4091\ : InMux
    port map (
            O => \N__26896\,
            I => \N__26886\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__26893\,
            I => \N__26883\
        );

    \I__4089\ : InMux
    port map (
            O => \N__26892\,
            I => \N__26878\
        );

    \I__4088\ : InMux
    port map (
            O => \N__26891\,
            I => \N__26878\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__26886\,
            I => \N__26875\
        );

    \I__4086\ : Span4Mux_h
    port map (
            O => \N__26883\,
            I => \N__26872\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__26878\,
            I => \N__26869\
        );

    \I__4084\ : Span4Mux_v
    port map (
            O => \N__26875\,
            I => \N__26866\
        );

    \I__4083\ : Odrv4
    port map (
            O => \N__26872\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__4082\ : Odrv12
    port map (
            O => \N__26869\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__4081\ : Odrv4
    port map (
            O => \N__26866\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__4080\ : InMux
    port map (
            O => \N__26859\,
            I => \N__26856\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__26856\,
            I => \N__26853\
        );

    \I__4078\ : Odrv4
    port map (
            O => \N__26853\,
            I => \current_shift_inst.PI_CTRL.integrator_i_21\
        );

    \I__4077\ : CascadeMux
    port map (
            O => \N__26850\,
            I => \N__26847\
        );

    \I__4076\ : InMux
    port map (
            O => \N__26847\,
            I => \N__26842\
        );

    \I__4075\ : InMux
    port map (
            O => \N__26846\,
            I => \N__26839\
        );

    \I__4074\ : InMux
    port map (
            O => \N__26845\,
            I => \N__26836\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__26842\,
            I => \N__26833\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__26839\,
            I => \N__26828\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__26836\,
            I => \N__26825\
        );

    \I__4070\ : Span4Mux_v
    port map (
            O => \N__26833\,
            I => \N__26822\
        );

    \I__4069\ : InMux
    port map (
            O => \N__26832\,
            I => \N__26817\
        );

    \I__4068\ : InMux
    port map (
            O => \N__26831\,
            I => \N__26817\
        );

    \I__4067\ : Span4Mux_v
    port map (
            O => \N__26828\,
            I => \N__26812\
        );

    \I__4066\ : Span4Mux_v
    port map (
            O => \N__26825\,
            I => \N__26812\
        );

    \I__4065\ : Odrv4
    port map (
            O => \N__26822\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__26817\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__4063\ : Odrv4
    port map (
            O => \N__26812\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__4062\ : CascadeMux
    port map (
            O => \N__26805\,
            I => \N__26802\
        );

    \I__4061\ : InMux
    port map (
            O => \N__26802\,
            I => \N__26799\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__26799\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34JZ0\
        );

    \I__4059\ : CascadeMux
    port map (
            O => \N__26796\,
            I => \N__26793\
        );

    \I__4058\ : InMux
    port map (
            O => \N__26793\,
            I => \N__26790\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__26790\,
            I => \N__26787\
        );

    \I__4056\ : Span4Mux_h
    port map (
            O => \N__26787\,
            I => \N__26784\
        );

    \I__4055\ : Odrv4
    port map (
            O => \N__26784\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI7T941Z0Z_10\
        );

    \I__4054\ : InMux
    port map (
            O => \N__26781\,
            I => \N__26778\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__26778\,
            I => \N__26775\
        );

    \I__4052\ : Span4Mux_h
    port map (
            O => \N__26775\,
            I => \N__26772\
        );

    \I__4051\ : Odrv4
    port map (
            O => \N__26772\,
            I => \current_shift_inst.PI_CTRL.integrator_i_6\
        );

    \I__4050\ : InMux
    port map (
            O => \N__26769\,
            I => \N__26766\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__26766\,
            I => \N__26763\
        );

    \I__4048\ : Odrv4
    port map (
            O => \N__26763\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__4047\ : CascadeMux
    port map (
            O => \N__26760\,
            I => \N__26756\
        );

    \I__4046\ : CascadeMux
    port map (
            O => \N__26759\,
            I => \N__26752\
        );

    \I__4045\ : InMux
    port map (
            O => \N__26756\,
            I => \N__26749\
        );

    \I__4044\ : CascadeMux
    port map (
            O => \N__26755\,
            I => \N__26746\
        );

    \I__4043\ : InMux
    port map (
            O => \N__26752\,
            I => \N__26743\
        );

    \I__4042\ : LocalMux
    port map (
            O => \N__26749\,
            I => \N__26740\
        );

    \I__4041\ : InMux
    port map (
            O => \N__26746\,
            I => \N__26737\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__26743\,
            I => \N__26734\
        );

    \I__4039\ : Span4Mux_v
    port map (
            O => \N__26740\,
            I => \N__26729\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__26737\,
            I => \N__26729\
        );

    \I__4037\ : Span4Mux_v
    port map (
            O => \N__26734\,
            I => \N__26722\
        );

    \I__4036\ : Span4Mux_h
    port map (
            O => \N__26729\,
            I => \N__26722\
        );

    \I__4035\ : InMux
    port map (
            O => \N__26728\,
            I => \N__26717\
        );

    \I__4034\ : InMux
    port map (
            O => \N__26727\,
            I => \N__26717\
        );

    \I__4033\ : Odrv4
    port map (
            O => \N__26722\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__26717\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4031\ : CascadeMux
    port map (
            O => \N__26712\,
            I => \N__26709\
        );

    \I__4030\ : InMux
    port map (
            O => \N__26709\,
            I => \N__26706\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__26706\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__4028\ : InMux
    port map (
            O => \N__26703\,
            I => \N__26700\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__26700\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__4026\ : InMux
    port map (
            O => \N__26697\,
            I => \N__26694\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__26694\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__4024\ : CascadeMux
    port map (
            O => \N__26691\,
            I => \N__26687\
        );

    \I__4023\ : InMux
    port map (
            O => \N__26690\,
            I => \N__26684\
        );

    \I__4022\ : InMux
    port map (
            O => \N__26687\,
            I => \N__26679\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__26684\,
            I => \N__26676\
        );

    \I__4020\ : InMux
    port map (
            O => \N__26683\,
            I => \N__26673\
        );

    \I__4019\ : InMux
    port map (
            O => \N__26682\,
            I => \N__26670\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__26679\,
            I => \N__26667\
        );

    \I__4017\ : Span4Mux_h
    port map (
            O => \N__26676\,
            I => \N__26664\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__26673\,
            I => \N__26659\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__26670\,
            I => \N__26659\
        );

    \I__4014\ : Span4Mux_h
    port map (
            O => \N__26667\,
            I => \N__26654\
        );

    \I__4013\ : Span4Mux_v
    port map (
            O => \N__26664\,
            I => \N__26654\
        );

    \I__4012\ : Odrv12
    port map (
            O => \N__26659\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__4011\ : Odrv4
    port map (
            O => \N__26654\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__4010\ : CascadeMux
    port map (
            O => \N__26649\,
            I => \N__26646\
        );

    \I__4009\ : InMux
    port map (
            O => \N__26646\,
            I => \N__26643\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__26643\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4IZ0\
        );

    \I__4007\ : CascadeMux
    port map (
            O => \N__26640\,
            I => \N__26637\
        );

    \I__4006\ : InMux
    port map (
            O => \N__26637\,
            I => \N__26633\
        );

    \I__4005\ : InMux
    port map (
            O => \N__26636\,
            I => \N__26630\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__26633\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_i_14\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__26630\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_i_14\
        );

    \I__4002\ : CascadeMux
    port map (
            O => \N__26625\,
            I => \N__26622\
        );

    \I__4001\ : InMux
    port map (
            O => \N__26622\,
            I => \N__26619\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__26619\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42IZ0\
        );

    \I__3999\ : CascadeMux
    port map (
            O => \N__26616\,
            I => \N__26613\
        );

    \I__3998\ : InMux
    port map (
            O => \N__26613\,
            I => \N__26610\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__26610\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20JZ0\
        );

    \I__3996\ : CascadeMux
    port map (
            O => \N__26607\,
            I => \N__26604\
        );

    \I__3995\ : InMux
    port map (
            O => \N__26604\,
            I => \N__26601\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__26601\,
            I => \N__26598\
        );

    \I__3993\ : Odrv4
    port map (
            O => \N__26598\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96JZ0\
        );

    \I__3992\ : CascadeMux
    port map (
            O => \N__26595\,
            I => \N__26592\
        );

    \I__3991\ : InMux
    port map (
            O => \N__26592\,
            I => \N__26589\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__26589\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65JZ0\
        );

    \I__3989\ : CascadeMux
    port map (
            O => \N__26586\,
            I => \N__26583\
        );

    \I__3988\ : InMux
    port map (
            O => \N__26583\,
            I => \N__26580\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__26580\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51JZ0\
        );

    \I__3986\ : CascadeMux
    port map (
            O => \N__26577\,
            I => \N__26574\
        );

    \I__3985\ : InMux
    port map (
            O => \N__26574\,
            I => \N__26571\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__26571\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJZ0\
        );

    \I__3983\ : InMux
    port map (
            O => \N__26568\,
            I => \N__26564\
        );

    \I__3982\ : CascadeMux
    port map (
            O => \N__26567\,
            I => \N__26561\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__26564\,
            I => \N__26558\
        );

    \I__3980\ : InMux
    port map (
            O => \N__26561\,
            I => \N__26555\
        );

    \I__3979\ : Span4Mux_v
    port map (
            O => \N__26558\,
            I => \N__26550\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__26555\,
            I => \N__26547\
        );

    \I__3977\ : InMux
    port map (
            O => \N__26554\,
            I => \N__26543\
        );

    \I__3976\ : InMux
    port map (
            O => \N__26553\,
            I => \N__26540\
        );

    \I__3975\ : Span4Mux_v
    port map (
            O => \N__26550\,
            I => \N__26535\
        );

    \I__3974\ : Span4Mux_h
    port map (
            O => \N__26547\,
            I => \N__26535\
        );

    \I__3973\ : InMux
    port map (
            O => \N__26546\,
            I => \N__26532\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__26543\,
            I => \N__26527\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__26540\,
            I => \N__26527\
        );

    \I__3970\ : Odrv4
    port map (
            O => \N__26535\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__26532\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__3968\ : Odrv12
    port map (
            O => \N__26527\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__3967\ : CascadeMux
    port map (
            O => \N__26520\,
            I => \N__26517\
        );

    \I__3966\ : InMux
    port map (
            O => \N__26517\,
            I => \N__26514\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__26514\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8JZ0\
        );

    \I__3964\ : InMux
    port map (
            O => \N__26511\,
            I => \N__26506\
        );

    \I__3963\ : InMux
    port map (
            O => \N__26510\,
            I => \N__26503\
        );

    \I__3962\ : InMux
    port map (
            O => \N__26509\,
            I => \N__26500\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__26506\,
            I => \N__26496\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__26503\,
            I => \N__26493\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__26500\,
            I => \N__26489\
        );

    \I__3958\ : InMux
    port map (
            O => \N__26499\,
            I => \N__26486\
        );

    \I__3957\ : Span4Mux_h
    port map (
            O => \N__26496\,
            I => \N__26481\
        );

    \I__3956\ : Span4Mux_h
    port map (
            O => \N__26493\,
            I => \N__26481\
        );

    \I__3955\ : InMux
    port map (
            O => \N__26492\,
            I => \N__26478\
        );

    \I__3954\ : Span4Mux_h
    port map (
            O => \N__26489\,
            I => \N__26473\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__26486\,
            I => \N__26473\
        );

    \I__3952\ : Odrv4
    port map (
            O => \N__26481\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__26478\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__3950\ : Odrv4
    port map (
            O => \N__26473\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__3949\ : CascadeMux
    port map (
            O => \N__26466\,
            I => \N__26463\
        );

    \I__3948\ : InMux
    port map (
            O => \N__26463\,
            I => \N__26460\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__26460\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIHA7UZ0Z_8\
        );

    \I__3946\ : CascadeMux
    port map (
            O => \N__26457\,
            I => \N__26454\
        );

    \I__3945\ : InMux
    port map (
            O => \N__26454\,
            I => \N__26451\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__26451\,
            I => \N__26448\
        );

    \I__3943\ : Span4Mux_h
    port map (
            O => \N__26448\,
            I => \N__26445\
        );

    \I__3942\ : Odrv4
    port map (
            O => \N__26445\,
            I => \current_shift_inst.PI_CTRL.integrator_i_30\
        );

    \I__3941\ : CascadeMux
    port map (
            O => \N__26442\,
            I => \N__26439\
        );

    \I__3940\ : InMux
    port map (
            O => \N__26439\,
            I => \N__26436\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__26436\,
            I => \N__26433\
        );

    \I__3938\ : Odrv4
    port map (
            O => \N__26433\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI905UZ0Z_6\
        );

    \I__3937\ : CascadeMux
    port map (
            O => \N__26430\,
            I => \N__26427\
        );

    \I__3936\ : InMux
    port map (
            O => \N__26427\,
            I => \N__26424\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__26424\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11IZ0\
        );

    \I__3934\ : InMux
    port map (
            O => \N__26421\,
            I => \N__26417\
        );

    \I__3933\ : CascadeMux
    port map (
            O => \N__26420\,
            I => \N__26412\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__26417\,
            I => \N__26408\
        );

    \I__3931\ : InMux
    port map (
            O => \N__26416\,
            I => \N__26405\
        );

    \I__3930\ : InMux
    port map (
            O => \N__26415\,
            I => \N__26402\
        );

    \I__3929\ : InMux
    port map (
            O => \N__26412\,
            I => \N__26399\
        );

    \I__3928\ : InMux
    port map (
            O => \N__26411\,
            I => \N__26396\
        );

    \I__3927\ : Span4Mux_h
    port map (
            O => \N__26408\,
            I => \N__26391\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__26405\,
            I => \N__26391\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__26402\,
            I => \N__26388\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__26399\,
            I => \N__26385\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__26396\,
            I => \N__26380\
        );

    \I__3922\ : Span4Mux_v
    port map (
            O => \N__26391\,
            I => \N__26380\
        );

    \I__3921\ : Odrv4
    port map (
            O => \N__26388\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__3920\ : Odrv4
    port map (
            O => \N__26385\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__3919\ : Odrv4
    port map (
            O => \N__26380\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__3918\ : CascadeMux
    port map (
            O => \N__26373\,
            I => \N__26370\
        );

    \I__3917\ : InMux
    port map (
            O => \N__26370\,
            I => \N__26367\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__26367\,
            I => \N__26364\
        );

    \I__3915\ : Odrv4
    port map (
            O => \N__26364\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82JZ0\
        );

    \I__3914\ : InMux
    port map (
            O => \N__26361\,
            I => \N__26358\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__26358\,
            I => \N__26354\
        );

    \I__3912\ : InMux
    port map (
            O => \N__26357\,
            I => \N__26351\
        );

    \I__3911\ : Span4Mux_h
    port map (
            O => \N__26354\,
            I => \N__26344\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__26351\,
            I => \N__26344\
        );

    \I__3909\ : InMux
    port map (
            O => \N__26350\,
            I => \N__26339\
        );

    \I__3908\ : InMux
    port map (
            O => \N__26349\,
            I => \N__26339\
        );

    \I__3907\ : Span4Mux_h
    port map (
            O => \N__26344\,
            I => \N__26335\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__26339\,
            I => \N__26332\
        );

    \I__3905\ : InMux
    port map (
            O => \N__26338\,
            I => \N__26329\
        );

    \I__3904\ : Odrv4
    port map (
            O => \N__26335\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__3903\ : Odrv12
    port map (
            O => \N__26332\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__26329\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__3901\ : CascadeMux
    port map (
            O => \N__26322\,
            I => \N__26319\
        );

    \I__3900\ : InMux
    port map (
            O => \N__26319\,
            I => \N__26316\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__26316\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5IZ0\
        );

    \I__3898\ : CascadeMux
    port map (
            O => \N__26313\,
            I => \N__26310\
        );

    \I__3897\ : InMux
    port map (
            O => \N__26310\,
            I => \N__26307\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__26307\,
            I => \N__26304\
        );

    \I__3895\ : Odrv4
    port map (
            O => \N__26304\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73IZ0\
        );

    \I__3894\ : CascadeMux
    port map (
            O => \N__26301\,
            I => \N__26295\
        );

    \I__3893\ : InMux
    port map (
            O => \N__26300\,
            I => \N__26292\
        );

    \I__3892\ : InMux
    port map (
            O => \N__26299\,
            I => \N__26288\
        );

    \I__3891\ : InMux
    port map (
            O => \N__26298\,
            I => \N__26285\
        );

    \I__3890\ : InMux
    port map (
            O => \N__26295\,
            I => \N__26282\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__26292\,
            I => \N__26279\
        );

    \I__3888\ : InMux
    port map (
            O => \N__26291\,
            I => \N__26276\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__26288\,
            I => \N__26273\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__26285\,
            I => \N__26268\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__26282\,
            I => \N__26268\
        );

    \I__3884\ : Span4Mux_h
    port map (
            O => \N__26279\,
            I => \N__26265\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__26276\,
            I => \N__26260\
        );

    \I__3882\ : Span4Mux_h
    port map (
            O => \N__26273\,
            I => \N__26260\
        );

    \I__3881\ : Odrv12
    port map (
            O => \N__26268\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__3880\ : Odrv4
    port map (
            O => \N__26265\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__3879\ : Odrv4
    port map (
            O => \N__26260\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__3878\ : CascadeMux
    port map (
            O => \N__26253\,
            I => \N__26250\
        );

    \I__3877\ : InMux
    port map (
            O => \N__26250\,
            I => \N__26247\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__26247\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIQ6T01Z0Z_13\
        );

    \I__3875\ : InMux
    port map (
            O => \N__26244\,
            I => \N__26241\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__26241\,
            I => \current_shift_inst.PI_CTRL.integrator_i_0\
        );

    \I__3873\ : CascadeMux
    port map (
            O => \N__26238\,
            I => \current_shift_inst.PI_CTRL.integrator_i_0_cascade_\
        );

    \I__3872\ : CascadeMux
    port map (
            O => \N__26235\,
            I => \N__26232\
        );

    \I__3871\ : InMux
    port map (
            O => \N__26232\,
            I => \N__26229\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__26229\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI1M2UZ0Z_4\
        );

    \I__3869\ : InMux
    port map (
            O => \N__26226\,
            I => \N__26223\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__26223\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1\
        );

    \I__3867\ : InMux
    port map (
            O => \N__26220\,
            I => \N__26217\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__26217\,
            I => \current_shift_inst.PI_CTRL.integrator_i_1\
        );

    \I__3865\ : CascadeMux
    port map (
            O => \N__26214\,
            I => \N__26211\
        );

    \I__3864\ : InMux
    port map (
            O => \N__26211\,
            I => \N__26208\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__26208\,
            I => \N__26205\
        );

    \I__3862\ : Span4Mux_v
    port map (
            O => \N__26205\,
            I => \N__26202\
        );

    \I__3861\ : Span4Mux_h
    port map (
            O => \N__26202\,
            I => \N__26197\
        );

    \I__3860\ : InMux
    port map (
            O => \N__26201\,
            I => \N__26192\
        );

    \I__3859\ : InMux
    port map (
            O => \N__26200\,
            I => \N__26192\
        );

    \I__3858\ : Odrv4
    port map (
            O => \N__26197\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__26192\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__3856\ : InMux
    port map (
            O => \N__26187\,
            I => \N__26184\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__26184\,
            I => \current_shift_inst.PI_CTRL.un1_enablelt3_0\
        );

    \I__3854\ : CascadeMux
    port map (
            O => \N__26181\,
            I => \N__26178\
        );

    \I__3853\ : InMux
    port map (
            O => \N__26178\,
            I => \N__26175\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__26175\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVHZ0\
        );

    \I__3851\ : CascadeMux
    port map (
            O => \N__26172\,
            I => \N__26169\
        );

    \I__3850\ : InMux
    port map (
            O => \N__26169\,
            I => \N__26163\
        );

    \I__3849\ : InMux
    port map (
            O => \N__26168\,
            I => \N__26160\
        );

    \I__3848\ : InMux
    port map (
            O => \N__26167\,
            I => \N__26157\
        );

    \I__3847\ : InMux
    port map (
            O => \N__26166\,
            I => \N__26154\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__26163\,
            I => \N__26151\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__26160\,
            I => \N__26146\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__26157\,
            I => \N__26146\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__26154\,
            I => \N__26143\
        );

    \I__3842\ : Span4Mux_v
    port map (
            O => \N__26151\,
            I => \N__26139\
        );

    \I__3841\ : Span12Mux_s10_v
    port map (
            O => \N__26146\,
            I => \N__26136\
        );

    \I__3840\ : Span4Mux_h
    port map (
            O => \N__26143\,
            I => \N__26133\
        );

    \I__3839\ : InMux
    port map (
            O => \N__26142\,
            I => \N__26130\
        );

    \I__3838\ : Odrv4
    port map (
            O => \N__26139\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__3837\ : Odrv12
    port map (
            O => \N__26136\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__3836\ : Odrv4
    port map (
            O => \N__26133\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__26130\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__3834\ : CascadeMux
    port map (
            O => \N__26121\,
            I => \N__26118\
        );

    \I__3833\ : InMux
    port map (
            O => \N__26118\,
            I => \N__26115\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__26115\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIM1S01Z0Z_12\
        );

    \I__3831\ : InMux
    port map (
            O => \N__26112\,
            I => \N__26109\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__26109\,
            I => \current_shift_inst.PI_CTRL.integrator_i_10\
        );

    \I__3829\ : InMux
    port map (
            O => \N__26106\,
            I => \N__26102\
        );

    \I__3828\ : InMux
    port map (
            O => \N__26105\,
            I => \N__26099\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__26102\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__26099\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__3825\ : InMux
    port map (
            O => \N__26094\,
            I => \N__26090\
        );

    \I__3824\ : InMux
    port map (
            O => \N__26093\,
            I => \N__26087\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__26090\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__26087\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__3821\ : InMux
    port map (
            O => \N__26082\,
            I => \N__26079\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__26079\,
            I => \N__26076\
        );

    \I__3819\ : Odrv4
    port map (
            O => \N__26076\,
            I => \phase_controller_inst1.stoper_hc.un4_running_df28\
        );

    \I__3818\ : InMux
    port map (
            O => \N__26073\,
            I => \N__26070\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__26070\,
            I => \N__26067\
        );

    \I__3816\ : Span4Mux_v
    port map (
            O => \N__26067\,
            I => \N__26064\
        );

    \I__3815\ : Odrv4
    port map (
            O => \N__26064\,
            I => \current_shift_inst.PI_CTRL.integrator_i_9\
        );

    \I__3814\ : InMux
    port map (
            O => \N__26061\,
            I => \N__26058\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__26058\,
            I => \N__26055\
        );

    \I__3812\ : Odrv12
    port map (
            O => \N__26055\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\
        );

    \I__3811\ : InMux
    port map (
            O => \N__26052\,
            I => \N__26049\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__26049\,
            I => \N__26046\
        );

    \I__3809\ : Odrv4
    port map (
            O => \N__26046\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\
        );

    \I__3808\ : CascadeMux
    port map (
            O => \N__26043\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14_cascade_\
        );

    \I__3807\ : InMux
    port map (
            O => \N__26040\,
            I => \N__26037\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__26037\,
            I => \N__26034\
        );

    \I__3805\ : Odrv4
    port map (
            O => \N__26034\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0\
        );

    \I__3804\ : CascadeMux
    port map (
            O => \N__26031\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_\
        );

    \I__3803\ : CascadeMux
    port map (
            O => \N__26028\,
            I => \N__26025\
        );

    \I__3802\ : InMux
    port map (
            O => \N__26025\,
            I => \N__26021\
        );

    \I__3801\ : InMux
    port map (
            O => \N__26024\,
            I => \N__26017\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__26021\,
            I => \N__26014\
        );

    \I__3799\ : InMux
    port map (
            O => \N__26020\,
            I => \N__26009\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__26017\,
            I => \N__26006\
        );

    \I__3797\ : Span4Mux_h
    port map (
            O => \N__26014\,
            I => \N__26003\
        );

    \I__3796\ : InMux
    port map (
            O => \N__26013\,
            I => \N__25998\
        );

    \I__3795\ : InMux
    port map (
            O => \N__26012\,
            I => \N__25998\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__26009\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3793\ : Odrv4
    port map (
            O => \N__26006\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3792\ : Odrv4
    port map (
            O => \N__26003\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__25998\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3790\ : InMux
    port map (
            O => \N__25989\,
            I => \N__25986\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__25986\,
            I => \current_shift_inst.PI_CTRL.N_71\
        );

    \I__3788\ : IoInMux
    port map (
            O => \N__25983\,
            I => \N__25980\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__25980\,
            I => \N__25977\
        );

    \I__3786\ : Span4Mux_s3_v
    port map (
            O => \N__25977\,
            I => \N__25974\
        );

    \I__3785\ : Span4Mux_h
    port map (
            O => \N__25974\,
            I => \N__25971\
        );

    \I__3784\ : Sp12to4
    port map (
            O => \N__25971\,
            I => \N__25968\
        );

    \I__3783\ : Span12Mux_s11_v
    port map (
            O => \N__25968\,
            I => \N__25965\
        );

    \I__3782\ : Span12Mux_v
    port map (
            O => \N__25965\,
            I => \N__25962\
        );

    \I__3781\ : Odrv12
    port map (
            O => \N__25962\,
            I => \pll_inst.red_c_i\
        );

    \I__3780\ : InMux
    port map (
            O => \N__25959\,
            I => \N__25956\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__25956\,
            I => \N__25953\
        );

    \I__3778\ : Span4Mux_v
    port map (
            O => \N__25953\,
            I => \N__25950\
        );

    \I__3777\ : Odrv4
    port map (
            O => \N__25950\,
            I => \current_shift_inst.PI_CTRL.integrator_i_20\
        );

    \I__3776\ : InMux
    port map (
            O => \N__25947\,
            I => \N__25944\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__25944\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt18\
        );

    \I__3774\ : InMux
    port map (
            O => \N__25941\,
            I => \N__25937\
        );

    \I__3773\ : InMux
    port map (
            O => \N__25940\,
            I => \N__25934\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__25937\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__25934\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__3770\ : InMux
    port map (
            O => \N__25929\,
            I => \N__25925\
        );

    \I__3769\ : InMux
    port map (
            O => \N__25928\,
            I => \N__25922\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__25925\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__25922\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__3766\ : InMux
    port map (
            O => \N__25917\,
            I => \N__25914\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__25914\,
            I => \phase_controller_inst1.stoper_hc.un4_running_df24\
        );

    \I__3764\ : CascadeMux
    port map (
            O => \N__25911\,
            I => \N__25908\
        );

    \I__3763\ : InMux
    port map (
            O => \N__25908\,
            I => \N__25905\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__25905\,
            I => \N__25902\
        );

    \I__3761\ : Span4Mux_v
    port map (
            O => \N__25902\,
            I => \N__25899\
        );

    \I__3760\ : Odrv4
    port map (
            O => \N__25899\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt16\
        );

    \I__3759\ : InMux
    port map (
            O => \N__25896\,
            I => \N__25891\
        );

    \I__3758\ : InMux
    port map (
            O => \N__25895\,
            I => \N__25886\
        );

    \I__3757\ : InMux
    port map (
            O => \N__25894\,
            I => \N__25886\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__25891\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__25886\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__3754\ : CascadeMux
    port map (
            O => \N__25881\,
            I => \N__25877\
        );

    \I__3753\ : InMux
    port map (
            O => \N__25880\,
            I => \N__25873\
        );

    \I__3752\ : InMux
    port map (
            O => \N__25877\,
            I => \N__25868\
        );

    \I__3751\ : InMux
    port map (
            O => \N__25876\,
            I => \N__25868\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__25873\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__25868\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__3748\ : CascadeMux
    port map (
            O => \N__25863\,
            I => \N__25860\
        );

    \I__3747\ : InMux
    port map (
            O => \N__25860\,
            I => \N__25857\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__25857\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\
        );

    \I__3745\ : InMux
    port map (
            O => \N__25854\,
            I => \N__25850\
        );

    \I__3744\ : InMux
    port map (
            O => \N__25853\,
            I => \N__25847\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__25850\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__25847\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__3741\ : InMux
    port map (
            O => \N__25842\,
            I => \N__25838\
        );

    \I__3740\ : InMux
    port map (
            O => \N__25841\,
            I => \N__25835\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__25838\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__25835\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__3737\ : InMux
    port map (
            O => \N__25830\,
            I => \N__25827\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__25827\,
            I => \phase_controller_inst1.stoper_hc.un4_running_df20\
        );

    \I__3735\ : InMux
    port map (
            O => \N__25824\,
            I => \N__25819\
        );

    \I__3734\ : InMux
    port map (
            O => \N__25823\,
            I => \N__25814\
        );

    \I__3733\ : InMux
    port map (
            O => \N__25822\,
            I => \N__25814\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__25819\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__25814\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__3730\ : CascadeMux
    port map (
            O => \N__25809\,
            I => \N__25805\
        );

    \I__3729\ : InMux
    port map (
            O => \N__25808\,
            I => \N__25800\
        );

    \I__3728\ : InMux
    port map (
            O => \N__25805\,
            I => \N__25800\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__25800\,
            I => \N__25797\
        );

    \I__3726\ : Span4Mux_v
    port map (
            O => \N__25797\,
            I => \N__25794\
        );

    \I__3725\ : Odrv4
    port map (
            O => \N__25794\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__3724\ : InMux
    port map (
            O => \N__25791\,
            I => \N__25786\
        );

    \I__3723\ : InMux
    port map (
            O => \N__25790\,
            I => \N__25781\
        );

    \I__3722\ : InMux
    port map (
            O => \N__25789\,
            I => \N__25781\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__25786\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__25781\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__3719\ : InMux
    port map (
            O => \N__25776\,
            I => \N__25773\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__25773\,
            I => \N__25770\
        );

    \I__3717\ : Odrv12
    port map (
            O => \N__25770\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\
        );

    \I__3716\ : InMux
    port map (
            O => \N__25767\,
            I => \N__25763\
        );

    \I__3715\ : InMux
    port map (
            O => \N__25766\,
            I => \N__25760\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__25763\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__25760\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__3712\ : InMux
    port map (
            O => \N__25755\,
            I => \N__25751\
        );

    \I__3711\ : InMux
    port map (
            O => \N__25754\,
            I => \N__25748\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__25751\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__25748\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__3708\ : InMux
    port map (
            O => \N__25743\,
            I => \N__25740\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__25740\,
            I => \phase_controller_inst1.stoper_hc.un4_running_df22\
        );

    \I__3706\ : InMux
    port map (
            O => \N__25737\,
            I => \N__25733\
        );

    \I__3705\ : InMux
    port map (
            O => \N__25736\,
            I => \N__25730\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__25733\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__25730\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__3702\ : InMux
    port map (
            O => \N__25725\,
            I => \N__25721\
        );

    \I__3701\ : InMux
    port map (
            O => \N__25724\,
            I => \N__25718\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__25721\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__25718\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__3698\ : InMux
    port map (
            O => \N__25713\,
            I => \N__25710\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__25710\,
            I => \N__25707\
        );

    \I__3696\ : Odrv4
    port map (
            O => \N__25707\,
            I => \phase_controller_inst1.stoper_hc.un4_running_df26\
        );

    \I__3695\ : InMux
    port map (
            O => \N__25704\,
            I => \N__25701\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__25701\,
            I => \N__25698\
        );

    \I__3693\ : Odrv4
    port map (
            O => \N__25698\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO\
        );

    \I__3692\ : InMux
    port map (
            O => \N__25695\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_28\
        );

    \I__3691\ : InMux
    port map (
            O => \N__25692\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30\
        );

    \I__3690\ : InMux
    port map (
            O => \N__25689\,
            I => \N__25685\
        );

    \I__3689\ : InMux
    port map (
            O => \N__25688\,
            I => \N__25682\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__25685\,
            I => \N__25679\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__25682\,
            I => \N__25676\
        );

    \I__3686\ : Span4Mux_v
    port map (
            O => \N__25679\,
            I => \N__25671\
        );

    \I__3685\ : Span4Mux_h
    port map (
            O => \N__25676\,
            I => \N__25671\
        );

    \I__3684\ : Odrv4
    port map (
            O => \N__25671\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__3683\ : CascadeMux
    port map (
            O => \N__25668\,
            I => \N__25665\
        );

    \I__3682\ : InMux
    port map (
            O => \N__25665\,
            I => \N__25660\
        );

    \I__3681\ : InMux
    port map (
            O => \N__25664\,
            I => \N__25656\
        );

    \I__3680\ : InMux
    port map (
            O => \N__25663\,
            I => \N__25653\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__25660\,
            I => \N__25650\
        );

    \I__3678\ : InMux
    port map (
            O => \N__25659\,
            I => \N__25647\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__25656\,
            I => \N__25644\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__25653\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__3675\ : Odrv4
    port map (
            O => \N__25650\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__25647\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__3673\ : Odrv12
    port map (
            O => \N__25644\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__3672\ : CascadeMux
    port map (
            O => \N__25635\,
            I => \N__25632\
        );

    \I__3671\ : InMux
    port map (
            O => \N__25632\,
            I => \N__25627\
        );

    \I__3670\ : InMux
    port map (
            O => \N__25631\,
            I => \N__25624\
        );

    \I__3669\ : InMux
    port map (
            O => \N__25630\,
            I => \N__25621\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__25627\,
            I => \N__25618\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__25624\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__25621\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__3665\ : Odrv12
    port map (
            O => \N__25618\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__3664\ : InMux
    port map (
            O => \N__25611\,
            I => \N__25608\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__25608\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\
        );

    \I__3662\ : InMux
    port map (
            O => \N__25605\,
            I => \N__25601\
        );

    \I__3661\ : InMux
    port map (
            O => \N__25604\,
            I => \N__25598\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__25601\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__25598\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__3658\ : CascadeMux
    port map (
            O => \N__25593\,
            I => \N__25590\
        );

    \I__3657\ : InMux
    port map (
            O => \N__25590\,
            I => \N__25587\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__25587\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__3655\ : CascadeMux
    port map (
            O => \N__25584\,
            I => \N__25581\
        );

    \I__3654\ : InMux
    port map (
            O => \N__25581\,
            I => \N__25578\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__25578\,
            I => \N__25575\
        );

    \I__3652\ : Odrv4
    port map (
            O => \N__25575\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\
        );

    \I__3651\ : InMux
    port map (
            O => \N__25572\,
            I => \N__25568\
        );

    \I__3650\ : InMux
    port map (
            O => \N__25571\,
            I => \N__25565\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__25568\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__25565\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__3647\ : InMux
    port map (
            O => \N__25560\,
            I => \N__25557\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__25557\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__3645\ : CascadeMux
    port map (
            O => \N__25554\,
            I => \N__25551\
        );

    \I__3644\ : InMux
    port map (
            O => \N__25551\,
            I => \N__25548\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__25548\,
            I => \N__25545\
        );

    \I__3642\ : Odrv4
    port map (
            O => \N__25545\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\
        );

    \I__3641\ : InMux
    port map (
            O => \N__25542\,
            I => \N__25538\
        );

    \I__3640\ : InMux
    port map (
            O => \N__25541\,
            I => \N__25535\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__25538\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__25535\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__3637\ : InMux
    port map (
            O => \N__25530\,
            I => \N__25527\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__25527\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__3635\ : InMux
    port map (
            O => \N__25524\,
            I => \N__25521\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__25521\,
            I => \N__25518\
        );

    \I__3633\ : Odrv4
    port map (
            O => \N__25518\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\
        );

    \I__3632\ : InMux
    port map (
            O => \N__25515\,
            I => \N__25511\
        );

    \I__3631\ : InMux
    port map (
            O => \N__25514\,
            I => \N__25508\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__25511\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__25508\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__3628\ : CascadeMux
    port map (
            O => \N__25503\,
            I => \N__25500\
        );

    \I__3627\ : InMux
    port map (
            O => \N__25500\,
            I => \N__25497\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__25497\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__3625\ : InMux
    port map (
            O => \N__25494\,
            I => \N__25491\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__25491\,
            I => \N__25488\
        );

    \I__3623\ : Odrv4
    port map (
            O => \N__25488\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\
        );

    \I__3622\ : InMux
    port map (
            O => \N__25485\,
            I => \N__25481\
        );

    \I__3621\ : InMux
    port map (
            O => \N__25484\,
            I => \N__25478\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__25481\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__25478\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__3618\ : CascadeMux
    port map (
            O => \N__25473\,
            I => \N__25470\
        );

    \I__3617\ : InMux
    port map (
            O => \N__25470\,
            I => \N__25467\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__25467\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__3615\ : CascadeMux
    port map (
            O => \N__25464\,
            I => \N__25461\
        );

    \I__3614\ : InMux
    port map (
            O => \N__25461\,
            I => \N__25458\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__25458\,
            I => \N__25455\
        );

    \I__3612\ : Odrv12
    port map (
            O => \N__25455\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\
        );

    \I__3611\ : InMux
    port map (
            O => \N__25452\,
            I => \N__25448\
        );

    \I__3610\ : InMux
    port map (
            O => \N__25451\,
            I => \N__25445\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__25448\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__25445\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__3607\ : InMux
    port map (
            O => \N__25440\,
            I => \N__25437\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__25437\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__3605\ : InMux
    port map (
            O => \N__25434\,
            I => \N__25431\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__25431\,
            I => \N__25428\
        );

    \I__3603\ : Odrv12
    port map (
            O => \N__25428\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\
        );

    \I__3602\ : CascadeMux
    port map (
            O => \N__25425\,
            I => \N__25422\
        );

    \I__3601\ : InMux
    port map (
            O => \N__25422\,
            I => \N__25418\
        );

    \I__3600\ : InMux
    port map (
            O => \N__25421\,
            I => \N__25415\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__25418\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__25415\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__3597\ : CascadeMux
    port map (
            O => \N__25410\,
            I => \N__25407\
        );

    \I__3596\ : InMux
    port map (
            O => \N__25407\,
            I => \N__25404\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__25404\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__3594\ : InMux
    port map (
            O => \N__25401\,
            I => \N__25398\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__25398\,
            I => \N__25395\
        );

    \I__3592\ : Span12Mux_s9_v
    port map (
            O => \N__25395\,
            I => \N__25392\
        );

    \I__3591\ : Odrv12
    port map (
            O => \N__25392\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\
        );

    \I__3590\ : InMux
    port map (
            O => \N__25389\,
            I => \N__25385\
        );

    \I__3589\ : InMux
    port map (
            O => \N__25388\,
            I => \N__25382\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__25385\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__25382\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__3586\ : CascadeMux
    port map (
            O => \N__25377\,
            I => \N__25374\
        );

    \I__3585\ : InMux
    port map (
            O => \N__25374\,
            I => \N__25371\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__25371\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__3583\ : InMux
    port map (
            O => \N__25368\,
            I => \N__25364\
        );

    \I__3582\ : InMux
    port map (
            O => \N__25367\,
            I => \N__25361\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__25364\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__25361\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__3579\ : InMux
    port map (
            O => \N__25356\,
            I => \N__25353\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__25353\,
            I => \N__25350\
        );

    \I__3577\ : Odrv12
    port map (
            O => \N__25350\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\
        );

    \I__3576\ : CascadeMux
    port map (
            O => \N__25347\,
            I => \N__25344\
        );

    \I__3575\ : InMux
    port map (
            O => \N__25344\,
            I => \N__25341\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__25341\,
            I => \N__25338\
        );

    \I__3573\ : Odrv4
    port map (
            O => \N__25338\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__3572\ : InMux
    port map (
            O => \N__25335\,
            I => \N__25332\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__25332\,
            I => \N__25329\
        );

    \I__3570\ : Span4Mux_v
    port map (
            O => \N__25329\,
            I => \N__25326\
        );

    \I__3569\ : Span4Mux_v
    port map (
            O => \N__25326\,
            I => \N__25323\
        );

    \I__3568\ : Odrv4
    port map (
            O => \N__25323\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\
        );

    \I__3567\ : InMux
    port map (
            O => \N__25320\,
            I => \N__25316\
        );

    \I__3566\ : InMux
    port map (
            O => \N__25319\,
            I => \N__25313\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__25316\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__25313\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__3563\ : CascadeMux
    port map (
            O => \N__25308\,
            I => \N__25305\
        );

    \I__3562\ : InMux
    port map (
            O => \N__25305\,
            I => \N__25302\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__25302\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__3560\ : InMux
    port map (
            O => \N__25299\,
            I => \N__25296\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__25296\,
            I => \N__25293\
        );

    \I__3558\ : Span4Mux_v
    port map (
            O => \N__25293\,
            I => \N__25290\
        );

    \I__3557\ : Span4Mux_h
    port map (
            O => \N__25290\,
            I => \N__25287\
        );

    \I__3556\ : Odrv4
    port map (
            O => \N__25287\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\
        );

    \I__3555\ : InMux
    port map (
            O => \N__25284\,
            I => \N__25280\
        );

    \I__3554\ : InMux
    port map (
            O => \N__25283\,
            I => \N__25277\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__25280\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__25277\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3551\ : CascadeMux
    port map (
            O => \N__25272\,
            I => \N__25269\
        );

    \I__3550\ : InMux
    port map (
            O => \N__25269\,
            I => \N__25266\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__25266\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__3548\ : InMux
    port map (
            O => \N__25263\,
            I => \N__25259\
        );

    \I__3547\ : InMux
    port map (
            O => \N__25262\,
            I => \N__25256\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__25259\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__25256\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__3544\ : CascadeMux
    port map (
            O => \N__25251\,
            I => \N__25248\
        );

    \I__3543\ : InMux
    port map (
            O => \N__25248\,
            I => \N__25245\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__25245\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__3541\ : InMux
    port map (
            O => \N__25242\,
            I => \N__25239\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__25239\,
            I => \N__25236\
        );

    \I__3539\ : Odrv4
    port map (
            O => \N__25236\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\
        );

    \I__3538\ : InMux
    port map (
            O => \N__25233\,
            I => \N__25229\
        );

    \I__3537\ : InMux
    port map (
            O => \N__25232\,
            I => \N__25226\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__25229\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__25226\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__3534\ : CascadeMux
    port map (
            O => \N__25221\,
            I => \N__25218\
        );

    \I__3533\ : InMux
    port map (
            O => \N__25218\,
            I => \N__25215\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__25215\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__3531\ : CascadeMux
    port map (
            O => \N__25212\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9_cascade_\
        );

    \I__3530\ : InMux
    port map (
            O => \N__25209\,
            I => \N__25206\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__25206\,
            I => \phase_controller_inst1.stoper_hc.N_267_iZ0Z_1\
        );

    \I__3528\ : CascadeMux
    port map (
            O => \N__25203\,
            I => \N__25198\
        );

    \I__3527\ : InMux
    port map (
            O => \N__25202\,
            I => \N__25195\
        );

    \I__3526\ : InMux
    port map (
            O => \N__25201\,
            I => \N__25192\
        );

    \I__3525\ : InMux
    port map (
            O => \N__25198\,
            I => \N__25189\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__25195\,
            I => \N__25186\
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__25192\,
            I => \N__25183\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__25189\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__3521\ : Odrv4
    port map (
            O => \N__25186\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__3520\ : Odrv4
    port map (
            O => \N__25183\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__3519\ : InMux
    port map (
            O => \N__25176\,
            I => \N__25173\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__25173\,
            I => \N__25170\
        );

    \I__3517\ : Span4Mux_v
    port map (
            O => \N__25170\,
            I => \N__25167\
        );

    \I__3516\ : Odrv4
    port map (
            O => \N__25167\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\
        );

    \I__3515\ : CascadeMux
    port map (
            O => \N__25164\,
            I => \N__25161\
        );

    \I__3514\ : InMux
    port map (
            O => \N__25161\,
            I => \N__25158\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__25158\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__3512\ : InMux
    port map (
            O => \N__25155\,
            I => \N__25151\
        );

    \I__3511\ : InMux
    port map (
            O => \N__25154\,
            I => \N__25148\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__25151\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__25148\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__3508\ : CascadeMux
    port map (
            O => \N__25143\,
            I => \N__25140\
        );

    \I__3507\ : InMux
    port map (
            O => \N__25140\,
            I => \N__25137\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__25137\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__3505\ : CascadeMux
    port map (
            O => \N__25134\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9_cascade_\
        );

    \I__3504\ : CascadeMux
    port map (
            O => \N__25131\,
            I => \delay_measurement_inst.delay_hc_timer.N_342_i_cascade_\
        );

    \I__3503\ : CascadeMux
    port map (
            O => \N__25128\,
            I => \elapsed_time_ns_1_RNIHHC6P1_0_18_cascade_\
        );

    \I__3502\ : InMux
    port map (
            O => \N__25125\,
            I => \N__25122\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__25122\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18\
        );

    \I__3500\ : InMux
    port map (
            O => \N__25119\,
            I => \N__25116\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__25116\,
            I => \N__25113\
        );

    \I__3498\ : Span4Mux_v
    port map (
            O => \N__25113\,
            I => \N__25110\
        );

    \I__3497\ : Odrv4
    port map (
            O => \N__25110\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17\
        );

    \I__3496\ : InMux
    port map (
            O => \N__25107\,
            I => \N__25101\
        );

    \I__3495\ : CascadeMux
    port map (
            O => \N__25106\,
            I => \N__25098\
        );

    \I__3494\ : InMux
    port map (
            O => \N__25105\,
            I => \N__25093\
        );

    \I__3493\ : InMux
    port map (
            O => \N__25104\,
            I => \N__25093\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__25101\,
            I => \N__25090\
        );

    \I__3491\ : InMux
    port map (
            O => \N__25098\,
            I => \N__25087\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__25093\,
            I => \N__25084\
        );

    \I__3489\ : Odrv4
    port map (
            O => \N__25090\,
            I => \elapsed_time_ns_1_RNIFFC6P1_0_16\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__25087\,
            I => \elapsed_time_ns_1_RNIFFC6P1_0_16\
        );

    \I__3487\ : Odrv12
    port map (
            O => \N__25084\,
            I => \elapsed_time_ns_1_RNIFFC6P1_0_16\
        );

    \I__3486\ : CascadeMux
    port map (
            O => \N__25077\,
            I => \phase_controller_inst1.stoper_hc.N_267_iZ0Z_1_cascade_\
        );

    \I__3485\ : CascadeMux
    port map (
            O => \N__25074\,
            I => \elapsed_time_ns_1_RNIFFC6P1_0_16_cascade_\
        );

    \I__3484\ : InMux
    port map (
            O => \N__25071\,
            I => \N__25065\
        );

    \I__3483\ : InMux
    port map (
            O => \N__25070\,
            I => \N__25065\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__25065\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\
        );

    \I__3481\ : InMux
    port map (
            O => \N__25062\,
            I => \N__25056\
        );

    \I__3480\ : InMux
    port map (
            O => \N__25061\,
            I => \N__25056\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__25056\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\
        );

    \I__3478\ : CascadeMux
    port map (
            O => \N__25053\,
            I => \elapsed_time_ns_1_RNILGKEE1_0_4_cascade_\
        );

    \I__3477\ : CascadeMux
    port map (
            O => \N__25050\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2_cascade_\
        );

    \I__3476\ : CascadeMux
    port map (
            O => \N__25047\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6_cascade_\
        );

    \I__3475\ : CascadeMux
    port map (
            O => \N__25044\,
            I => \elapsed_time_ns_1_RNIUE3CP1_0_6_cascade_\
        );

    \I__3474\ : CascadeMux
    port map (
            O => \N__25041\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_\
        );

    \I__3473\ : InMux
    port map (
            O => \N__25038\,
            I => \N__25035\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__25035\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__3471\ : InMux
    port map (
            O => \N__25032\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\
        );

    \I__3470\ : CascadeMux
    port map (
            O => \N__25029\,
            I => \N__25026\
        );

    \I__3469\ : InMux
    port map (
            O => \N__25026\,
            I => \N__25023\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__25023\,
            I => \N__25020\
        );

    \I__3467\ : Odrv4
    port map (
            O => \N__25020\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__3466\ : InMux
    port map (
            O => \N__25017\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\
        );

    \I__3465\ : InMux
    port map (
            O => \N__25014\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\
        );

    \I__3464\ : InMux
    port map (
            O => \N__25011\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\
        );

    \I__3463\ : InMux
    port map (
            O => \N__25008\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\
        );

    \I__3462\ : InMux
    port map (
            O => \N__25005\,
            I => \bfn_9_13_0_\
        );

    \I__3461\ : CascadeMux
    port map (
            O => \N__25002\,
            I => \N__24999\
        );

    \I__3460\ : InMux
    port map (
            O => \N__24999\,
            I => \N__24996\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__24996\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\
        );

    \I__3458\ : InMux
    port map (
            O => \N__24993\,
            I => \N__24990\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__24990\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3\
        );

    \I__3456\ : InMux
    port map (
            O => \N__24987\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\
        );

    \I__3455\ : InMux
    port map (
            O => \N__24984\,
            I => \N__24981\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__24981\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__3453\ : InMux
    port map (
            O => \N__24978\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\
        );

    \I__3452\ : InMux
    port map (
            O => \N__24975\,
            I => \N__24972\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__24972\,
            I => \N__24969\
        );

    \I__3450\ : Odrv4
    port map (
            O => \N__24969\,
            I => \current_shift_inst.PI_CTRL.integrator_i_19\
        );

    \I__3449\ : CascadeMux
    port map (
            O => \N__24966\,
            I => \N__24963\
        );

    \I__3448\ : InMux
    port map (
            O => \N__24963\,
            I => \N__24960\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__24960\,
            I => \N__24957\
        );

    \I__3446\ : Odrv12
    port map (
            O => \N__24957\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__3445\ : InMux
    port map (
            O => \N__24954\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\
        );

    \I__3444\ : CascadeMux
    port map (
            O => \N__24951\,
            I => \N__24948\
        );

    \I__3443\ : InMux
    port map (
            O => \N__24948\,
            I => \N__24945\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__24945\,
            I => \N__24942\
        );

    \I__3441\ : Odrv4
    port map (
            O => \N__24942\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__3440\ : InMux
    port map (
            O => \N__24939\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\
        );

    \I__3439\ : CascadeMux
    port map (
            O => \N__24936\,
            I => \N__24933\
        );

    \I__3438\ : InMux
    port map (
            O => \N__24933\,
            I => \N__24930\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__24930\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__3436\ : InMux
    port map (
            O => \N__24927\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\
        );

    \I__3435\ : InMux
    port map (
            O => \N__24924\,
            I => \N__24921\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__24921\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__3433\ : InMux
    port map (
            O => \N__24918\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\
        );

    \I__3432\ : InMux
    port map (
            O => \N__24915\,
            I => \N__24912\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__24912\,
            I => \N__24909\
        );

    \I__3430\ : Span4Mux_v
    port map (
            O => \N__24909\,
            I => \N__24906\
        );

    \I__3429\ : Span4Mux_v
    port map (
            O => \N__24906\,
            I => \N__24903\
        );

    \I__3428\ : Odrv4
    port map (
            O => \N__24903\,
            I => \current_shift_inst.PI_CTRL.integrator_i_23\
        );

    \I__3427\ : InMux
    port map (
            O => \N__24900\,
            I => \N__24897\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__24897\,
            I => \N__24894\
        );

    \I__3425\ : Odrv4
    port map (
            O => \N__24894\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__3424\ : InMux
    port map (
            O => \N__24891\,
            I => \bfn_9_12_0_\
        );

    \I__3423\ : InMux
    port map (
            O => \N__24888\,
            I => \N__24885\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__24885\,
            I => \N__24882\
        );

    \I__3421\ : Odrv4
    port map (
            O => \N__24882\,
            I => \current_shift_inst.PI_CTRL.integrator_i_24\
        );

    \I__3420\ : CascadeMux
    port map (
            O => \N__24879\,
            I => \N__24876\
        );

    \I__3419\ : InMux
    port map (
            O => \N__24876\,
            I => \N__24873\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__24873\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__3417\ : InMux
    port map (
            O => \N__24870\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\
        );

    \I__3416\ : CascadeMux
    port map (
            O => \N__24867\,
            I => \N__24864\
        );

    \I__3415\ : InMux
    port map (
            O => \N__24864\,
            I => \N__24861\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__24861\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__3413\ : InMux
    port map (
            O => \N__24858\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\
        );

    \I__3412\ : CascadeMux
    port map (
            O => \N__24855\,
            I => \N__24852\
        );

    \I__3411\ : InMux
    port map (
            O => \N__24852\,
            I => \N__24849\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__24849\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__3409\ : InMux
    port map (
            O => \N__24846\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\
        );

    \I__3408\ : InMux
    port map (
            O => \N__24843\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\
        );

    \I__3407\ : CascadeMux
    port map (
            O => \N__24840\,
            I => \N__24837\
        );

    \I__3406\ : InMux
    port map (
            O => \N__24837\,
            I => \N__24834\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__24834\,
            I => \N__24831\
        );

    \I__3404\ : Odrv4
    port map (
            O => \N__24831\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__3403\ : InMux
    port map (
            O => \N__24828\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\
        );

    \I__3402\ : InMux
    port map (
            O => \N__24825\,
            I => \N__24822\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__24822\,
            I => \N__24819\
        );

    \I__3400\ : Odrv4
    port map (
            O => \N__24819\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__3399\ : InMux
    port map (
            O => \N__24816\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\
        );

    \I__3398\ : CascadeMux
    port map (
            O => \N__24813\,
            I => \N__24810\
        );

    \I__3397\ : InMux
    port map (
            O => \N__24810\,
            I => \N__24807\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__24807\,
            I => \N__24804\
        );

    \I__3395\ : Odrv4
    port map (
            O => \N__24804\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__3394\ : InMux
    port map (
            O => \N__24801\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\
        );

    \I__3393\ : InMux
    port map (
            O => \N__24798\,
            I => \N__24795\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__24795\,
            I => \N__24792\
        );

    \I__3391\ : Odrv4
    port map (
            O => \N__24792\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__3390\ : InMux
    port map (
            O => \N__24789\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\
        );

    \I__3389\ : InMux
    port map (
            O => \N__24786\,
            I => \N__24783\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__24783\,
            I => \N__24780\
        );

    \I__3387\ : Odrv12
    port map (
            O => \N__24780\,
            I => \current_shift_inst.PI_CTRL.integrator_i_15\
        );

    \I__3386\ : CascadeMux
    port map (
            O => \N__24777\,
            I => \N__24774\
        );

    \I__3385\ : InMux
    port map (
            O => \N__24774\,
            I => \N__24771\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__24771\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__3383\ : InMux
    port map (
            O => \N__24768\,
            I => \bfn_9_11_0_\
        );

    \I__3382\ : InMux
    port map (
            O => \N__24765\,
            I => \N__24762\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__24762\,
            I => \N__24759\
        );

    \I__3380\ : Odrv4
    port map (
            O => \N__24759\,
            I => \current_shift_inst.PI_CTRL.integrator_i_16\
        );

    \I__3379\ : CascadeMux
    port map (
            O => \N__24756\,
            I => \N__24753\
        );

    \I__3378\ : InMux
    port map (
            O => \N__24753\,
            I => \N__24750\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__24750\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6IZ0\
        );

    \I__3376\ : InMux
    port map (
            O => \N__24747\,
            I => \N__24744\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__24744\,
            I => \N__24741\
        );

    \I__3374\ : Span4Mux_v
    port map (
            O => \N__24741\,
            I => \N__24738\
        );

    \I__3373\ : Odrv4
    port map (
            O => \N__24738\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__3372\ : InMux
    port map (
            O => \N__24735\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\
        );

    \I__3371\ : CascadeMux
    port map (
            O => \N__24732\,
            I => \N__24729\
        );

    \I__3370\ : InMux
    port map (
            O => \N__24729\,
            I => \N__24726\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__24726\,
            I => \N__24723\
        );

    \I__3368\ : Span4Mux_v
    port map (
            O => \N__24723\,
            I => \N__24720\
        );

    \I__3367\ : Odrv4
    port map (
            O => \N__24720\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__3366\ : InMux
    port map (
            O => \N__24717\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\
        );

    \I__3365\ : InMux
    port map (
            O => \N__24714\,
            I => \N__24711\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__24711\,
            I => \N__24708\
        );

    \I__3363\ : Odrv4
    port map (
            O => \N__24708\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\
        );

    \I__3362\ : InMux
    port map (
            O => \N__24705\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\
        );

    \I__3361\ : InMux
    port map (
            O => \N__24702\,
            I => \N__24699\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__24699\,
            I => \current_shift_inst.PI_CTRL.integrator_i_3\
        );

    \I__3359\ : CascadeMux
    port map (
            O => \N__24696\,
            I => \N__24693\
        );

    \I__3358\ : InMux
    port map (
            O => \N__24693\,
            I => \N__24690\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__24690\,
            I => \current_shift_inst.PI_CTRL.error_control_RNID56UZ0Z_7\
        );

    \I__3356\ : InMux
    port map (
            O => \N__24687\,
            I => \N__24684\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__24684\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\
        );

    \I__3354\ : InMux
    port map (
            O => \N__24681\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\
        );

    \I__3353\ : InMux
    port map (
            O => \N__24678\,
            I => \N__24675\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__24675\,
            I => \N__24672\
        );

    \I__3351\ : Odrv12
    port map (
            O => \N__24672\,
            I => \current_shift_inst.PI_CTRL.integrator_i_4\
        );

    \I__3350\ : InMux
    port map (
            O => \N__24669\,
            I => \N__24666\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__24666\,
            I => \N__24663\
        );

    \I__3348\ : Odrv4
    port map (
            O => \N__24663\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__3347\ : InMux
    port map (
            O => \N__24660\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\
        );

    \I__3346\ : InMux
    port map (
            O => \N__24657\,
            I => \N__24654\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__24654\,
            I => \N__24651\
        );

    \I__3344\ : Span4Mux_h
    port map (
            O => \N__24651\,
            I => \N__24648\
        );

    \I__3343\ : Odrv4
    port map (
            O => \N__24648\,
            I => \current_shift_inst.PI_CTRL.integrator_i_5\
        );

    \I__3342\ : CascadeMux
    port map (
            O => \N__24645\,
            I => \N__24642\
        );

    \I__3341\ : InMux
    port map (
            O => \N__24642\,
            I => \N__24639\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__24639\,
            I => \N__24636\
        );

    \I__3339\ : Odrv4
    port map (
            O => \N__24636\,
            I => \current_shift_inst.PI_CTRL.error_control_RNILF8UZ0Z_9\
        );

    \I__3338\ : InMux
    port map (
            O => \N__24633\,
            I => \N__24630\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__24630\,
            I => \N__24627\
        );

    \I__3336\ : Odrv4
    port map (
            O => \N__24627\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__3335\ : InMux
    port map (
            O => \N__24624\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\
        );

    \I__3334\ : InMux
    port map (
            O => \N__24621\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\
        );

    \I__3333\ : InMux
    port map (
            O => \N__24618\,
            I => \N__24615\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__24615\,
            I => \current_shift_inst.PI_CTRL.integrator_i_7\
        );

    \I__3331\ : CascadeMux
    port map (
            O => \N__24612\,
            I => \N__24609\
        );

    \I__3330\ : InMux
    port map (
            O => \N__24609\,
            I => \N__24606\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__24606\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIISQ01Z0Z_11\
        );

    \I__3328\ : InMux
    port map (
            O => \N__24603\,
            I => \N__24600\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__24600\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__3326\ : InMux
    port map (
            O => \N__24597\,
            I => \bfn_9_10_0_\
        );

    \I__3325\ : InMux
    port map (
            O => \N__24594\,
            I => \N__24591\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__24591\,
            I => \current_shift_inst.PI_CTRL.integrator_i_8\
        );

    \I__3323\ : InMux
    port map (
            O => \N__24588\,
            I => \N__24585\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__24585\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__3321\ : InMux
    port map (
            O => \N__24582\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\
        );

    \I__3320\ : InMux
    port map (
            O => \N__24579\,
            I => \N__24576\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__24576\,
            I => \N__24573\
        );

    \I__3318\ : Odrv4
    port map (
            O => \N__24573\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0\
        );

    \I__3317\ : InMux
    port map (
            O => \N__24570\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\
        );

    \I__3316\ : InMux
    port map (
            O => \N__24567\,
            I => \N__24564\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__24564\,
            I => \N__24561\
        );

    \I__3314\ : Span4Mux_h
    port map (
            O => \N__24561\,
            I => \N__24555\
        );

    \I__3313\ : InMux
    port map (
            O => \N__24560\,
            I => \N__24552\
        );

    \I__3312\ : CascadeMux
    port map (
            O => \N__24559\,
            I => \N__24549\
        );

    \I__3311\ : CascadeMux
    port map (
            O => \N__24558\,
            I => \N__24546\
        );

    \I__3310\ : Sp12to4
    port map (
            O => \N__24555\,
            I => \N__24543\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__24552\,
            I => \N__24540\
        );

    \I__3308\ : InMux
    port map (
            O => \N__24549\,
            I => \N__24535\
        );

    \I__3307\ : InMux
    port map (
            O => \N__24546\,
            I => \N__24535\
        );

    \I__3306\ : Span12Mux_s10_v
    port map (
            O => \N__24543\,
            I => \N__24532\
        );

    \I__3305\ : Span4Mux_h
    port map (
            O => \N__24540\,
            I => \N__24529\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__24535\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__3303\ : Odrv12
    port map (
            O => \N__24532\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__3302\ : Odrv4
    port map (
            O => \N__24529\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__3301\ : IoInMux
    port map (
            O => \N__24522\,
            I => \N__24519\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__24519\,
            I => s3_phy_c
        );

    \I__3299\ : InMux
    port map (
            O => \N__24516\,
            I => \N__24513\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__24513\,
            I => \N__24510\
        );

    \I__3297\ : Odrv12
    port map (
            O => \N__24510\,
            I => il_min_comp1_c
        );

    \I__3296\ : InMux
    port map (
            O => \N__24507\,
            I => \N__24504\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__24504\,
            I => \N__24500\
        );

    \I__3294\ : InMux
    port map (
            O => \N__24503\,
            I => \N__24497\
        );

    \I__3293\ : Span4Mux_h
    port map (
            O => \N__24500\,
            I => \N__24490\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__24497\,
            I => \N__24490\
        );

    \I__3291\ : InMux
    port map (
            O => \N__24496\,
            I => \N__24487\
        );

    \I__3290\ : InMux
    port map (
            O => \N__24495\,
            I => \N__24484\
        );

    \I__3289\ : Span4Mux_v
    port map (
            O => \N__24490\,
            I => \N__24481\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__24487\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__24484\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__3286\ : Odrv4
    port map (
            O => \N__24481\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__3285\ : ClkMux
    port map (
            O => \N__24474\,
            I => \N__24468\
        );

    \I__3284\ : ClkMux
    port map (
            O => \N__24473\,
            I => \N__24468\
        );

    \I__3283\ : GlobalMux
    port map (
            O => \N__24468\,
            I => \N__24465\
        );

    \I__3282\ : gio2CtrlBuf
    port map (
            O => \N__24465\,
            I => delay_hc_input_c_g
        );

    \I__3281\ : InMux
    port map (
            O => \N__24462\,
            I => \N__24459\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__24459\,
            I => \N__24456\
        );

    \I__3279\ : Span4Mux_v
    port map (
            O => \N__24456\,
            I => \N__24453\
        );

    \I__3278\ : Span4Mux_h
    port map (
            O => \N__24453\,
            I => \N__24450\
        );

    \I__3277\ : Odrv4
    port map (
            O => \N__24450\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__3276\ : InMux
    port map (
            O => \N__24447\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\
        );

    \I__3275\ : InMux
    port map (
            O => \N__24444\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\
        );

    \I__3274\ : InMux
    port map (
            O => \N__24441\,
            I => \bfn_8_26_0_\
        );

    \I__3273\ : InMux
    port map (
            O => \N__24438\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\
        );

    \I__3272\ : InMux
    port map (
            O => \N__24435\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\
        );

    \I__3271\ : InMux
    port map (
            O => \N__24432\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\
        );

    \I__3270\ : InMux
    port map (
            O => \N__24429\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\
        );

    \I__3269\ : InMux
    port map (
            O => \N__24426\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\
        );

    \I__3268\ : InMux
    port map (
            O => \N__24423\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\
        );

    \I__3267\ : InMux
    port map (
            O => \N__24420\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__3266\ : InMux
    port map (
            O => \N__24417\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__3265\ : InMux
    port map (
            O => \N__24414\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__3264\ : InMux
    port map (
            O => \N__24411\,
            I => \bfn_8_25_0_\
        );

    \I__3263\ : InMux
    port map (
            O => \N__24408\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__3262\ : InMux
    port map (
            O => \N__24405\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__3261\ : InMux
    port map (
            O => \N__24402\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\
        );

    \I__3260\ : InMux
    port map (
            O => \N__24399\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__3259\ : InMux
    port map (
            O => \N__24396\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\
        );

    \I__3258\ : InMux
    port map (
            O => \N__24393\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__3257\ : InMux
    port map (
            O => \N__24390\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__3256\ : InMux
    port map (
            O => \N__24387\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__3255\ : InMux
    port map (
            O => \N__24384\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__3254\ : InMux
    port map (
            O => \N__24381\,
            I => \bfn_8_24_0_\
        );

    \I__3253\ : InMux
    port map (
            O => \N__24378\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__3252\ : InMux
    port map (
            O => \N__24375\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__3251\ : InMux
    port map (
            O => \N__24372\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__3250\ : InMux
    port map (
            O => \N__24369\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__3249\ : CascadeMux
    port map (
            O => \N__24366\,
            I => \N__24363\
        );

    \I__3248\ : InMux
    port map (
            O => \N__24363\,
            I => \N__24359\
        );

    \I__3247\ : InMux
    port map (
            O => \N__24362\,
            I => \N__24356\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__24359\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__24356\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__3244\ : InMux
    port map (
            O => \N__24351\,
            I => \N__24347\
        );

    \I__3243\ : InMux
    port map (
            O => \N__24350\,
            I => \N__24344\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__24347\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__24344\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\
        );

    \I__3240\ : InMux
    port map (
            O => \N__24339\,
            I => \N__24336\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__24336\,
            I => \N__24329\
        );

    \I__3238\ : InMux
    port map (
            O => \N__24335\,
            I => \N__24324\
        );

    \I__3237\ : InMux
    port map (
            O => \N__24334\,
            I => \N__24324\
        );

    \I__3236\ : InMux
    port map (
            O => \N__24333\,
            I => \N__24319\
        );

    \I__3235\ : InMux
    port map (
            O => \N__24332\,
            I => \N__24319\
        );

    \I__3234\ : Odrv4
    port map (
            O => \N__24329\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__24324\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__24319\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__3231\ : CascadeMux
    port map (
            O => \N__24312\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\
        );

    \I__3230\ : CascadeMux
    port map (
            O => \N__24309\,
            I => \N__24306\
        );

    \I__3229\ : InMux
    port map (
            O => \N__24306\,
            I => \N__24303\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__24303\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\
        );

    \I__3227\ : InMux
    port map (
            O => \N__24300\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__3226\ : InMux
    port map (
            O => \N__24297\,
            I => \N__24294\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__24294\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIM9HS1Z0Z_28\
        );

    \I__3224\ : InMux
    port map (
            O => \N__24291\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__3223\ : InMux
    port map (
            O => \N__24288\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__3222\ : InMux
    port map (
            O => \N__24285\,
            I => \bfn_8_18_0_\
        );

    \I__3221\ : InMux
    port map (
            O => \N__24282\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__3220\ : InMux
    port map (
            O => \N__24279\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__3219\ : InMux
    port map (
            O => \N__24276\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__3218\ : InMux
    port map (
            O => \N__24273\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__3217\ : InMux
    port map (
            O => \N__24270\,
            I => \N__24232\
        );

    \I__3216\ : InMux
    port map (
            O => \N__24269\,
            I => \N__24232\
        );

    \I__3215\ : InMux
    port map (
            O => \N__24268\,
            I => \N__24232\
        );

    \I__3214\ : InMux
    port map (
            O => \N__24267\,
            I => \N__24232\
        );

    \I__3213\ : InMux
    port map (
            O => \N__24266\,
            I => \N__24223\
        );

    \I__3212\ : InMux
    port map (
            O => \N__24265\,
            I => \N__24223\
        );

    \I__3211\ : InMux
    port map (
            O => \N__24264\,
            I => \N__24223\
        );

    \I__3210\ : InMux
    port map (
            O => \N__24263\,
            I => \N__24223\
        );

    \I__3209\ : InMux
    port map (
            O => \N__24262\,
            I => \N__24218\
        );

    \I__3208\ : InMux
    port map (
            O => \N__24261\,
            I => \N__24218\
        );

    \I__3207\ : InMux
    port map (
            O => \N__24260\,
            I => \N__24209\
        );

    \I__3206\ : InMux
    port map (
            O => \N__24259\,
            I => \N__24209\
        );

    \I__3205\ : InMux
    port map (
            O => \N__24258\,
            I => \N__24209\
        );

    \I__3204\ : InMux
    port map (
            O => \N__24257\,
            I => \N__24209\
        );

    \I__3203\ : InMux
    port map (
            O => \N__24256\,
            I => \N__24200\
        );

    \I__3202\ : InMux
    port map (
            O => \N__24255\,
            I => \N__24200\
        );

    \I__3201\ : InMux
    port map (
            O => \N__24254\,
            I => \N__24200\
        );

    \I__3200\ : InMux
    port map (
            O => \N__24253\,
            I => \N__24200\
        );

    \I__3199\ : InMux
    port map (
            O => \N__24252\,
            I => \N__24191\
        );

    \I__3198\ : InMux
    port map (
            O => \N__24251\,
            I => \N__24191\
        );

    \I__3197\ : InMux
    port map (
            O => \N__24250\,
            I => \N__24191\
        );

    \I__3196\ : InMux
    port map (
            O => \N__24249\,
            I => \N__24191\
        );

    \I__3195\ : InMux
    port map (
            O => \N__24248\,
            I => \N__24182\
        );

    \I__3194\ : InMux
    port map (
            O => \N__24247\,
            I => \N__24182\
        );

    \I__3193\ : InMux
    port map (
            O => \N__24246\,
            I => \N__24182\
        );

    \I__3192\ : InMux
    port map (
            O => \N__24245\,
            I => \N__24182\
        );

    \I__3191\ : InMux
    port map (
            O => \N__24244\,
            I => \N__24173\
        );

    \I__3190\ : InMux
    port map (
            O => \N__24243\,
            I => \N__24173\
        );

    \I__3189\ : InMux
    port map (
            O => \N__24242\,
            I => \N__24173\
        );

    \I__3188\ : InMux
    port map (
            O => \N__24241\,
            I => \N__24173\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__24232\,
            I => \N__24162\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__24223\,
            I => \N__24162\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__24218\,
            I => \N__24162\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__24209\,
            I => \N__24162\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__24200\,
            I => \N__24162\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__24191\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__24182\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__24173\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__3179\ : Odrv4
    port map (
            O => \N__24162\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__3178\ : InMux
    port map (
            O => \N__24153\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__3177\ : CEMux
    port map (
            O => \N__24150\,
            I => \N__24147\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__24147\,
            I => \N__24141\
        );

    \I__3175\ : CEMux
    port map (
            O => \N__24146\,
            I => \N__24138\
        );

    \I__3174\ : CEMux
    port map (
            O => \N__24145\,
            I => \N__24135\
        );

    \I__3173\ : CEMux
    port map (
            O => \N__24144\,
            I => \N__24132\
        );

    \I__3172\ : Span4Mux_v
    port map (
            O => \N__24141\,
            I => \N__24129\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__24138\,
            I => \N__24126\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__24135\,
            I => \N__24123\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__24132\,
            I => \N__24120\
        );

    \I__3168\ : Span4Mux_h
    port map (
            O => \N__24129\,
            I => \N__24113\
        );

    \I__3167\ : Span4Mux_v
    port map (
            O => \N__24126\,
            I => \N__24113\
        );

    \I__3166\ : Span4Mux_h
    port map (
            O => \N__24123\,
            I => \N__24113\
        );

    \I__3165\ : Odrv12
    port map (
            O => \N__24120\,
            I => \delay_measurement_inst.delay_hc_timer.N_394_i\
        );

    \I__3164\ : Odrv4
    port map (
            O => \N__24113\,
            I => \delay_measurement_inst.delay_hc_timer.N_394_i\
        );

    \I__3163\ : InMux
    port map (
            O => \N__24108\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__3162\ : InMux
    port map (
            O => \N__24105\,
            I => \bfn_8_17_0_\
        );

    \I__3161\ : InMux
    port map (
            O => \N__24102\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__3160\ : InMux
    port map (
            O => \N__24099\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__3159\ : InMux
    port map (
            O => \N__24096\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__3158\ : InMux
    port map (
            O => \N__24093\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__3157\ : InMux
    port map (
            O => \N__24090\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__3156\ : InMux
    port map (
            O => \N__24087\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__3155\ : InMux
    port map (
            O => \N__24084\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__3154\ : InMux
    port map (
            O => \N__24081\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__3153\ : InMux
    port map (
            O => \N__24078\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__3152\ : InMux
    port map (
            O => \N__24075\,
            I => \bfn_8_16_0_\
        );

    \I__3151\ : InMux
    port map (
            O => \N__24072\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__3150\ : InMux
    port map (
            O => \N__24069\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__3149\ : InMux
    port map (
            O => \N__24066\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__3148\ : InMux
    port map (
            O => \N__24063\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__3147\ : InMux
    port map (
            O => \N__24060\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__3146\ : InMux
    port map (
            O => \N__24057\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__3145\ : InMux
    port map (
            O => \N__24054\,
            I => \N__24046\
        );

    \I__3144\ : InMux
    port map (
            O => \N__24053\,
            I => \N__24046\
        );

    \I__3143\ : InMux
    port map (
            O => \N__24052\,
            I => \N__24043\
        );

    \I__3142\ : InMux
    port map (
            O => \N__24051\,
            I => \N__24040\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__24046\,
            I => \N__24037\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__24043\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__24040\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__3138\ : Odrv4
    port map (
            O => \N__24037\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__3137\ : InMux
    port map (
            O => \N__24030\,
            I => \N__24025\
        );

    \I__3136\ : InMux
    port map (
            O => \N__24029\,
            I => \N__24022\
        );

    \I__3135\ : InMux
    port map (
            O => \N__24028\,
            I => \N__24019\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__24025\,
            I => \N__24016\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__24022\,
            I => \N__24009\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__24019\,
            I => \N__24009\
        );

    \I__3131\ : Span4Mux_v
    port map (
            O => \N__24016\,
            I => \N__24009\
        );

    \I__3130\ : Span4Mux_v
    port map (
            O => \N__24009\,
            I => \N__24006\
        );

    \I__3129\ : Odrv4
    port map (
            O => \N__24006\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__3128\ : CascadeMux
    port map (
            O => \N__24003\,
            I => \N__24000\
        );

    \I__3127\ : InMux
    port map (
            O => \N__24000\,
            I => \N__23996\
        );

    \I__3126\ : InMux
    port map (
            O => \N__23999\,
            I => \N__23993\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__23996\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__23993\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__3123\ : InMux
    port map (
            O => \N__23988\,
            I => \N__23984\
        );

    \I__3122\ : InMux
    port map (
            O => \N__23987\,
            I => \N__23981\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__23984\,
            I => \phase_controller_inst2.state_RNI9M3OZ0Z_0\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__23981\,
            I => \phase_controller_inst2.state_RNI9M3OZ0Z_0\
        );

    \I__3119\ : InMux
    port map (
            O => \N__23976\,
            I => \bfn_8_15_0_\
        );

    \I__3118\ : InMux
    port map (
            O => \N__23973\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__3117\ : InMux
    port map (
            O => \N__23970\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__3116\ : InMux
    port map (
            O => \N__23967\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__3115\ : InMux
    port map (
            O => \N__23964\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__3114\ : InMux
    port map (
            O => \N__23961\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__3113\ : CascadeMux
    port map (
            O => \N__23958\,
            I => \N__23955\
        );

    \I__3112\ : InMux
    port map (
            O => \N__23955\,
            I => \N__23952\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__23952\,
            I => \N__23949\
        );

    \I__3110\ : Odrv12
    port map (
            O => \N__23949\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\
        );

    \I__3109\ : CascadeMux
    port map (
            O => \N__23946\,
            I => \N__23943\
        );

    \I__3108\ : InMux
    port map (
            O => \N__23943\,
            I => \N__23938\
        );

    \I__3107\ : InMux
    port map (
            O => \N__23942\,
            I => \N__23935\
        );

    \I__3106\ : InMux
    port map (
            O => \N__23941\,
            I => \N__23932\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__23938\,
            I => \N__23928\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__23935\,
            I => \N__23925\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__23932\,
            I => \N__23922\
        );

    \I__3102\ : InMux
    port map (
            O => \N__23931\,
            I => \N__23918\
        );

    \I__3101\ : Span4Mux_v
    port map (
            O => \N__23928\,
            I => \N__23911\
        );

    \I__3100\ : Span4Mux_v
    port map (
            O => \N__23925\,
            I => \N__23911\
        );

    \I__3099\ : Span4Mux_v
    port map (
            O => \N__23922\,
            I => \N__23911\
        );

    \I__3098\ : InMux
    port map (
            O => \N__23921\,
            I => \N__23908\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__23918\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__3096\ : Odrv4
    port map (
            O => \N__23911\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__23908\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__3094\ : CascadeMux
    port map (
            O => \N__23901\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20_cascade_\
        );

    \I__3093\ : CascadeMux
    port map (
            O => \N__23898\,
            I => \N__23887\
        );

    \I__3092\ : CascadeMux
    port map (
            O => \N__23897\,
            I => \N__23883\
        );

    \I__3091\ : CascadeMux
    port map (
            O => \N__23896\,
            I => \N__23879\
        );

    \I__3090\ : CascadeMux
    port map (
            O => \N__23895\,
            I => \N__23875\
        );

    \I__3089\ : CascadeMux
    port map (
            O => \N__23894\,
            I => \N__23871\
        );

    \I__3088\ : CascadeMux
    port map (
            O => \N__23893\,
            I => \N__23867\
        );

    \I__3087\ : CascadeMux
    port map (
            O => \N__23892\,
            I => \N__23863\
        );

    \I__3086\ : InMux
    port map (
            O => \N__23891\,
            I => \N__23844\
        );

    \I__3085\ : InMux
    port map (
            O => \N__23890\,
            I => \N__23844\
        );

    \I__3084\ : InMux
    port map (
            O => \N__23887\,
            I => \N__23844\
        );

    \I__3083\ : InMux
    port map (
            O => \N__23886\,
            I => \N__23844\
        );

    \I__3082\ : InMux
    port map (
            O => \N__23883\,
            I => \N__23844\
        );

    \I__3081\ : InMux
    port map (
            O => \N__23882\,
            I => \N__23844\
        );

    \I__3080\ : InMux
    port map (
            O => \N__23879\,
            I => \N__23844\
        );

    \I__3079\ : InMux
    port map (
            O => \N__23878\,
            I => \N__23844\
        );

    \I__3078\ : InMux
    port map (
            O => \N__23875\,
            I => \N__23827\
        );

    \I__3077\ : InMux
    port map (
            O => \N__23874\,
            I => \N__23827\
        );

    \I__3076\ : InMux
    port map (
            O => \N__23871\,
            I => \N__23827\
        );

    \I__3075\ : InMux
    port map (
            O => \N__23870\,
            I => \N__23827\
        );

    \I__3074\ : InMux
    port map (
            O => \N__23867\,
            I => \N__23827\
        );

    \I__3073\ : InMux
    port map (
            O => \N__23866\,
            I => \N__23827\
        );

    \I__3072\ : InMux
    port map (
            O => \N__23863\,
            I => \N__23827\
        );

    \I__3071\ : InMux
    port map (
            O => \N__23862\,
            I => \N__23827\
        );

    \I__3070\ : CascadeMux
    port map (
            O => \N__23861\,
            I => \N__23824\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__23844\,
            I => \N__23818\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__23827\,
            I => \N__23818\
        );

    \I__3067\ : InMux
    port map (
            O => \N__23824\,
            I => \N__23813\
        );

    \I__3066\ : InMux
    port map (
            O => \N__23823\,
            I => \N__23813\
        );

    \I__3065\ : Span12Mux_v
    port map (
            O => \N__23818\,
            I => \N__23808\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__23813\,
            I => \N__23808\
        );

    \I__3063\ : Odrv12
    port map (
            O => \N__23808\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__3062\ : CascadeMux
    port map (
            O => \N__23805\,
            I => \N__23802\
        );

    \I__3061\ : InMux
    port map (
            O => \N__23802\,
            I => \N__23798\
        );

    \I__3060\ : InMux
    port map (
            O => \N__23801\,
            I => \N__23794\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__23798\,
            I => \N__23791\
        );

    \I__3058\ : InMux
    port map (
            O => \N__23797\,
            I => \N__23788\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__23794\,
            I => \N__23783\
        );

    \I__3056\ : Span4Mux_v
    port map (
            O => \N__23791\,
            I => \N__23780\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__23788\,
            I => \N__23777\
        );

    \I__3054\ : InMux
    port map (
            O => \N__23787\,
            I => \N__23772\
        );

    \I__3053\ : InMux
    port map (
            O => \N__23786\,
            I => \N__23772\
        );

    \I__3052\ : Odrv4
    port map (
            O => \N__23783\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__3051\ : Odrv4
    port map (
            O => \N__23780\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__3050\ : Odrv12
    port map (
            O => \N__23777\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__23772\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__3048\ : InMux
    port map (
            O => \N__23763\,
            I => \N__23760\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__23760\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\
        );

    \I__3046\ : InMux
    port map (
            O => \N__23757\,
            I => \N__23754\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__23754\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\
        );

    \I__3044\ : CascadeMux
    port map (
            O => \N__23751\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13_cascade_\
        );

    \I__3043\ : CascadeMux
    port map (
            O => \N__23748\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_\
        );

    \I__3042\ : InMux
    port map (
            O => \N__23745\,
            I => \N__23742\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__23742\,
            I => \current_shift_inst.PI_CTRL.N_72\
        );

    \I__3040\ : InMux
    port map (
            O => \N__23739\,
            I => \N__23736\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__23736\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\
        );

    \I__3038\ : CascadeMux
    port map (
            O => \N__23733\,
            I => \N__23730\
        );

    \I__3037\ : InMux
    port map (
            O => \N__23730\,
            I => \N__23726\
        );

    \I__3036\ : InMux
    port map (
            O => \N__23729\,
            I => \N__23722\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__23726\,
            I => \N__23717\
        );

    \I__3034\ : InMux
    port map (
            O => \N__23725\,
            I => \N__23714\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__23722\,
            I => \N__23711\
        );

    \I__3032\ : InMux
    port map (
            O => \N__23721\,
            I => \N__23706\
        );

    \I__3031\ : InMux
    port map (
            O => \N__23720\,
            I => \N__23706\
        );

    \I__3030\ : Odrv12
    port map (
            O => \N__23717\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__23714\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__3028\ : Odrv4
    port map (
            O => \N__23711\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__23706\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__3026\ : CascadeMux
    port map (
            O => \N__23697\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_\
        );

    \I__3025\ : CascadeMux
    port map (
            O => \N__23694\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12_cascade_\
        );

    \I__3024\ : InMux
    port map (
            O => \N__23691\,
            I => \N__23688\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__23688\,
            I => \N__23685\
        );

    \I__3022\ : Odrv4
    port map (
            O => \N__23685\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10\
        );

    \I__3021\ : InMux
    port map (
            O => \N__23682\,
            I => \N__23679\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__23679\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\
        );

    \I__3019\ : InMux
    port map (
            O => \N__23676\,
            I => \N__23673\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__23673\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\
        );

    \I__3017\ : InMux
    port map (
            O => \N__23670\,
            I => \N__23667\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__23667\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\
        );

    \I__3015\ : InMux
    port map (
            O => \N__23664\,
            I => \N__23661\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__23661\,
            I => \phase_controller_inst2.start_timer_hc_RNO_0_0\
        );

    \I__3013\ : InMux
    port map (
            O => \N__23658\,
            I => \N__23655\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__23655\,
            I => \N__23652\
        );

    \I__3011\ : Odrv4
    port map (
            O => \N__23652\,
            I => \phase_controller_inst2.start_timer_hc_0_sqmuxa\
        );

    \I__3010\ : CascadeMux
    port map (
            O => \N__23649\,
            I => \N__23646\
        );

    \I__3009\ : InMux
    port map (
            O => \N__23646\,
            I => \N__23638\
        );

    \I__3008\ : InMux
    port map (
            O => \N__23645\,
            I => \N__23638\
        );

    \I__3007\ : InMux
    port map (
            O => \N__23644\,
            I => \N__23635\
        );

    \I__3006\ : InMux
    port map (
            O => \N__23643\,
            I => \N__23632\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__23638\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__23635\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__23632\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__3002\ : InMux
    port map (
            O => \N__23625\,
            I => \N__23622\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__23622\,
            I => \N__23618\
        );

    \I__3000\ : InMux
    port map (
            O => \N__23621\,
            I => \N__23615\
        );

    \I__2999\ : Span4Mux_s1_v
    port map (
            O => \N__23618\,
            I => \N__23610\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__23615\,
            I => \N__23610\
        );

    \I__2997\ : Span4Mux_v
    port map (
            O => \N__23610\,
            I => \N__23605\
        );

    \I__2996\ : InMux
    port map (
            O => \N__23609\,
            I => \N__23602\
        );

    \I__2995\ : InMux
    port map (
            O => \N__23608\,
            I => \N__23599\
        );

    \I__2994\ : Span4Mux_h
    port map (
            O => \N__23605\,
            I => \N__23596\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__23602\,
            I => \N__23591\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__23599\,
            I => \N__23591\
        );

    \I__2991\ : Sp12to4
    port map (
            O => \N__23596\,
            I => \N__23588\
        );

    \I__2990\ : Span4Mux_v
    port map (
            O => \N__23591\,
            I => \N__23585\
        );

    \I__2989\ : Span12Mux_v
    port map (
            O => \N__23588\,
            I => \N__23582\
        );

    \I__2988\ : Sp12to4
    port map (
            O => \N__23585\,
            I => \N__23579\
        );

    \I__2987\ : Span12Mux_v
    port map (
            O => \N__23582\,
            I => \N__23576\
        );

    \I__2986\ : Span12Mux_h
    port map (
            O => \N__23579\,
            I => \N__23573\
        );

    \I__2985\ : Span12Mux_h
    port map (
            O => \N__23576\,
            I => \N__23570\
        );

    \I__2984\ : Span12Mux_v
    port map (
            O => \N__23573\,
            I => \N__23567\
        );

    \I__2983\ : Odrv12
    port map (
            O => \N__23570\,
            I => start_stop_c
        );

    \I__2982\ : Odrv12
    port map (
            O => \N__23567\,
            I => start_stop_c
        );

    \I__2981\ : InMux
    port map (
            O => \N__23562\,
            I => \N__23559\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__23559\,
            I => \N__23555\
        );

    \I__2979\ : InMux
    port map (
            O => \N__23558\,
            I => \N__23550\
        );

    \I__2978\ : Span12Mux_s6_v
    port map (
            O => \N__23555\,
            I => \N__23547\
        );

    \I__2977\ : InMux
    port map (
            O => \N__23554\,
            I => \N__23542\
        );

    \I__2976\ : InMux
    port map (
            O => \N__23553\,
            I => \N__23542\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__23550\,
            I => \N__23539\
        );

    \I__2974\ : Odrv12
    port map (
            O => \N__23547\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__23542\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__2972\ : Odrv4
    port map (
            O => \N__23539\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__2971\ : IoInMux
    port map (
            O => \N__23532\,
            I => \N__23529\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__23529\,
            I => \N__23526\
        );

    \I__2969\ : Span4Mux_s3_v
    port map (
            O => \N__23526\,
            I => \N__23523\
        );

    \I__2968\ : Odrv4
    port map (
            O => \N__23523\,
            I => s4_phy_c
        );

    \I__2967\ : InMux
    port map (
            O => \N__23520\,
            I => \N__23517\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__23517\,
            I => \N__23514\
        );

    \I__2965\ : Odrv12
    port map (
            O => \N__23514\,
            I => il_max_comp1_c
        );

    \I__2964\ : InMux
    port map (
            O => \N__23511\,
            I => \N__23508\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__23508\,
            I => \il_max_comp1_D1\
        );

    \I__2962\ : InMux
    port map (
            O => \N__23505\,
            I => \N__23498\
        );

    \I__2961\ : InMux
    port map (
            O => \N__23504\,
            I => \N__23498\
        );

    \I__2960\ : InMux
    port map (
            O => \N__23503\,
            I => \N__23495\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__23498\,
            I => \N__23492\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__23495\,
            I => \N__23489\
        );

    \I__2957\ : Odrv4
    port map (
            O => \N__23492\,
            I => \il_max_comp2_D2\
        );

    \I__2956\ : Odrv4
    port map (
            O => \N__23489\,
            I => \il_max_comp2_D2\
        );

    \I__2955\ : InMux
    port map (
            O => \N__23484\,
            I => \N__23478\
        );

    \I__2954\ : InMux
    port map (
            O => \N__23483\,
            I => \N__23478\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__23478\,
            I => \N__23474\
        );

    \I__2952\ : InMux
    port map (
            O => \N__23477\,
            I => \N__23471\
        );

    \I__2951\ : Odrv4
    port map (
            O => \N__23474\,
            I => \il_min_comp2_D2\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__23471\,
            I => \il_min_comp2_D2\
        );

    \I__2949\ : InMux
    port map (
            O => \N__23466\,
            I => \N__23459\
        );

    \I__2948\ : InMux
    port map (
            O => \N__23465\,
            I => \N__23459\
        );

    \I__2947\ : InMux
    port map (
            O => \N__23464\,
            I => \N__23456\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__23459\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__23456\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__2944\ : IoInMux
    port map (
            O => \N__23451\,
            I => \N__23448\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__23448\,
            I => \N__23445\
        );

    \I__2942\ : Span4Mux_s3_v
    port map (
            O => \N__23445\,
            I => \N__23442\
        );

    \I__2941\ : Span4Mux_v
    port map (
            O => \N__23442\,
            I => \N__23439\
        );

    \I__2940\ : Span4Mux_v
    port map (
            O => \N__23439\,
            I => \N__23436\
        );

    \I__2939\ : Span4Mux_v
    port map (
            O => \N__23436\,
            I => \N__23433\
        );

    \I__2938\ : Odrv4
    port map (
            O => \N__23433\,
            I => \delay_measurement_inst.delay_hc_timer.N_393_i\
        );

    \I__2937\ : InMux
    port map (
            O => \N__23430\,
            I => \N__23427\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__23427\,
            I => \N__23424\
        );

    \I__2935\ : Span4Mux_h
    port map (
            O => \N__23424\,
            I => \N__23421\
        );

    \I__2934\ : Odrv4
    port map (
            O => \N__23421\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__2933\ : InMux
    port map (
            O => \N__23418\,
            I => \N__23415\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__23415\,
            I => \N__23411\
        );

    \I__2931\ : InMux
    port map (
            O => \N__23414\,
            I => \N__23408\
        );

    \I__2930\ : Odrv4
    port map (
            O => \N__23411\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__23408\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2928\ : CascadeMux
    port map (
            O => \N__23403\,
            I => \N__23400\
        );

    \I__2927\ : InMux
    port map (
            O => \N__23400\,
            I => \N__23396\
        );

    \I__2926\ : InMux
    port map (
            O => \N__23399\,
            I => \N__23393\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__23396\,
            I => \N__23388\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__23393\,
            I => \N__23388\
        );

    \I__2923\ : Odrv4
    port map (
            O => \N__23388\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2922\ : InMux
    port map (
            O => \N__23385\,
            I => \N__23382\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__23382\,
            I => \N__23379\
        );

    \I__2920\ : Span4Mux_h
    port map (
            O => \N__23379\,
            I => \N__23376\
        );

    \I__2919\ : Odrv4
    port map (
            O => \N__23376\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\
        );

    \I__2918\ : InMux
    port map (
            O => \N__23373\,
            I => \N__23370\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__23370\,
            I => \N__23367\
        );

    \I__2916\ : Odrv12
    port map (
            O => \N__23367\,
            I => \il_min_comp2_D1\
        );

    \I__2915\ : InMux
    port map (
            O => \N__23364\,
            I => \N__23361\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__23361\,
            I => \phase_controller_inst2.start_timer_tr_0_sqmuxa\
        );

    \I__2913\ : InMux
    port map (
            O => \N__23358\,
            I => \N__23355\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__23355\,
            I => \N__23352\
        );

    \I__2911\ : Span4Mux_h
    port map (
            O => \N__23352\,
            I => \N__23349\
        );

    \I__2910\ : Odrv4
    port map (
            O => \N__23349\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__2909\ : InMux
    port map (
            O => \N__23346\,
            I => \N__23343\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__23343\,
            I => \N__23340\
        );

    \I__2907\ : Odrv4
    port map (
            O => \N__23340\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__2906\ : InMux
    port map (
            O => \N__23337\,
            I => \N__23334\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__23334\,
            I => \N__23331\
        );

    \I__2904\ : Odrv4
    port map (
            O => \N__23331\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\
        );

    \I__2903\ : CascadeMux
    port map (
            O => \N__23328\,
            I => \N__23325\
        );

    \I__2902\ : InMux
    port map (
            O => \N__23325\,
            I => \N__23322\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__23322\,
            I => \N__23319\
        );

    \I__2900\ : Odrv4
    port map (
            O => \N__23319\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\
        );

    \I__2899\ : InMux
    port map (
            O => \N__23316\,
            I => \N__23313\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__23313\,
            I => \N__23310\
        );

    \I__2897\ : Odrv4
    port map (
            O => \N__23310\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\
        );

    \I__2896\ : CascadeMux
    port map (
            O => \N__23307\,
            I => \N__23304\
        );

    \I__2895\ : InMux
    port map (
            O => \N__23304\,
            I => \N__23301\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__23301\,
            I => \N__23298\
        );

    \I__2893\ : Odrv4
    port map (
            O => \N__23298\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__2892\ : InMux
    port map (
            O => \N__23295\,
            I => \N__23292\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__23292\,
            I => \N__23289\
        );

    \I__2890\ : Odrv4
    port map (
            O => \N__23289\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__2889\ : InMux
    port map (
            O => \N__23286\,
            I => \N__23283\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__23283\,
            I => \N__23280\
        );

    \I__2887\ : Odrv4
    port map (
            O => \N__23280\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__2886\ : CascadeMux
    port map (
            O => \N__23277\,
            I => \N__23274\
        );

    \I__2885\ : InMux
    port map (
            O => \N__23274\,
            I => \N__23271\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__23271\,
            I => \N__23268\
        );

    \I__2883\ : Odrv4
    port map (
            O => \N__23268\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__2882\ : InMux
    port map (
            O => \N__23265\,
            I => \N__23262\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__23262\,
            I => \N__23259\
        );

    \I__2880\ : Span12Mux_v
    port map (
            O => \N__23259\,
            I => \N__23256\
        );

    \I__2879\ : Odrv12
    port map (
            O => \N__23256\,
            I => \il_max_comp2_D1\
        );

    \I__2878\ : InMux
    port map (
            O => \N__23253\,
            I => \N__23250\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__23250\,
            I => \N__23247\
        );

    \I__2876\ : Odrv12
    port map (
            O => \N__23247\,
            I => il_min_comp2_c
        );

    \I__2875\ : CascadeMux
    port map (
            O => \N__23244\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\
        );

    \I__2874\ : InMux
    port map (
            O => \N__23241\,
            I => \N__23235\
        );

    \I__2873\ : InMux
    port map (
            O => \N__23240\,
            I => \N__23235\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__23235\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__2871\ : InMux
    port map (
            O => \N__23232\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__2870\ : CascadeMux
    port map (
            O => \N__23229\,
            I => \N__23225\
        );

    \I__2869\ : CascadeMux
    port map (
            O => \N__23228\,
            I => \N__23222\
        );

    \I__2868\ : InMux
    port map (
            O => \N__23225\,
            I => \N__23219\
        );

    \I__2867\ : InMux
    port map (
            O => \N__23222\,
            I => \N__23216\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__23219\,
            I => \N__23211\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__23216\,
            I => \N__23211\
        );

    \I__2864\ : Odrv4
    port map (
            O => \N__23211\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__2863\ : InMux
    port map (
            O => \N__23208\,
            I => \bfn_5_12_0_\
        );

    \I__2862\ : CascadeMux
    port map (
            O => \N__23205\,
            I => \N__23201\
        );

    \I__2861\ : InMux
    port map (
            O => \N__23204\,
            I => \N__23198\
        );

    \I__2860\ : InMux
    port map (
            O => \N__23201\,
            I => \N__23195\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__23198\,
            I => \N__23192\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__23195\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__2857\ : Odrv4
    port map (
            O => \N__23192\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__2856\ : InMux
    port map (
            O => \N__23187\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\
        );

    \I__2855\ : InMux
    port map (
            O => \N__23184\,
            I => \N__23180\
        );

    \I__2854\ : InMux
    port map (
            O => \N__23183\,
            I => \N__23177\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__23180\,
            I => \N__23174\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__23177\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__2851\ : Odrv4
    port map (
            O => \N__23174\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__2850\ : InMux
    port map (
            O => \N__23169\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__2849\ : InMux
    port map (
            O => \N__23166\,
            I => \N__23160\
        );

    \I__2848\ : InMux
    port map (
            O => \N__23165\,
            I => \N__23160\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__23160\,
            I => \N__23157\
        );

    \I__2846\ : Odrv4
    port map (
            O => \N__23157\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2845\ : InMux
    port map (
            O => \N__23154\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__2844\ : InMux
    port map (
            O => \N__23151\,
            I => \N__23147\
        );

    \I__2843\ : InMux
    port map (
            O => \N__23150\,
            I => \N__23144\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__23147\,
            I => \N__23141\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__23144\,
            I => \N__23138\
        );

    \I__2840\ : Span4Mux_h
    port map (
            O => \N__23141\,
            I => \N__23135\
        );

    \I__2839\ : Odrv4
    port map (
            O => \N__23138\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2838\ : Odrv4
    port map (
            O => \N__23135\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2837\ : InMux
    port map (
            O => \N__23130\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\
        );

    \I__2836\ : InMux
    port map (
            O => \N__23127\,
            I => \N__23121\
        );

    \I__2835\ : InMux
    port map (
            O => \N__23126\,
            I => \N__23121\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__23121\,
            I => \N__23118\
        );

    \I__2833\ : Odrv4
    port map (
            O => \N__23118\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2832\ : InMux
    port map (
            O => \N__23115\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__2831\ : InMux
    port map (
            O => \N__23112\,
            I => \N__23106\
        );

    \I__2830\ : InMux
    port map (
            O => \N__23111\,
            I => \N__23106\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__23106\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2828\ : InMux
    port map (
            O => \N__23103\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__2827\ : InMux
    port map (
            O => \N__23100\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__2826\ : InMux
    port map (
            O => \N__23097\,
            I => \N__23091\
        );

    \I__2825\ : InMux
    port map (
            O => \N__23096\,
            I => \N__23091\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__23091\,
            I => \N__23083\
        );

    \I__2823\ : InMux
    port map (
            O => \N__23090\,
            I => \N__23078\
        );

    \I__2822\ : InMux
    port map (
            O => \N__23089\,
            I => \N__23078\
        );

    \I__2821\ : InMux
    port map (
            O => \N__23088\,
            I => \N__23075\
        );

    \I__2820\ : InMux
    port map (
            O => \N__23087\,
            I => \N__23072\
        );

    \I__2819\ : InMux
    port map (
            O => \N__23086\,
            I => \N__23069\
        );

    \I__2818\ : Span4Mux_s2_h
    port map (
            O => \N__23083\,
            I => \N__23055\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__23078\,
            I => \N__23055\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__23075\,
            I => \N__23055\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__23072\,
            I => \N__23055\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__23069\,
            I => \N__23055\
        );

    \I__2813\ : InMux
    port map (
            O => \N__23068\,
            I => \N__23050\
        );

    \I__2812\ : InMux
    port map (
            O => \N__23067\,
            I => \N__23050\
        );

    \I__2811\ : InMux
    port map (
            O => \N__23066\,
            I => \N__23047\
        );

    \I__2810\ : Sp12to4
    port map (
            O => \N__23055\,
            I => \N__23040\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__23050\,
            I => \N__23040\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__23047\,
            I => \N__23040\
        );

    \I__2807\ : Span12Mux_s11_v
    port map (
            O => \N__23040\,
            I => \N__23037\
        );

    \I__2806\ : Odrv12
    port map (
            O => \N__23037\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2805\ : InMux
    port map (
            O => \N__23034\,
            I => \N__23030\
        );

    \I__2804\ : InMux
    port map (
            O => \N__23033\,
            I => \N__23027\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__23030\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__23027\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2801\ : InMux
    port map (
            O => \N__23022\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__2800\ : CascadeMux
    port map (
            O => \N__23019\,
            I => \N__23015\
        );

    \I__2799\ : InMux
    port map (
            O => \N__23018\,
            I => \N__23012\
        );

    \I__2798\ : InMux
    port map (
            O => \N__23015\,
            I => \N__23009\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__23012\,
            I => \N__23006\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__23009\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2795\ : Odrv4
    port map (
            O => \N__23006\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2794\ : InMux
    port map (
            O => \N__23001\,
            I => \bfn_5_11_0_\
        );

    \I__2793\ : InMux
    port map (
            O => \N__22998\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\
        );

    \I__2792\ : InMux
    port map (
            O => \N__22995\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__2791\ : CascadeMux
    port map (
            O => \N__22992\,
            I => \N__22988\
        );

    \I__2790\ : InMux
    port map (
            O => \N__22991\,
            I => \N__22985\
        );

    \I__2789\ : InMux
    port map (
            O => \N__22988\,
            I => \N__22982\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__22985\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__22982\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2786\ : InMux
    port map (
            O => \N__22977\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__2785\ : InMux
    port map (
            O => \N__22974\,
            I => \N__22970\
        );

    \I__2784\ : InMux
    port map (
            O => \N__22973\,
            I => \N__22967\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__22970\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__22967\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2781\ : InMux
    port map (
            O => \N__22962\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\
        );

    \I__2780\ : InMux
    port map (
            O => \N__22959\,
            I => \N__22955\
        );

    \I__2779\ : InMux
    port map (
            O => \N__22958\,
            I => \N__22952\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__22955\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__22952\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2776\ : InMux
    port map (
            O => \N__22947\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__2775\ : InMux
    port map (
            O => \N__22944\,
            I => \N__22940\
        );

    \I__2774\ : InMux
    port map (
            O => \N__22943\,
            I => \N__22937\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__22940\,
            I => \N__22934\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__22937\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2771\ : Odrv4
    port map (
            O => \N__22934\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2770\ : InMux
    port map (
            O => \N__22929\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__2769\ : InMux
    port map (
            O => \N__22926\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__2768\ : CascadeMux
    port map (
            O => \N__22923\,
            I => \N__22920\
        );

    \I__2767\ : InMux
    port map (
            O => \N__22920\,
            I => \N__22915\
        );

    \I__2766\ : InMux
    port map (
            O => \N__22919\,
            I => \N__22912\
        );

    \I__2765\ : InMux
    port map (
            O => \N__22918\,
            I => \N__22909\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__22915\,
            I => \N__22906\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__22912\,
            I => \N__22901\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__22909\,
            I => \N__22901\
        );

    \I__2761\ : Span4Mux_h
    port map (
            O => \N__22906\,
            I => \N__22898\
        );

    \I__2760\ : Span12Mux_s8_v
    port map (
            O => \N__22901\,
            I => \N__22895\
        );

    \I__2759\ : Odrv4
    port map (
            O => \N__22898\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2758\ : Odrv12
    port map (
            O => \N__22895\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2757\ : InMux
    port map (
            O => \N__22890\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__2756\ : InMux
    port map (
            O => \N__22887\,
            I => \N__22882\
        );

    \I__2755\ : InMux
    port map (
            O => \N__22886\,
            I => \N__22879\
        );

    \I__2754\ : InMux
    port map (
            O => \N__22885\,
            I => \N__22876\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__22882\,
            I => \N__22873\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__22879\,
            I => \N__22868\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__22876\,
            I => \N__22868\
        );

    \I__2750\ : Span4Mux_h
    port map (
            O => \N__22873\,
            I => \N__22865\
        );

    \I__2749\ : Span4Mux_h
    port map (
            O => \N__22868\,
            I => \N__22862\
        );

    \I__2748\ : Odrv4
    port map (
            O => \N__22865\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2747\ : Odrv4
    port map (
            O => \N__22862\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2746\ : InMux
    port map (
            O => \N__22857\,
            I => \bfn_5_10_0_\
        );

    \I__2745\ : InMux
    port map (
            O => \N__22854\,
            I => \N__22850\
        );

    \I__2744\ : InMux
    port map (
            O => \N__22853\,
            I => \N__22847\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__22850\,
            I => \N__22841\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__22847\,
            I => \N__22841\
        );

    \I__2741\ : InMux
    port map (
            O => \N__22846\,
            I => \N__22838\
        );

    \I__2740\ : Span4Mux_v
    port map (
            O => \N__22841\,
            I => \N__22833\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__22838\,
            I => \N__22833\
        );

    \I__2738\ : Span4Mux_h
    port map (
            O => \N__22833\,
            I => \N__22830\
        );

    \I__2737\ : Odrv4
    port map (
            O => \N__22830\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2736\ : InMux
    port map (
            O => \N__22827\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\
        );

    \I__2735\ : InMux
    port map (
            O => \N__22824\,
            I => \N__22818\
        );

    \I__2734\ : InMux
    port map (
            O => \N__22823\,
            I => \N__22818\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__22818\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__2732\ : InMux
    port map (
            O => \N__22815\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__2731\ : InMux
    port map (
            O => \N__22812\,
            I => \N__22806\
        );

    \I__2730\ : InMux
    port map (
            O => \N__22811\,
            I => \N__22806\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__22806\,
            I => \N__22803\
        );

    \I__2728\ : Odrv4
    port map (
            O => \N__22803\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2727\ : InMux
    port map (
            O => \N__22800\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__2726\ : CascadeMux
    port map (
            O => \N__22797\,
            I => \N__22794\
        );

    \I__2725\ : InMux
    port map (
            O => \N__22794\,
            I => \N__22788\
        );

    \I__2724\ : InMux
    port map (
            O => \N__22793\,
            I => \N__22788\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__22788\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2722\ : InMux
    port map (
            O => \N__22785\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\
        );

    \I__2721\ : InMux
    port map (
            O => \N__22782\,
            I => \N__22776\
        );

    \I__2720\ : InMux
    port map (
            O => \N__22781\,
            I => \N__22776\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__22776\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2718\ : InMux
    port map (
            O => \N__22773\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__2717\ : InMux
    port map (
            O => \N__22770\,
            I => \N__22764\
        );

    \I__2716\ : InMux
    port map (
            O => \N__22769\,
            I => \N__22764\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__22764\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2714\ : InMux
    port map (
            O => \N__22761\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__2713\ : InMux
    port map (
            O => \N__22758\,
            I => \N__22755\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__22755\,
            I => \N__22752\
        );

    \I__2711\ : Span4Mux_h
    port map (
            O => \N__22752\,
            I => \N__22749\
        );

    \I__2710\ : Odrv4
    port map (
            O => \N__22749\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__2709\ : InMux
    port map (
            O => \N__22746\,
            I => \N__22743\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__22743\,
            I => \N__22740\
        );

    \I__2707\ : Odrv12
    port map (
            O => \N__22740\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__2706\ : InMux
    port map (
            O => \N__22737\,
            I => \N__22734\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__22734\,
            I => \N__22731\
        );

    \I__2704\ : Span4Mux_h
    port map (
            O => \N__22731\,
            I => \N__22728\
        );

    \I__2703\ : Odrv4
    port map (
            O => \N__22728\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__2702\ : InMux
    port map (
            O => \N__22725\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\
        );

    \I__2701\ : InMux
    port map (
            O => \N__22722\,
            I => \N__22719\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__22719\,
            I => \N__22716\
        );

    \I__2699\ : Span4Mux_h
    port map (
            O => \N__22716\,
            I => \N__22713\
        );

    \I__2698\ : Odrv4
    port map (
            O => \N__22713\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__2697\ : InMux
    port map (
            O => \N__22710\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\
        );

    \I__2696\ : InMux
    port map (
            O => \N__22707\,
            I => \N__22704\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__22704\,
            I => \N__22699\
        );

    \I__2694\ : InMux
    port map (
            O => \N__22703\,
            I => \N__22696\
        );

    \I__2693\ : InMux
    port map (
            O => \N__22702\,
            I => \N__22693\
        );

    \I__2692\ : Span4Mux_s2_h
    port map (
            O => \N__22699\,
            I => \N__22688\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__22696\,
            I => \N__22688\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__22693\,
            I => \N__22685\
        );

    \I__2689\ : Span4Mux_h
    port map (
            O => \N__22688\,
            I => \N__22682\
        );

    \I__2688\ : Span4Mux_h
    port map (
            O => \N__22685\,
            I => \N__22679\
        );

    \I__2687\ : Odrv4
    port map (
            O => \N__22682\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2686\ : Odrv4
    port map (
            O => \N__22679\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2685\ : InMux
    port map (
            O => \N__22674\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__22671\,
            I => \N__22668\
        );

    \I__2683\ : InMux
    port map (
            O => \N__22668\,
            I => \N__22665\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__22665\,
            I => \N__22661\
        );

    \I__2681\ : InMux
    port map (
            O => \N__22664\,
            I => \N__22658\
        );

    \I__2680\ : Span4Mux_v
    port map (
            O => \N__22661\,
            I => \N__22651\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__22658\,
            I => \N__22651\
        );

    \I__2678\ : InMux
    port map (
            O => \N__22657\,
            I => \N__22646\
        );

    \I__2677\ : InMux
    port map (
            O => \N__22656\,
            I => \N__22646\
        );

    \I__2676\ : Span4Mux_s2_h
    port map (
            O => \N__22651\,
            I => \N__22641\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__22646\,
            I => \N__22641\
        );

    \I__2674\ : Span4Mux_h
    port map (
            O => \N__22641\,
            I => \N__22638\
        );

    \I__2673\ : Odrv4
    port map (
            O => \N__22638\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2672\ : InMux
    port map (
            O => \N__22635\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\
        );

    \I__2671\ : CascadeMux
    port map (
            O => \N__22632\,
            I => \N__22629\
        );

    \I__2670\ : InMux
    port map (
            O => \N__22629\,
            I => \N__22626\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__22626\,
            I => \N__22621\
        );

    \I__2668\ : InMux
    port map (
            O => \N__22625\,
            I => \N__22618\
        );

    \I__2667\ : InMux
    port map (
            O => \N__22624\,
            I => \N__22615\
        );

    \I__2666\ : Span4Mux_v
    port map (
            O => \N__22621\,
            I => \N__22610\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__22618\,
            I => \N__22610\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__22615\,
            I => \N__22607\
        );

    \I__2663\ : Span4Mux_h
    port map (
            O => \N__22610\,
            I => \N__22604\
        );

    \I__2662\ : Span4Mux_h
    port map (
            O => \N__22607\,
            I => \N__22601\
        );

    \I__2661\ : Odrv4
    port map (
            O => \N__22604\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2660\ : Odrv4
    port map (
            O => \N__22601\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2659\ : InMux
    port map (
            O => \N__22596\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__2658\ : CascadeMux
    port map (
            O => \N__22593\,
            I => \N__22590\
        );

    \I__2657\ : InMux
    port map (
            O => \N__22590\,
            I => \N__22586\
        );

    \I__2656\ : InMux
    port map (
            O => \N__22589\,
            I => \N__22582\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__22586\,
            I => \N__22579\
        );

    \I__2654\ : InMux
    port map (
            O => \N__22585\,
            I => \N__22576\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__22582\,
            I => \N__22573\
        );

    \I__2652\ : Span4Mux_v
    port map (
            O => \N__22579\,
            I => \N__22568\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__22576\,
            I => \N__22568\
        );

    \I__2650\ : Span4Mux_h
    port map (
            O => \N__22573\,
            I => \N__22565\
        );

    \I__2649\ : Span4Mux_h
    port map (
            O => \N__22568\,
            I => \N__22562\
        );

    \I__2648\ : Odrv4
    port map (
            O => \N__22565\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2647\ : Odrv4
    port map (
            O => \N__22562\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2646\ : InMux
    port map (
            O => \N__22557\,
            I => \N__22552\
        );

    \I__2645\ : InMux
    port map (
            O => \N__22556\,
            I => \N__22549\
        );

    \I__2644\ : InMux
    port map (
            O => \N__22555\,
            I => \N__22546\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__22552\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__22549\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__22546\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2640\ : InMux
    port map (
            O => \N__22539\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__2639\ : InMux
    port map (
            O => \N__22536\,
            I => \N__22531\
        );

    \I__2638\ : InMux
    port map (
            O => \N__22535\,
            I => \N__22528\
        );

    \I__2637\ : InMux
    port map (
            O => \N__22534\,
            I => \N__22525\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__22531\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__22528\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__22525\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2633\ : InMux
    port map (
            O => \N__22518\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__2632\ : InMux
    port map (
            O => \N__22515\,
            I => \N__22510\
        );

    \I__2631\ : InMux
    port map (
            O => \N__22514\,
            I => \N__22507\
        );

    \I__2630\ : InMux
    port map (
            O => \N__22513\,
            I => \N__22504\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__22510\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__22507\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__22504\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2626\ : InMux
    port map (
            O => \N__22497\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__2625\ : InMux
    port map (
            O => \N__22494\,
            I => \N__22489\
        );

    \I__2624\ : InMux
    port map (
            O => \N__22493\,
            I => \N__22486\
        );

    \I__2623\ : InMux
    port map (
            O => \N__22492\,
            I => \N__22483\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__22489\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__22486\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__22483\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2619\ : InMux
    port map (
            O => \N__22476\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__2618\ : InMux
    port map (
            O => \N__22473\,
            I => \N__22468\
        );

    \I__2617\ : InMux
    port map (
            O => \N__22472\,
            I => \N__22465\
        );

    \I__2616\ : InMux
    port map (
            O => \N__22471\,
            I => \N__22462\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__22468\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__22465\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__22462\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2612\ : InMux
    port map (
            O => \N__22455\,
            I => \bfn_4_13_0_\
        );

    \I__2611\ : InMux
    port map (
            O => \N__22452\,
            I => \N__22434\
        );

    \I__2610\ : InMux
    port map (
            O => \N__22451\,
            I => \N__22434\
        );

    \I__2609\ : InMux
    port map (
            O => \N__22450\,
            I => \N__22434\
        );

    \I__2608\ : InMux
    port map (
            O => \N__22449\,
            I => \N__22434\
        );

    \I__2607\ : InMux
    port map (
            O => \N__22448\,
            I => \N__22429\
        );

    \I__2606\ : InMux
    port map (
            O => \N__22447\,
            I => \N__22429\
        );

    \I__2605\ : InMux
    port map (
            O => \N__22446\,
            I => \N__22420\
        );

    \I__2604\ : InMux
    port map (
            O => \N__22445\,
            I => \N__22420\
        );

    \I__2603\ : InMux
    port map (
            O => \N__22444\,
            I => \N__22420\
        );

    \I__2602\ : InMux
    port map (
            O => \N__22443\,
            I => \N__22420\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__22434\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__22429\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__22420\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__2598\ : InMux
    port map (
            O => \N__22413\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__2597\ : InMux
    port map (
            O => \N__22410\,
            I => \N__22405\
        );

    \I__2596\ : InMux
    port map (
            O => \N__22409\,
            I => \N__22402\
        );

    \I__2595\ : InMux
    port map (
            O => \N__22408\,
            I => \N__22399\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__22405\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__22402\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__22399\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2591\ : CascadeMux
    port map (
            O => \N__22392\,
            I => \N__22389\
        );

    \I__2590\ : InMux
    port map (
            O => \N__22389\,
            I => \N__22386\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__22386\,
            I => \N__22382\
        );

    \I__2588\ : InMux
    port map (
            O => \N__22385\,
            I => \N__22379\
        );

    \I__2587\ : Span4Mux_h
    port map (
            O => \N__22382\,
            I => \N__22374\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__22379\,
            I => \N__22374\
        );

    \I__2585\ : Span4Mux_v
    port map (
            O => \N__22374\,
            I => \N__22371\
        );

    \I__2584\ : Span4Mux_h
    port map (
            O => \N__22371\,
            I => \N__22368\
        );

    \I__2583\ : Span4Mux_v
    port map (
            O => \N__22368\,
            I => \N__22365\
        );

    \I__2582\ : Odrv4
    port map (
            O => \N__22365\,
            I => \pwm_generator_inst.O_10\
        );

    \I__2581\ : InMux
    port map (
            O => \N__22362\,
            I => \N__22358\
        );

    \I__2580\ : InMux
    port map (
            O => \N__22361\,
            I => \N__22354\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__22358\,
            I => \N__22351\
        );

    \I__2578\ : InMux
    port map (
            O => \N__22357\,
            I => \N__22348\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__22354\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__2576\ : Odrv12
    port map (
            O => \N__22351\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__22348\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__2574\ : InMux
    port map (
            O => \N__22341\,
            I => \N__22338\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__22338\,
            I => \N__22335\
        );

    \I__2572\ : Odrv12
    port map (
            O => \N__22335\,
            I => il_max_comp2_c
        );

    \I__2571\ : InMux
    port map (
            O => \N__22332\,
            I => \N__22329\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__22329\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__2569\ : CascadeMux
    port map (
            O => \N__22326\,
            I => \N__22323\
        );

    \I__2568\ : InMux
    port map (
            O => \N__22323\,
            I => \N__22320\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__22320\,
            I => \N__22317\
        );

    \I__2566\ : Odrv4
    port map (
            O => \N__22317\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\
        );

    \I__2565\ : InMux
    port map (
            O => \N__22314\,
            I => \N__22311\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__22311\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\
        );

    \I__2563\ : CascadeMux
    port map (
            O => \N__22308\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_\
        );

    \I__2562\ : InMux
    port map (
            O => \N__22305\,
            I => \N__22302\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__22302\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\
        );

    \I__2560\ : InMux
    port map (
            O => \N__22299\,
            I => \N__22294\
        );

    \I__2559\ : InMux
    port map (
            O => \N__22298\,
            I => \N__22291\
        );

    \I__2558\ : InMux
    port map (
            O => \N__22297\,
            I => \N__22288\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__22294\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__22291\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__22288\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2554\ : InMux
    port map (
            O => \N__22281\,
            I => \bfn_4_12_0_\
        );

    \I__2553\ : InMux
    port map (
            O => \N__22278\,
            I => \N__22273\
        );

    \I__2552\ : InMux
    port map (
            O => \N__22277\,
            I => \N__22270\
        );

    \I__2551\ : InMux
    port map (
            O => \N__22276\,
            I => \N__22267\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__22273\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__22270\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__22267\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2547\ : InMux
    port map (
            O => \N__22260\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__2546\ : InMux
    port map (
            O => \N__22257\,
            I => \N__22252\
        );

    \I__2545\ : InMux
    port map (
            O => \N__22256\,
            I => \N__22249\
        );

    \I__2544\ : InMux
    port map (
            O => \N__22255\,
            I => \N__22246\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__22252\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__22249\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__22246\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2540\ : InMux
    port map (
            O => \N__22239\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__2539\ : InMux
    port map (
            O => \N__22236\,
            I => \N__22231\
        );

    \I__2538\ : InMux
    port map (
            O => \N__22235\,
            I => \N__22228\
        );

    \I__2537\ : InMux
    port map (
            O => \N__22234\,
            I => \N__22225\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__22231\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__22228\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__22225\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2533\ : InMux
    port map (
            O => \N__22218\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__2532\ : CascadeMux
    port map (
            O => \N__22215\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\
        );

    \I__2531\ : InMux
    port map (
            O => \N__22212\,
            I => \N__22209\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__22209\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\
        );

    \I__2529\ : CascadeMux
    port map (
            O => \N__22206\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_\
        );

    \I__2528\ : InMux
    port map (
            O => \N__22203\,
            I => \N__22195\
        );

    \I__2527\ : InMux
    port map (
            O => \N__22202\,
            I => \N__22195\
        );

    \I__2526\ : CascadeMux
    port map (
            O => \N__22201\,
            I => \N__22190\
        );

    \I__2525\ : CascadeMux
    port map (
            O => \N__22200\,
            I => \N__22187\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__22195\,
            I => \N__22181\
        );

    \I__2523\ : InMux
    port map (
            O => \N__22194\,
            I => \N__22174\
        );

    \I__2522\ : InMux
    port map (
            O => \N__22193\,
            I => \N__22174\
        );

    \I__2521\ : InMux
    port map (
            O => \N__22190\,
            I => \N__22174\
        );

    \I__2520\ : InMux
    port map (
            O => \N__22187\,
            I => \N__22171\
        );

    \I__2519\ : InMux
    port map (
            O => \N__22186\,
            I => \N__22168\
        );

    \I__2518\ : InMux
    port map (
            O => \N__22185\,
            I => \N__22165\
        );

    \I__2517\ : InMux
    port map (
            O => \N__22184\,
            I => \N__22162\
        );

    \I__2516\ : Span4Mux_v
    port map (
            O => \N__22181\,
            I => \N__22159\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__22174\,
            I => \N__22154\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__22171\,
            I => \N__22154\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__22168\,
            I => \N__22151\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__22165\,
            I => \N__22146\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__22162\,
            I => \N__22146\
        );

    \I__2510\ : Span4Mux_h
    port map (
            O => \N__22159\,
            I => \N__22143\
        );

    \I__2509\ : Span4Mux_h
    port map (
            O => \N__22154\,
            I => \N__22140\
        );

    \I__2508\ : Span4Mux_h
    port map (
            O => \N__22151\,
            I => \N__22137\
        );

    \I__2507\ : Span4Mux_h
    port map (
            O => \N__22146\,
            I => \N__22134\
        );

    \I__2506\ : Odrv4
    port map (
            O => \N__22143\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2505\ : Odrv4
    port map (
            O => \N__22140\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2504\ : Odrv4
    port map (
            O => \N__22137\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2503\ : Odrv4
    port map (
            O => \N__22134\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2502\ : InMux
    port map (
            O => \N__22125\,
            I => \N__22122\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__22122\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\
        );

    \I__2500\ : CascadeMux
    port map (
            O => \N__22119\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\
        );

    \I__2499\ : InMux
    port map (
            O => \N__22116\,
            I => \N__22113\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__22113\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\
        );

    \I__2497\ : InMux
    port map (
            O => \N__22110\,
            I => \N__22107\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__22107\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\
        );

    \I__2495\ : InMux
    port map (
            O => \N__22104\,
            I => \N__22101\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__22101\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\
        );

    \I__2493\ : InMux
    port map (
            O => \N__22098\,
            I => \N__22095\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__22095\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\
        );

    \I__2491\ : InMux
    port map (
            O => \N__22092\,
            I => \N__22089\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__22089\,
            I => \N__22086\
        );

    \I__2489\ : Odrv12
    port map (
            O => \N__22086\,
            I => \pwm_generator_inst.thresholdZ0Z_5\
        );

    \I__2488\ : InMux
    port map (
            O => \N__22083\,
            I => \N__22080\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__22080\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_0\
        );

    \I__2486\ : InMux
    port map (
            O => \N__22077\,
            I => \N__22074\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__22074\,
            I => \N__22071\
        );

    \I__2484\ : Span12Mux_s11_v
    port map (
            O => \N__22071\,
            I => \N__22068\
        );

    \I__2483\ : Odrv12
    port map (
            O => \N__22068\,
            I => \pwm_generator_inst.thresholdZ0Z_0\
        );

    \I__2482\ : InMux
    port map (
            O => \N__22065\,
            I => \N__22062\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__22062\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\
        );

    \I__2480\ : InMux
    port map (
            O => \N__22059\,
            I => \N__22056\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__22056\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_5\
        );

    \I__2478\ : CascadeMux
    port map (
            O => \N__22053\,
            I => \N__22050\
        );

    \I__2477\ : InMux
    port map (
            O => \N__22050\,
            I => \N__22047\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__22047\,
            I => \N__22044\
        );

    \I__2475\ : Odrv12
    port map (
            O => \N__22044\,
            I => \pwm_generator_inst.thresholdZ0Z_9\
        );

    \I__2474\ : InMux
    port map (
            O => \N__22041\,
            I => \N__22038\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__22038\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\
        );

    \I__2472\ : InMux
    port map (
            O => \N__22035\,
            I => \N__22032\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__22032\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_9\
        );

    \I__2470\ : InMux
    port map (
            O => \N__22029\,
            I => \N__22026\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__22026\,
            I => \N__22023\
        );

    \I__2468\ : Odrv12
    port map (
            O => \N__22023\,
            I => \pwm_generator_inst.thresholdZ0Z_8\
        );

    \I__2467\ : InMux
    port map (
            O => \N__22020\,
            I => \N__22013\
        );

    \I__2466\ : InMux
    port map (
            O => \N__22019\,
            I => \N__22013\
        );

    \I__2465\ : InMux
    port map (
            O => \N__22018\,
            I => \N__22010\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__22013\,
            I => \N__22005\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__22010\,
            I => \N__22002\
        );

    \I__2462\ : InMux
    port map (
            O => \N__22009\,
            I => \N__21997\
        );

    \I__2461\ : InMux
    port map (
            O => \N__22008\,
            I => \N__21997\
        );

    \I__2460\ : Span4Mux_v
    port map (
            O => \N__22005\,
            I => \N__21990\
        );

    \I__2459\ : Span4Mux_s3_h
    port map (
            O => \N__22002\,
            I => \N__21990\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__21997\,
            I => \N__21990\
        );

    \I__2457\ : Span4Mux_v
    port map (
            O => \N__21990\,
            I => \N__21982\
        );

    \I__2456\ : InMux
    port map (
            O => \N__21989\,
            I => \N__21979\
        );

    \I__2455\ : InMux
    port map (
            O => \N__21988\,
            I => \N__21976\
        );

    \I__2454\ : InMux
    port map (
            O => \N__21987\,
            I => \N__21969\
        );

    \I__2453\ : InMux
    port map (
            O => \N__21986\,
            I => \N__21969\
        );

    \I__2452\ : InMux
    port map (
            O => \N__21985\,
            I => \N__21969\
        );

    \I__2451\ : Span4Mux_v
    port map (
            O => \N__21982\,
            I => \N__21966\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__21979\,
            I => \N__21961\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__21976\,
            I => \N__21961\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__21969\,
            I => \N__21958\
        );

    \I__2447\ : Odrv4
    port map (
            O => \N__21966\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2446\ : Odrv12
    port map (
            O => \N__21961\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2445\ : Odrv4
    port map (
            O => \N__21958\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2444\ : CascadeMux
    port map (
            O => \N__21951\,
            I => \N__21944\
        );

    \I__2443\ : CascadeMux
    port map (
            O => \N__21950\,
            I => \N__21940\
        );

    \I__2442\ : CascadeMux
    port map (
            O => \N__21949\,
            I => \N__21936\
        );

    \I__2441\ : CascadeMux
    port map (
            O => \N__21948\,
            I => \N__21933\
        );

    \I__2440\ : InMux
    port map (
            O => \N__21947\,
            I => \N__21928\
        );

    \I__2439\ : InMux
    port map (
            O => \N__21944\,
            I => \N__21928\
        );

    \I__2438\ : InMux
    port map (
            O => \N__21943\,
            I => \N__21908\
        );

    \I__2437\ : InMux
    port map (
            O => \N__21940\,
            I => \N__21905\
        );

    \I__2436\ : CascadeMux
    port map (
            O => \N__21939\,
            I => \N__21902\
        );

    \I__2435\ : InMux
    port map (
            O => \N__21936\,
            I => \N__21897\
        );

    \I__2434\ : InMux
    port map (
            O => \N__21933\,
            I => \N__21897\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__21928\,
            I => \N__21894\
        );

    \I__2432\ : InMux
    port map (
            O => \N__21927\,
            I => \N__21888\
        );

    \I__2431\ : InMux
    port map (
            O => \N__21926\,
            I => \N__21871\
        );

    \I__2430\ : InMux
    port map (
            O => \N__21925\,
            I => \N__21871\
        );

    \I__2429\ : InMux
    port map (
            O => \N__21924\,
            I => \N__21871\
        );

    \I__2428\ : InMux
    port map (
            O => \N__21923\,
            I => \N__21871\
        );

    \I__2427\ : InMux
    port map (
            O => \N__21922\,
            I => \N__21871\
        );

    \I__2426\ : InMux
    port map (
            O => \N__21921\,
            I => \N__21871\
        );

    \I__2425\ : InMux
    port map (
            O => \N__21920\,
            I => \N__21871\
        );

    \I__2424\ : InMux
    port map (
            O => \N__21919\,
            I => \N__21871\
        );

    \I__2423\ : InMux
    port map (
            O => \N__21918\,
            I => \N__21856\
        );

    \I__2422\ : InMux
    port map (
            O => \N__21917\,
            I => \N__21856\
        );

    \I__2421\ : InMux
    port map (
            O => \N__21916\,
            I => \N__21856\
        );

    \I__2420\ : InMux
    port map (
            O => \N__21915\,
            I => \N__21856\
        );

    \I__2419\ : InMux
    port map (
            O => \N__21914\,
            I => \N__21856\
        );

    \I__2418\ : InMux
    port map (
            O => \N__21913\,
            I => \N__21856\
        );

    \I__2417\ : InMux
    port map (
            O => \N__21912\,
            I => \N__21856\
        );

    \I__2416\ : CascadeMux
    port map (
            O => \N__21911\,
            I => \N__21848\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__21908\,
            I => \N__21843\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__21905\,
            I => \N__21843\
        );

    \I__2413\ : InMux
    port map (
            O => \N__21902\,
            I => \N__21840\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__21897\,
            I => \N__21837\
        );

    \I__2411\ : Span4Mux_h
    port map (
            O => \N__21894\,
            I => \N__21834\
        );

    \I__2410\ : CascadeMux
    port map (
            O => \N__21893\,
            I => \N__21831\
        );

    \I__2409\ : InMux
    port map (
            O => \N__21892\,
            I => \N__21826\
        );

    \I__2408\ : InMux
    port map (
            O => \N__21891\,
            I => \N__21826\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__21888\,
            I => \N__21819\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__21871\,
            I => \N__21819\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__21856\,
            I => \N__21819\
        );

    \I__2404\ : InMux
    port map (
            O => \N__21855\,
            I => \N__21812\
        );

    \I__2403\ : InMux
    port map (
            O => \N__21854\,
            I => \N__21812\
        );

    \I__2402\ : InMux
    port map (
            O => \N__21853\,
            I => \N__21812\
        );

    \I__2401\ : InMux
    port map (
            O => \N__21852\,
            I => \N__21805\
        );

    \I__2400\ : InMux
    port map (
            O => \N__21851\,
            I => \N__21805\
        );

    \I__2399\ : InMux
    port map (
            O => \N__21848\,
            I => \N__21805\
        );

    \I__2398\ : Span4Mux_v
    port map (
            O => \N__21843\,
            I => \N__21802\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__21840\,
            I => \N__21795\
        );

    \I__2396\ : Span12Mux_h
    port map (
            O => \N__21837\,
            I => \N__21795\
        );

    \I__2395\ : Sp12to4
    port map (
            O => \N__21834\,
            I => \N__21795\
        );

    \I__2394\ : InMux
    port map (
            O => \N__21831\,
            I => \N__21792\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__21826\,
            I => \N__21789\
        );

    \I__2392\ : Span4Mux_v
    port map (
            O => \N__21819\,
            I => \N__21784\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__21812\,
            I => \N__21784\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__21805\,
            I => \N_19_1\
        );

    \I__2389\ : Odrv4
    port map (
            O => \N__21802\,
            I => \N_19_1\
        );

    \I__2388\ : Odrv12
    port map (
            O => \N__21795\,
            I => \N_19_1\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__21792\,
            I => \N_19_1\
        );

    \I__2386\ : Odrv4
    port map (
            O => \N__21789\,
            I => \N_19_1\
        );

    \I__2385\ : Odrv4
    port map (
            O => \N__21784\,
            I => \N_19_1\
        );

    \I__2384\ : CascadeMux
    port map (
            O => \N__21771\,
            I => \N__21768\
        );

    \I__2383\ : InMux
    port map (
            O => \N__21768\,
            I => \N__21765\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__21765\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\
        );

    \I__2381\ : InMux
    port map (
            O => \N__21762\,
            I => \N__21753\
        );

    \I__2380\ : InMux
    port map (
            O => \N__21761\,
            I => \N__21753\
        );

    \I__2379\ : InMux
    port map (
            O => \N__21760\,
            I => \N__21748\
        );

    \I__2378\ : InMux
    port map (
            O => \N__21759\,
            I => \N__21748\
        );

    \I__2377\ : InMux
    port map (
            O => \N__21758\,
            I => \N__21745\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__21753\,
            I => \N__21742\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__21748\,
            I => \N__21737\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__21745\,
            I => \N__21732\
        );

    \I__2373\ : Span4Mux_h
    port map (
            O => \N__21742\,
            I => \N__21732\
        );

    \I__2372\ : InMux
    port map (
            O => \N__21741\,
            I => \N__21729\
        );

    \I__2371\ : InMux
    port map (
            O => \N__21740\,
            I => \N__21726\
        );

    \I__2370\ : Span12Mux_s6_h
    port map (
            O => \N__21737\,
            I => \N__21720\
        );

    \I__2369\ : Span4Mux_v
    port map (
            O => \N__21732\,
            I => \N__21713\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__21729\,
            I => \N__21713\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__21726\,
            I => \N__21713\
        );

    \I__2366\ : InMux
    port map (
            O => \N__21725\,
            I => \N__21706\
        );

    \I__2365\ : InMux
    port map (
            O => \N__21724\,
            I => \N__21706\
        );

    \I__2364\ : InMux
    port map (
            O => \N__21723\,
            I => \N__21706\
        );

    \I__2363\ : Span12Mux_v
    port map (
            O => \N__21720\,
            I => \N__21703\
        );

    \I__2362\ : Span4Mux_v
    port map (
            O => \N__21713\,
            I => \N__21698\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__21706\,
            I => \N__21698\
        );

    \I__2360\ : Odrv12
    port map (
            O => \N__21703\,
            I => \pwm_generator_inst.N_17\
        );

    \I__2359\ : Odrv4
    port map (
            O => \N__21698\,
            I => \pwm_generator_inst.N_17\
        );

    \I__2358\ : InMux
    port map (
            O => \N__21693\,
            I => \N__21690\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__21690\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_8\
        );

    \I__2356\ : InMux
    port map (
            O => \N__21687\,
            I => \N__21682\
        );

    \I__2355\ : InMux
    port map (
            O => \N__21686\,
            I => \N__21679\
        );

    \I__2354\ : InMux
    port map (
            O => \N__21685\,
            I => \N__21676\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__21682\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__21679\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__21676\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__2350\ : InMux
    port map (
            O => \N__21669\,
            I => \N__21666\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__21666\,
            I => \N__21663\
        );

    \I__2348\ : Span4Mux_v
    port map (
            O => \N__21663\,
            I => \N__21660\
        );

    \I__2347\ : Odrv4
    port map (
            O => \N__21660\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\
        );

    \I__2346\ : InMux
    port map (
            O => \N__21657\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_11\
        );

    \I__2345\ : InMux
    port map (
            O => \N__21654\,
            I => \N__21650\
        );

    \I__2344\ : InMux
    port map (
            O => \N__21653\,
            I => \N__21646\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__21650\,
            I => \N__21643\
        );

    \I__2342\ : InMux
    port map (
            O => \N__21649\,
            I => \N__21640\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__21646\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__2340\ : Odrv4
    port map (
            O => \N__21643\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__21640\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__2338\ : InMux
    port map (
            O => \N__21633\,
            I => \N__21630\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__21630\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\
        );

    \I__2336\ : InMux
    port map (
            O => \N__21627\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_12\
        );

    \I__2335\ : InMux
    port map (
            O => \N__21624\,
            I => \N__21621\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__21621\,
            I => \N__21616\
        );

    \I__2333\ : InMux
    port map (
            O => \N__21620\,
            I => \N__21613\
        );

    \I__2332\ : InMux
    port map (
            O => \N__21619\,
            I => \N__21610\
        );

    \I__2331\ : Span4Mux_s3_h
    port map (
            O => \N__21616\,
            I => \N__21605\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__21613\,
            I => \N__21605\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__21610\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__2328\ : Odrv4
    port map (
            O => \N__21605\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__2327\ : InMux
    port map (
            O => \N__21600\,
            I => \N__21597\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__21597\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\
        );

    \I__2325\ : InMux
    port map (
            O => \N__21594\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_13\
        );

    \I__2324\ : InMux
    port map (
            O => \N__21591\,
            I => \N__21587\
        );

    \I__2323\ : InMux
    port map (
            O => \N__21590\,
            I => \N__21584\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__21587\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__21584\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__2320\ : InMux
    port map (
            O => \N__21579\,
            I => \N__21576\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__21576\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\
        );

    \I__2318\ : InMux
    port map (
            O => \N__21573\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_14\
        );

    \I__2317\ : InMux
    port map (
            O => \N__21570\,
            I => \N__21566\
        );

    \I__2316\ : InMux
    port map (
            O => \N__21569\,
            I => \N__21563\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__21566\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__21563\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__2313\ : InMux
    port map (
            O => \N__21558\,
            I => \N__21555\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__21555\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\
        );

    \I__2311\ : InMux
    port map (
            O => \N__21552\,
            I => \bfn_3_17_0_\
        );

    \I__2310\ : InMux
    port map (
            O => \N__21549\,
            I => \N__21545\
        );

    \I__2309\ : InMux
    port map (
            O => \N__21548\,
            I => \N__21542\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__21545\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__21542\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__2306\ : InMux
    port map (
            O => \N__21537\,
            I => \N__21534\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__21534\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\
        );

    \I__2304\ : InMux
    port map (
            O => \N__21531\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_16\
        );

    \I__2303\ : InMux
    port map (
            O => \N__21528\,
            I => \N__21523\
        );

    \I__2302\ : InMux
    port map (
            O => \N__21527\,
            I => \N__21520\
        );

    \I__2301\ : InMux
    port map (
            O => \N__21526\,
            I => \N__21517\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__21523\,
            I => \N__21514\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__21520\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__21517\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__2297\ : Odrv4
    port map (
            O => \N__21514\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__2296\ : InMux
    port map (
            O => \N__21507\,
            I => \N__21504\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__21504\,
            I => \N__21501\
        );

    \I__2294\ : Odrv4
    port map (
            O => \N__21501\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\
        );

    \I__2293\ : InMux
    port map (
            O => \N__21498\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_17\
        );

    \I__2292\ : InMux
    port map (
            O => \N__21495\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_18\
        );

    \I__2291\ : InMux
    port map (
            O => \N__21492\,
            I => \N__21489\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__21489\,
            I => \N__21486\
        );

    \I__2289\ : Odrv4
    port map (
            O => \N__21486\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\
        );

    \I__2288\ : InMux
    port map (
            O => \N__21483\,
            I => \N__21480\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__21480\,
            I => \N__21477\
        );

    \I__2286\ : Sp12to4
    port map (
            O => \N__21477\,
            I => \N__21474\
        );

    \I__2285\ : Span12Mux_v
    port map (
            O => \N__21474\,
            I => \N__21471\
        );

    \I__2284\ : Odrv12
    port map (
            O => \N__21471\,
            I => \pwm_generator_inst.O_4\
        );

    \I__2283\ : InMux
    port map (
            O => \N__21468\,
            I => \N__21465\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__21465\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_4\
        );

    \I__2281\ : InMux
    port map (
            O => \N__21462\,
            I => \N__21459\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__21459\,
            I => \N__21456\
        );

    \I__2279\ : Span12Mux_v
    port map (
            O => \N__21456\,
            I => \N__21453\
        );

    \I__2278\ : Odrv12
    port map (
            O => \N__21453\,
            I => \pwm_generator_inst.O_5\
        );

    \I__2277\ : InMux
    port map (
            O => \N__21450\,
            I => \N__21447\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__21447\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_5\
        );

    \I__2275\ : InMux
    port map (
            O => \N__21444\,
            I => \N__21441\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__21441\,
            I => \N__21438\
        );

    \I__2273\ : Span4Mux_v
    port map (
            O => \N__21438\,
            I => \N__21435\
        );

    \I__2272\ : Span4Mux_h
    port map (
            O => \N__21435\,
            I => \N__21432\
        );

    \I__2271\ : Span4Mux_v
    port map (
            O => \N__21432\,
            I => \N__21429\
        );

    \I__2270\ : Odrv4
    port map (
            O => \N__21429\,
            I => \pwm_generator_inst.O_6\
        );

    \I__2269\ : InMux
    port map (
            O => \N__21426\,
            I => \N__21423\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__21423\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_6\
        );

    \I__2267\ : InMux
    port map (
            O => \N__21420\,
            I => \N__21417\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__21417\,
            I => \N__21414\
        );

    \I__2265\ : Span4Mux_v
    port map (
            O => \N__21414\,
            I => \N__21411\
        );

    \I__2264\ : Span4Mux_h
    port map (
            O => \N__21411\,
            I => \N__21408\
        );

    \I__2263\ : Span4Mux_v
    port map (
            O => \N__21408\,
            I => \N__21405\
        );

    \I__2262\ : Odrv4
    port map (
            O => \N__21405\,
            I => \pwm_generator_inst.O_7\
        );

    \I__2261\ : InMux
    port map (
            O => \N__21402\,
            I => \N__21399\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__21399\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_7\
        );

    \I__2259\ : InMux
    port map (
            O => \N__21396\,
            I => \N__21393\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__21393\,
            I => \N__21390\
        );

    \I__2257\ : Span4Mux_h
    port map (
            O => \N__21390\,
            I => \N__21387\
        );

    \I__2256\ : Span4Mux_v
    port map (
            O => \N__21387\,
            I => \N__21384\
        );

    \I__2255\ : Span4Mux_v
    port map (
            O => \N__21384\,
            I => \N__21381\
        );

    \I__2254\ : Odrv4
    port map (
            O => \N__21381\,
            I => \pwm_generator_inst.O_8\
        );

    \I__2253\ : InMux
    port map (
            O => \N__21378\,
            I => \N__21375\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__21375\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_8\
        );

    \I__2251\ : InMux
    port map (
            O => \N__21372\,
            I => \N__21369\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__21369\,
            I => \N__21366\
        );

    \I__2249\ : Span4Mux_h
    port map (
            O => \N__21366\,
            I => \N__21363\
        );

    \I__2248\ : Sp12to4
    port map (
            O => \N__21363\,
            I => \N__21360\
        );

    \I__2247\ : Odrv12
    port map (
            O => \N__21360\,
            I => \pwm_generator_inst.O_9\
        );

    \I__2246\ : InMux
    port map (
            O => \N__21357\,
            I => \N__21354\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__21354\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_9\
        );

    \I__2244\ : InMux
    port map (
            O => \N__21351\,
            I => \N__21348\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__21348\,
            I => \N__21345\
        );

    \I__2242\ : Span4Mux_s3_h
    port map (
            O => \N__21345\,
            I => \N__21342\
        );

    \I__2241\ : Odrv4
    port map (
            O => \N__21342\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\
        );

    \I__2240\ : InMux
    port map (
            O => \N__21339\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_9\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__21336\,
            I => \N__21332\
        );

    \I__2238\ : CascadeMux
    port map (
            O => \N__21335\,
            I => \N__21328\
        );

    \I__2237\ : InMux
    port map (
            O => \N__21332\,
            I => \N__21324\
        );

    \I__2236\ : InMux
    port map (
            O => \N__21331\,
            I => \N__21319\
        );

    \I__2235\ : InMux
    port map (
            O => \N__21328\,
            I => \N__21316\
        );

    \I__2234\ : InMux
    port map (
            O => \N__21327\,
            I => \N__21313\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__21324\,
            I => \N__21309\
        );

    \I__2232\ : InMux
    port map (
            O => \N__21323\,
            I => \N__21304\
        );

    \I__2231\ : InMux
    port map (
            O => \N__21322\,
            I => \N__21304\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__21319\,
            I => \N__21297\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__21316\,
            I => \N__21297\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__21313\,
            I => \N__21297\
        );

    \I__2227\ : InMux
    port map (
            O => \N__21312\,
            I => \N__21289\
        );

    \I__2226\ : Span4Mux_v
    port map (
            O => \N__21309\,
            I => \N__21284\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__21304\,
            I => \N__21284\
        );

    \I__2224\ : Span4Mux_v
    port map (
            O => \N__21297\,
            I => \N__21281\
        );

    \I__2223\ : InMux
    port map (
            O => \N__21296\,
            I => \N__21274\
        );

    \I__2222\ : InMux
    port map (
            O => \N__21295\,
            I => \N__21274\
        );

    \I__2221\ : InMux
    port map (
            O => \N__21294\,
            I => \N__21274\
        );

    \I__2220\ : InMux
    port map (
            O => \N__21293\,
            I => \N__21269\
        );

    \I__2219\ : InMux
    port map (
            O => \N__21292\,
            I => \N__21269\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__21289\,
            I => \N__21266\
        );

    \I__2217\ : Odrv4
    port map (
            O => \N__21284\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2216\ : Odrv4
    port map (
            O => \N__21281\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__21274\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__21269\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2213\ : Odrv12
    port map (
            O => \N__21266\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2212\ : InMux
    port map (
            O => \N__21255\,
            I => \N__21252\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__21252\,
            I => \N__21248\
        );

    \I__2210\ : InMux
    port map (
            O => \N__21251\,
            I => \N__21245\
        );

    \I__2209\ : Span4Mux_v
    port map (
            O => \N__21248\,
            I => \N__21240\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__21245\,
            I => \N__21240\
        );

    \I__2207\ : Span4Mux_v
    port map (
            O => \N__21240\,
            I => \N__21237\
        );

    \I__2206\ : Span4Mux_v
    port map (
            O => \N__21237\,
            I => \N__21234\
        );

    \I__2205\ : Odrv4
    port map (
            O => \N__21234\,
            I => \pwm_generator_inst.un3_threshold_acc\
        );

    \I__2204\ : InMux
    port map (
            O => \N__21231\,
            I => \N__21228\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__21228\,
            I => \N__21225\
        );

    \I__2202\ : Odrv4
    port map (
            O => \N__21225\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_1\
        );

    \I__2201\ : InMux
    port map (
            O => \N__21222\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_10\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__21219\,
            I => \pwm_generator_inst.un1_counterlto2_0_cascade_\
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__21216\,
            I => \pwm_generator_inst.un1_counterlto9_2_cascade_\
        );

    \I__2198\ : InMux
    port map (
            O => \N__21213\,
            I => \N__21210\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__21210\,
            I => \pwm_generator_inst.un1_counterlt9\
        );

    \I__2196\ : CascadeMux
    port map (
            O => \N__21207\,
            I => \N__21204\
        );

    \I__2195\ : InMux
    port map (
            O => \N__21204\,
            I => \N__21201\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__21201\,
            I => \N__21198\
        );

    \I__2193\ : Span4Mux_v
    port map (
            O => \N__21198\,
            I => \N__21194\
        );

    \I__2192\ : InMux
    port map (
            O => \N__21197\,
            I => \N__21191\
        );

    \I__2191\ : Odrv4
    port map (
            O => \N__21194\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__21191\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\
        );

    \I__2189\ : InMux
    port map (
            O => \N__21186\,
            I => \N__21183\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__21183\,
            I => \N__21180\
        );

    \I__2187\ : Span4Mux_h
    port map (
            O => \N__21180\,
            I => \N__21177\
        );

    \I__2186\ : Span4Mux_v
    port map (
            O => \N__21177\,
            I => \N__21174\
        );

    \I__2185\ : Span4Mux_v
    port map (
            O => \N__21174\,
            I => \N__21171\
        );

    \I__2184\ : Odrv4
    port map (
            O => \N__21171\,
            I => \pwm_generator_inst.O_0\
        );

    \I__2183\ : InMux
    port map (
            O => \N__21168\,
            I => \N__21165\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__21165\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_0\
        );

    \I__2181\ : InMux
    port map (
            O => \N__21162\,
            I => \N__21159\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__21159\,
            I => \N__21156\
        );

    \I__2179\ : Span4Mux_h
    port map (
            O => \N__21156\,
            I => \N__21153\
        );

    \I__2178\ : Sp12to4
    port map (
            O => \N__21153\,
            I => \N__21150\
        );

    \I__2177\ : Odrv12
    port map (
            O => \N__21150\,
            I => \pwm_generator_inst.O_1\
        );

    \I__2176\ : InMux
    port map (
            O => \N__21147\,
            I => \N__21144\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__21144\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_1\
        );

    \I__2174\ : InMux
    port map (
            O => \N__21141\,
            I => \N__21138\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__21138\,
            I => \N__21135\
        );

    \I__2172\ : Span12Mux_h
    port map (
            O => \N__21135\,
            I => \N__21132\
        );

    \I__2171\ : Odrv12
    port map (
            O => \N__21132\,
            I => \pwm_generator_inst.O_2\
        );

    \I__2170\ : InMux
    port map (
            O => \N__21129\,
            I => \N__21126\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__21126\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_2\
        );

    \I__2168\ : InMux
    port map (
            O => \N__21123\,
            I => \N__21120\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__21120\,
            I => \N__21117\
        );

    \I__2166\ : Span4Mux_h
    port map (
            O => \N__21117\,
            I => \N__21114\
        );

    \I__2165\ : Sp12to4
    port map (
            O => \N__21114\,
            I => \N__21111\
        );

    \I__2164\ : Odrv12
    port map (
            O => \N__21111\,
            I => \pwm_generator_inst.O_3\
        );

    \I__2163\ : InMux
    port map (
            O => \N__21108\,
            I => \N__21105\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__21105\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_3\
        );

    \I__2161\ : InMux
    port map (
            O => \N__21102\,
            I => \N__21099\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__21099\,
            I => \pwm_generator_inst.thresholdZ0Z_3\
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__21096\,
            I => \N__21093\
        );

    \I__2158\ : InMux
    port map (
            O => \N__21093\,
            I => \N__21090\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__21090\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__2156\ : InMux
    port map (
            O => \N__21087\,
            I => \N__21084\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__21084\,
            I => \N__21081\
        );

    \I__2154\ : Odrv4
    port map (
            O => \N__21081\,
            I => \pwm_generator_inst.thresholdZ0Z_4\
        );

    \I__2153\ : CascadeMux
    port map (
            O => \N__21078\,
            I => \N__21075\
        );

    \I__2152\ : InMux
    port map (
            O => \N__21075\,
            I => \N__21072\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__21072\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__2150\ : CascadeMux
    port map (
            O => \N__21069\,
            I => \N__21066\
        );

    \I__2149\ : InMux
    port map (
            O => \N__21066\,
            I => \N__21063\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__21063\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__2147\ : CascadeMux
    port map (
            O => \N__21060\,
            I => \N__21057\
        );

    \I__2146\ : InMux
    port map (
            O => \N__21057\,
            I => \N__21054\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__21054\,
            I => \pwm_generator_inst.thresholdZ0Z_6\
        );

    \I__2144\ : InMux
    port map (
            O => \N__21051\,
            I => \N__21048\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__21048\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__2142\ : InMux
    port map (
            O => \N__21045\,
            I => \N__21042\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__21042\,
            I => \N__21039\
        );

    \I__2140\ : Odrv4
    port map (
            O => \N__21039\,
            I => \pwm_generator_inst.thresholdZ0Z_7\
        );

    \I__2139\ : CascadeMux
    port map (
            O => \N__21036\,
            I => \N__21033\
        );

    \I__2138\ : InMux
    port map (
            O => \N__21033\,
            I => \N__21030\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__21030\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__2136\ : CascadeMux
    port map (
            O => \N__21027\,
            I => \N__21024\
        );

    \I__2135\ : InMux
    port map (
            O => \N__21024\,
            I => \N__21021\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__21021\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__2133\ : InMux
    port map (
            O => \N__21018\,
            I => \N__21015\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__21015\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__2131\ : InMux
    port map (
            O => \N__21012\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__2130\ : IoInMux
    port map (
            O => \N__21009\,
            I => \N__21006\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__21006\,
            I => \N__21003\
        );

    \I__2128\ : Span4Mux_s1_v
    port map (
            O => \N__21003\,
            I => \N__21000\
        );

    \I__2127\ : Sp12to4
    port map (
            O => \N__21000\,
            I => \N__20997\
        );

    \I__2126\ : Span12Mux_s10_h
    port map (
            O => \N__20997\,
            I => \N__20994\
        );

    \I__2125\ : Span12Mux_h
    port map (
            O => \N__20994\,
            I => \N__20991\
        );

    \I__2124\ : Odrv12
    port map (
            O => \N__20991\,
            I => pwm_output_c
        );

    \I__2123\ : CascadeMux
    port map (
            O => \N__20988\,
            I => \N__20985\
        );

    \I__2122\ : InMux
    port map (
            O => \N__20985\,
            I => \N__20982\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__20982\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4\
        );

    \I__2120\ : InMux
    port map (
            O => \N__20979\,
            I => \N__20972\
        );

    \I__2119\ : InMux
    port map (
            O => \N__20978\,
            I => \N__20972\
        );

    \I__2118\ : CascadeMux
    port map (
            O => \N__20977\,
            I => \N__20969\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__20972\,
            I => \N__20963\
        );

    \I__2116\ : InMux
    port map (
            O => \N__20969\,
            I => \N__20960\
        );

    \I__2115\ : InMux
    port map (
            O => \N__20968\,
            I => \N__20953\
        );

    \I__2114\ : InMux
    port map (
            O => \N__20967\,
            I => \N__20953\
        );

    \I__2113\ : InMux
    port map (
            O => \N__20966\,
            I => \N__20953\
        );

    \I__2112\ : Span4Mux_v
    port map (
            O => \N__20963\,
            I => \N__20947\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__20960\,
            I => \N__20947\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__20953\,
            I => \N__20944\
        );

    \I__2109\ : InMux
    port map (
            O => \N__20952\,
            I => \N__20941\
        );

    \I__2108\ : Span4Mux_v
    port map (
            O => \N__20947\,
            I => \N__20938\
        );

    \I__2107\ : Span4Mux_s3_h
    port map (
            O => \N__20944\,
            I => \N__20935\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__20941\,
            I => \N__20932\
        );

    \I__2105\ : Odrv4
    port map (
            O => \N__20938\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2104\ : Odrv4
    port map (
            O => \N__20935\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2103\ : Odrv4
    port map (
            O => \N__20932\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2102\ : InMux
    port map (
            O => \N__20925\,
            I => \N__20922\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__20922\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_1\
        );

    \I__2100\ : InMux
    port map (
            O => \N__20919\,
            I => \N__20916\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__20916\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_3\
        );

    \I__2098\ : InMux
    port map (
            O => \N__20913\,
            I => \N__20910\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__20910\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_2\
        );

    \I__2096\ : CascadeMux
    port map (
            O => \N__20907\,
            I => \N__20904\
        );

    \I__2095\ : InMux
    port map (
            O => \N__20904\,
            I => \N__20901\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__20901\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__2093\ : InMux
    port map (
            O => \N__20898\,
            I => \N__20895\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__20895\,
            I => \pwm_generator_inst.thresholdZ0Z_1\
        );

    \I__2091\ : CascadeMux
    port map (
            O => \N__20892\,
            I => \N__20889\
        );

    \I__2090\ : InMux
    port map (
            O => \N__20889\,
            I => \N__20886\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__20886\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__2088\ : InMux
    port map (
            O => \N__20883\,
            I => \N__20880\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__20880\,
            I => \N__20877\
        );

    \I__2086\ : Odrv4
    port map (
            O => \N__20877\,
            I => \pwm_generator_inst.thresholdZ0Z_2\
        );

    \I__2085\ : CascadeMux
    port map (
            O => \N__20874\,
            I => \N__20871\
        );

    \I__2084\ : InMux
    port map (
            O => \N__20871\,
            I => \N__20868\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__20868\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__2082\ : InMux
    port map (
            O => \N__20865\,
            I => \N__20862\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__20862\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_3\
        );

    \I__2080\ : InMux
    port map (
            O => \N__20859\,
            I => \N__20856\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__20856\,
            I => \N__20853\
        );

    \I__2078\ : Odrv12
    port map (
            O => \N__20853\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\
        );

    \I__2077\ : InMux
    port map (
            O => \N__20850\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_2\
        );

    \I__2076\ : InMux
    port map (
            O => \N__20847\,
            I => \N__20844\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__20844\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_4\
        );

    \I__2074\ : InMux
    port map (
            O => \N__20841\,
            I => \N__20838\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__20838\,
            I => \N__20835\
        );

    \I__2072\ : Odrv12
    port map (
            O => \N__20835\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\
        );

    \I__2071\ : InMux
    port map (
            O => \N__20832\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_3\
        );

    \I__2070\ : InMux
    port map (
            O => \N__20829\,
            I => \N__20826\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__20826\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_5\
        );

    \I__2068\ : InMux
    port map (
            O => \N__20823\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_4\
        );

    \I__2067\ : InMux
    port map (
            O => \N__20820\,
            I => \N__20817\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__20817\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_6\
        );

    \I__2065\ : CascadeMux
    port map (
            O => \N__20814\,
            I => \N__20811\
        );

    \I__2064\ : InMux
    port map (
            O => \N__20811\,
            I => \N__20808\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__20808\,
            I => \N__20805\
        );

    \I__2062\ : Span4Mux_v
    port map (
            O => \N__20805\,
            I => \N__20802\
        );

    \I__2061\ : Odrv4
    port map (
            O => \N__20802\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\
        );

    \I__2060\ : InMux
    port map (
            O => \N__20799\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_5\
        );

    \I__2059\ : InMux
    port map (
            O => \N__20796\,
            I => \N__20793\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__20793\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_7\
        );

    \I__2057\ : InMux
    port map (
            O => \N__20790\,
            I => \N__20787\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__20787\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\
        );

    \I__2055\ : InMux
    port map (
            O => \N__20784\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_6\
        );

    \I__2054\ : InMux
    port map (
            O => \N__20781\,
            I => \bfn_2_19_0_\
        );

    \I__2053\ : InMux
    port map (
            O => \N__20778\,
            I => \N__20775\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__20775\,
            I => \N__20772\
        );

    \I__2051\ : Odrv12
    port map (
            O => \N__20772\,
            I => \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\
        );

    \I__2050\ : InMux
    port map (
            O => \N__20769\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_8\
        );

    \I__2049\ : CascadeMux
    port map (
            O => \N__20766\,
            I => \N__20763\
        );

    \I__2048\ : InMux
    port map (
            O => \N__20763\,
            I => \N__20760\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__20760\,
            I => \N__20756\
        );

    \I__2046\ : InMux
    port map (
            O => \N__20759\,
            I => \N__20753\
        );

    \I__2045\ : Span4Mux_v
    port map (
            O => \N__20756\,
            I => \N__20748\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__20753\,
            I => \N__20748\
        );

    \I__2043\ : Odrv4
    port map (
            O => \N__20748\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\
        );

    \I__2042\ : InMux
    port map (
            O => \N__20745\,
            I => \N__20742\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__20742\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_8\
        );

    \I__2040\ : CascadeMux
    port map (
            O => \N__20739\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_\
        );

    \I__2039\ : InMux
    port map (
            O => \N__20736\,
            I => \N__20730\
        );

    \I__2038\ : InMux
    port map (
            O => \N__20735\,
            I => \N__20730\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__20730\,
            I => \N__20727\
        );

    \I__2036\ : Odrv4
    port map (
            O => \N__20727\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\
        );

    \I__2035\ : InMux
    port map (
            O => \N__20724\,
            I => \N__20718\
        );

    \I__2034\ : InMux
    port map (
            O => \N__20723\,
            I => \N__20718\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__20718\,
            I => \N__20715\
        );

    \I__2032\ : Odrv4
    port map (
            O => \N__20715\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\
        );

    \I__2031\ : CascadeMux
    port map (
            O => \N__20712\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_\
        );

    \I__2030\ : InMux
    port map (
            O => \N__20709\,
            I => \N__20703\
        );

    \I__2029\ : InMux
    port map (
            O => \N__20708\,
            I => \N__20703\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__20703\,
            I => \N__20700\
        );

    \I__2027\ : Odrv4
    port map (
            O => \N__20700\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\
        );

    \I__2026\ : CascadeMux
    port map (
            O => \N__20697\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_\
        );

    \I__2025\ : CascadeMux
    port map (
            O => \N__20694\,
            I => \N__20691\
        );

    \I__2024\ : InMux
    port map (
            O => \N__20691\,
            I => \N__20687\
        );

    \I__2023\ : InMux
    port map (
            O => \N__20690\,
            I => \N__20684\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__20687\,
            I => \N__20679\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__20684\,
            I => \N__20679\
        );

    \I__2020\ : Odrv4
    port map (
            O => \N__20679\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\
        );

    \I__2019\ : InMux
    port map (
            O => \N__20676\,
            I => \N__20673\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__20673\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_0\
        );

    \I__2017\ : CascadeMux
    port map (
            O => \N__20670\,
            I => \N__20667\
        );

    \I__2016\ : InMux
    port map (
            O => \N__20667\,
            I => \N__20664\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__20664\,
            I => \N__20661\
        );

    \I__2014\ : Odrv12
    port map (
            O => \N__20661\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\
        );

    \I__2013\ : InMux
    port map (
            O => \N__20658\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_0\
        );

    \I__2012\ : InMux
    port map (
            O => \N__20655\,
            I => \N__20652\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__20652\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_2\
        );

    \I__2010\ : CascadeMux
    port map (
            O => \N__20649\,
            I => \N__20646\
        );

    \I__2009\ : InMux
    port map (
            O => \N__20646\,
            I => \N__20643\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__20643\,
            I => \N__20640\
        );

    \I__2007\ : Odrv12
    port map (
            O => \N__20640\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\
        );

    \I__2006\ : InMux
    port map (
            O => \N__20637\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_1\
        );

    \I__2005\ : InMux
    port map (
            O => \N__20634\,
            I => \N__20631\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__20631\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\
        );

    \I__2003\ : InMux
    port map (
            O => \N__20628\,
            I => \N__20625\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__20625\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\
        );

    \I__2001\ : InMux
    port map (
            O => \N__20622\,
            I => \N__20619\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__20619\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\
        );

    \I__1999\ : InMux
    port map (
            O => \N__20616\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_19\
        );

    \I__1998\ : InMux
    port map (
            O => \N__20613\,
            I => \N__20610\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__20610\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\
        );

    \I__1996\ : CascadeMux
    port map (
            O => \N__20607\,
            I => \N__20604\
        );

    \I__1995\ : InMux
    port map (
            O => \N__20604\,
            I => \N__20601\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__20601\,
            I => \N__20597\
        );

    \I__1993\ : InMux
    port map (
            O => \N__20600\,
            I => \N__20594\
        );

    \I__1992\ : Span4Mux_v
    port map (
            O => \N__20597\,
            I => \N__20589\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__20594\,
            I => \N__20589\
        );

    \I__1990\ : Odrv4
    port map (
            O => \N__20589\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\
        );

    \I__1989\ : InMux
    port map (
            O => \N__20586\,
            I => \N__20583\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__20583\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\
        );

    \I__1987\ : InMux
    port map (
            O => \N__20580\,
            I => \bfn_2_15_0_\
        );

    \I__1986\ : InMux
    port map (
            O => \N__20577\,
            I => \N__20574\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__20574\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\
        );

    \I__1984\ : InMux
    port map (
            O => \N__20571\,
            I => \N__20568\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__20568\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\
        );

    \I__1982\ : InMux
    port map (
            O => \N__20565\,
            I => \N__20562\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__20562\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\
        );

    \I__1980\ : InMux
    port map (
            O => \N__20559\,
            I => \N__20556\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__20556\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\
        );

    \I__1978\ : InMux
    port map (
            O => \N__20553\,
            I => \N__20550\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__20550\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\
        );

    \I__1976\ : InMux
    port map (
            O => \N__20547\,
            I => \N__20544\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__20544\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\
        );

    \I__1974\ : InMux
    port map (
            O => \N__20541\,
            I => \N__20538\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__20538\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\
        );

    \I__1972\ : InMux
    port map (
            O => \N__20535\,
            I => \N__20532\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__20532\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\
        );

    \I__1970\ : InMux
    port map (
            O => \N__20529\,
            I => \N__20526\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__20526\,
            I => \N__20523\
        );

    \I__1968\ : Span4Mux_v
    port map (
            O => \N__20523\,
            I => \N__20520\
        );

    \I__1967\ : Span4Mux_v
    port map (
            O => \N__20520\,
            I => \N__20517\
        );

    \I__1966\ : Odrv4
    port map (
            O => \N__20517\,
            I => \pwm_generator_inst.O_12\
        );

    \I__1965\ : InMux
    port map (
            O => \N__20514\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0\
        );

    \I__1964\ : InMux
    port map (
            O => \N__20511\,
            I => \N__20508\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__20508\,
            I => \N__20505\
        );

    \I__1962\ : Span4Mux_v
    port map (
            O => \N__20505\,
            I => \N__20502\
        );

    \I__1961\ : Span4Mux_v
    port map (
            O => \N__20502\,
            I => \N__20499\
        );

    \I__1960\ : Odrv4
    port map (
            O => \N__20499\,
            I => \pwm_generator_inst.O_13\
        );

    \I__1959\ : InMux
    port map (
            O => \N__20496\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1\
        );

    \I__1958\ : InMux
    port map (
            O => \N__20493\,
            I => \N__20490\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__20490\,
            I => \N__20487\
        );

    \I__1956\ : Span12Mux_v
    port map (
            O => \N__20487\,
            I => \N__20484\
        );

    \I__1955\ : Odrv12
    port map (
            O => \N__20484\,
            I => \pwm_generator_inst.O_14\
        );

    \I__1954\ : InMux
    port map (
            O => \N__20481\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2\
        );

    \I__1953\ : InMux
    port map (
            O => \N__20478\,
            I => \N__20475\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__20475\,
            I => \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\
        );

    \I__1951\ : InMux
    port map (
            O => \N__20472\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3\
        );

    \I__1950\ : CascadeMux
    port map (
            O => \N__20469\,
            I => \N__20466\
        );

    \I__1949\ : InMux
    port map (
            O => \N__20466\,
            I => \N__20463\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__20463\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\
        );

    \I__1947\ : InMux
    port map (
            O => \N__20460\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4\
        );

    \I__1946\ : CascadeMux
    port map (
            O => \N__20457\,
            I => \N__20454\
        );

    \I__1945\ : InMux
    port map (
            O => \N__20454\,
            I => \N__20451\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__20451\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\
        );

    \I__1943\ : InMux
    port map (
            O => \N__20448\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5\
        );

    \I__1942\ : CascadeMux
    port map (
            O => \N__20445\,
            I => \N__20442\
        );

    \I__1941\ : InMux
    port map (
            O => \N__20442\,
            I => \N__20439\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__20439\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\
        );

    \I__1939\ : InMux
    port map (
            O => \N__20436\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6\
        );

    \I__1938\ : CascadeMux
    port map (
            O => \N__20433\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\
        );

    \I__1937\ : CascadeMux
    port map (
            O => \N__20430\,
            I => \N__20426\
        );

    \I__1936\ : CascadeMux
    port map (
            O => \N__20429\,
            I => \N__20423\
        );

    \I__1935\ : InMux
    port map (
            O => \N__20426\,
            I => \N__20420\
        );

    \I__1934\ : InMux
    port map (
            O => \N__20423\,
            I => \N__20417\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__20420\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__20417\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__1931\ : CascadeMux
    port map (
            O => \N__20412\,
            I => \current_shift_inst.PI_CTRL.N_31_cascade_\
        );

    \I__1930\ : InMux
    port map (
            O => \N__20409\,
            I => \N__20405\
        );

    \I__1929\ : InMux
    port map (
            O => \N__20408\,
            I => \N__20402\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__20405\,
            I => \N__20397\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__20402\,
            I => \N__20397\
        );

    \I__1926\ : Odrv4
    port map (
            O => \N__20397\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\
        );

    \I__1925\ : InMux
    port map (
            O => \N__20394\,
            I => \N__20391\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__20391\,
            I => \N__20388\
        );

    \I__1923\ : Span12Mux_v
    port map (
            O => \N__20388\,
            I => \N__20385\
        );

    \I__1922\ : Odrv12
    port map (
            O => \N__20385\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_7\
        );

    \I__1921\ : InMux
    port map (
            O => \N__20382\,
            I => \N__20379\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__20379\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_6\
        );

    \I__1919\ : InMux
    port map (
            O => \N__20376\,
            I => \N__20373\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__20373\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_4\
        );

    \I__1917\ : InMux
    port map (
            O => \N__20370\,
            I => \N__20363\
        );

    \I__1916\ : InMux
    port map (
            O => \N__20369\,
            I => \N__20363\
        );

    \I__1915\ : InMux
    port map (
            O => \N__20368\,
            I => \N__20360\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__20363\,
            I => pwm_duty_input_8
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__20360\,
            I => pwm_duty_input_8
        );

    \I__1912\ : InMux
    port map (
            O => \N__20355\,
            I => \N__20348\
        );

    \I__1911\ : InMux
    port map (
            O => \N__20354\,
            I => \N__20348\
        );

    \I__1910\ : InMux
    port map (
            O => \N__20353\,
            I => \N__20345\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__20348\,
            I => pwm_duty_input_9
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__20345\,
            I => pwm_duty_input_9
        );

    \I__1907\ : CascadeMux
    port map (
            O => \N__20340\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\
        );

    \I__1906\ : InMux
    port map (
            O => \N__20337\,
            I => \N__20334\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__20334\,
            I => \N__20329\
        );

    \I__1904\ : InMux
    port map (
            O => \N__20333\,
            I => \N__20324\
        );

    \I__1903\ : InMux
    port map (
            O => \N__20332\,
            I => \N__20324\
        );

    \I__1902\ : Span4Mux_s1_h
    port map (
            O => \N__20329\,
            I => \N__20321\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__20324\,
            I => pwm_duty_input_6
        );

    \I__1900\ : Odrv4
    port map (
            O => \N__20321\,
            I => pwm_duty_input_6
        );

    \I__1899\ : InMux
    port map (
            O => \N__20316\,
            I => \N__20313\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__20313\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__1897\ : CascadeMux
    port map (
            O => \N__20310\,
            I => \current_shift_inst.PI_CTRL.N_27_cascade_\
        );

    \I__1896\ : CascadeMux
    port map (
            O => \N__20307\,
            I => \N__20301\
        );

    \I__1895\ : CascadeMux
    port map (
            O => \N__20306\,
            I => \N__20298\
        );

    \I__1894\ : CascadeMux
    port map (
            O => \N__20305\,
            I => \N__20295\
        );

    \I__1893\ : CascadeMux
    port map (
            O => \N__20304\,
            I => \N__20292\
        );

    \I__1892\ : InMux
    port map (
            O => \N__20301\,
            I => \N__20287\
        );

    \I__1891\ : InMux
    port map (
            O => \N__20298\,
            I => \N__20287\
        );

    \I__1890\ : InMux
    port map (
            O => \N__20295\,
            I => \N__20283\
        );

    \I__1889\ : InMux
    port map (
            O => \N__20292\,
            I => \N__20280\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__20287\,
            I => \N__20277\
        );

    \I__1887\ : InMux
    port map (
            O => \N__20286\,
            I => \N__20274\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__20283\,
            I => \current_shift_inst.PI_CTRL.N_153\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__20280\,
            I => \current_shift_inst.PI_CTRL.N_153\
        );

    \I__1884\ : Odrv4
    port map (
            O => \N__20277\,
            I => \current_shift_inst.PI_CTRL.N_153\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__20274\,
            I => \current_shift_inst.PI_CTRL.N_153\
        );

    \I__1882\ : CascadeMux
    port map (
            O => \N__20265\,
            I => \N__20262\
        );

    \I__1881\ : InMux
    port map (
            O => \N__20262\,
            I => \N__20258\
        );

    \I__1880\ : InMux
    port map (
            O => \N__20261\,
            I => \N__20255\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__20258\,
            I => \N__20251\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__20255\,
            I => \N__20248\
        );

    \I__1877\ : InMux
    port map (
            O => \N__20254\,
            I => \N__20245\
        );

    \I__1876\ : Span4Mux_h
    port map (
            O => \N__20251\,
            I => \N__20240\
        );

    \I__1875\ : Span4Mux_s1_h
    port map (
            O => \N__20248\,
            I => \N__20240\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__20245\,
            I => pwm_duty_input_5
        );

    \I__1873\ : Odrv4
    port map (
            O => \N__20240\,
            I => pwm_duty_input_5
        );

    \I__1872\ : InMux
    port map (
            O => \N__20235\,
            I => \N__20232\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__20232\,
            I => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\
        );

    \I__1870\ : InMux
    port map (
            O => \N__20229\,
            I => \N__20226\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__20226\,
            I => \N__20223\
        );

    \I__1868\ : Odrv4
    port map (
            O => \N__20223\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\
        );

    \I__1867\ : InMux
    port map (
            O => \N__20220\,
            I => \N__20213\
        );

    \I__1866\ : InMux
    port map (
            O => \N__20219\,
            I => \N__20213\
        );

    \I__1865\ : InMux
    port map (
            O => \N__20218\,
            I => \N__20210\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__20213\,
            I => pwm_duty_input_4
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__20210\,
            I => pwm_duty_input_4
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__20205\,
            I => \N__20201\
        );

    \I__1861\ : InMux
    port map (
            O => \N__20204\,
            I => \N__20197\
        );

    \I__1860\ : InMux
    port map (
            O => \N__20201\,
            I => \N__20192\
        );

    \I__1859\ : InMux
    port map (
            O => \N__20200\,
            I => \N__20192\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__20197\,
            I => \N__20189\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__20192\,
            I => pwm_duty_input_3
        );

    \I__1856\ : Odrv4
    port map (
            O => \N__20189\,
            I => pwm_duty_input_3
        );

    \I__1855\ : InMux
    port map (
            O => \N__20184\,
            I => \N__20181\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__20181\,
            I => \N__20178\
        );

    \I__1853\ : Odrv4
    port map (
            O => \N__20178\,
            I => \pwm_generator_inst.un1_duty_inputlt3\
        );

    \I__1852\ : InMux
    port map (
            O => \N__20175\,
            I => \N__20169\
        );

    \I__1851\ : InMux
    port map (
            O => \N__20174\,
            I => \N__20169\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__20169\,
            I => \N__20165\
        );

    \I__1849\ : InMux
    port map (
            O => \N__20168\,
            I => \N__20162\
        );

    \I__1848\ : Odrv4
    port map (
            O => \N__20165\,
            I => \current_shift_inst.PI_CTRL.N_154\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__20162\,
            I => \current_shift_inst.PI_CTRL.N_154\
        );

    \I__1846\ : InMux
    port map (
            O => \N__20157\,
            I => \N__20154\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__20154\,
            I => \current_shift_inst.PI_CTRL.N_155\
        );

    \I__1844\ : InMux
    port map (
            O => \N__20151\,
            I => \bfn_1_16_0_\
        );

    \I__1843\ : InMux
    port map (
            O => \N__20148\,
            I => \N__20145\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__20145\,
            I => un7_start_stop_0_a2
        );

    \I__1841\ : InMux
    port map (
            O => \N__20142\,
            I => \N__20139\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__20139\,
            I => \N_38_i_i\
        );

    \I__1839\ : InMux
    port map (
            O => \N__20136\,
            I => \N__20132\
        );

    \I__1838\ : InMux
    port map (
            O => \N__20135\,
            I => \N__20129\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__20132\,
            I => \N__20126\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__20129\,
            I => pwm_duty_input_0
        );

    \I__1835\ : Odrv4
    port map (
            O => \N__20126\,
            I => pwm_duty_input_0
        );

    \I__1834\ : InMux
    port map (
            O => \N__20121\,
            I => \N__20117\
        );

    \I__1833\ : InMux
    port map (
            O => \N__20120\,
            I => \N__20114\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__20117\,
            I => \N__20111\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__20114\,
            I => pwm_duty_input_1
        );

    \I__1830\ : Odrv4
    port map (
            O => \N__20111\,
            I => pwm_duty_input_1
        );

    \I__1829\ : InMux
    port map (
            O => \N__20106\,
            I => \N__20102\
        );

    \I__1828\ : InMux
    port map (
            O => \N__20105\,
            I => \N__20099\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__20102\,
            I => pwm_duty_input_2
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__20099\,
            I => pwm_duty_input_2
        );

    \I__1825\ : InMux
    port map (
            O => \N__20094\,
            I => \N__20087\
        );

    \I__1824\ : InMux
    port map (
            O => \N__20093\,
            I => \N__20087\
        );

    \I__1823\ : InMux
    port map (
            O => \N__20092\,
            I => \N__20084\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__20087\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_3\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__20084\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_3\
        );

    \I__1820\ : InMux
    port map (
            O => \N__20079\,
            I => \N__20075\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__20078\,
            I => \N__20072\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__20075\,
            I => \N__20068\
        );

    \I__1817\ : InMux
    port map (
            O => \N__20072\,
            I => \N__20063\
        );

    \I__1816\ : InMux
    port map (
            O => \N__20071\,
            I => \N__20063\
        );

    \I__1815\ : Span4Mux_s2_h
    port map (
            O => \N__20068\,
            I => \N__20060\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__20063\,
            I => pwm_duty_input_7
        );

    \I__1813\ : Odrv4
    port map (
            O => \N__20060\,
            I => pwm_duty_input_7
        );

    \I__1812\ : InMux
    port map (
            O => \N__20055\,
            I => \N__20052\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__20052\,
            I => \N__20049\
        );

    \I__1810\ : Span4Mux_v
    port map (
            O => \N__20049\,
            I => \N__20046\
        );

    \I__1809\ : Odrv4
    port map (
            O => \N__20046\,
            I => \pwm_generator_inst.un2_threshold_acc_2_8\
        );

    \I__1808\ : CascadeMux
    port map (
            O => \N__20043\,
            I => \N__20040\
        );

    \I__1807\ : InMux
    port map (
            O => \N__20040\,
            I => \N__20037\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__20037\,
            I => \N__20034\
        );

    \I__1805\ : Span4Mux_v
    port map (
            O => \N__20034\,
            I => \N__20031\
        );

    \I__1804\ : Span4Mux_v
    port map (
            O => \N__20031\,
            I => \N__20028\
        );

    \I__1803\ : Odrv4
    port map (
            O => \N__20028\,
            I => \pwm_generator_inst.un2_threshold_acc_1_23\
        );

    \I__1802\ : InMux
    port map (
            O => \N__20025\,
            I => \bfn_1_15_0_\
        );

    \I__1801\ : InMux
    port map (
            O => \N__20022\,
            I => \N__20019\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__20019\,
            I => \N__20016\
        );

    \I__1799\ : Span4Mux_v
    port map (
            O => \N__20016\,
            I => \N__20013\
        );

    \I__1798\ : Odrv4
    port map (
            O => \N__20013\,
            I => \pwm_generator_inst.un2_threshold_acc_2_9\
        );

    \I__1797\ : CascadeMux
    port map (
            O => \N__20010\,
            I => \N__20007\
        );

    \I__1796\ : InMux
    port map (
            O => \N__20007\,
            I => \N__20004\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__20004\,
            I => \N__20001\
        );

    \I__1794\ : Span4Mux_v
    port map (
            O => \N__20001\,
            I => \N__19998\
        );

    \I__1793\ : Span4Mux_v
    port map (
            O => \N__19998\,
            I => \N__19995\
        );

    \I__1792\ : Odrv4
    port map (
            O => \N__19995\,
            I => \pwm_generator_inst.un2_threshold_acc_1_24\
        );

    \I__1791\ : InMux
    port map (
            O => \N__19992\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\
        );

    \I__1790\ : InMux
    port map (
            O => \N__19989\,
            I => \N__19986\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__19986\,
            I => \N__19983\
        );

    \I__1788\ : Span4Mux_v
    port map (
            O => \N__19983\,
            I => \N__19980\
        );

    \I__1787\ : Odrv4
    port map (
            O => \N__19980\,
            I => \pwm_generator_inst.un2_threshold_acc_2_10\
        );

    \I__1786\ : InMux
    port map (
            O => \N__19977\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\
        );

    \I__1785\ : CascadeMux
    port map (
            O => \N__19974\,
            I => \N__19971\
        );

    \I__1784\ : InMux
    port map (
            O => \N__19971\,
            I => \N__19968\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__19968\,
            I => \N__19965\
        );

    \I__1782\ : Span4Mux_v
    port map (
            O => \N__19965\,
            I => \N__19962\
        );

    \I__1781\ : Odrv4
    port map (
            O => \N__19962\,
            I => \pwm_generator_inst.un2_threshold_acc_2_11\
        );

    \I__1780\ : InMux
    port map (
            O => \N__19959\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\
        );

    \I__1779\ : InMux
    port map (
            O => \N__19956\,
            I => \N__19953\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__19953\,
            I => \N__19950\
        );

    \I__1777\ : Span4Mux_v
    port map (
            O => \N__19950\,
            I => \N__19947\
        );

    \I__1776\ : Odrv4
    port map (
            O => \N__19947\,
            I => \pwm_generator_inst.un2_threshold_acc_2_12\
        );

    \I__1775\ : InMux
    port map (
            O => \N__19944\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__19941\,
            I => \N__19938\
        );

    \I__1773\ : InMux
    port map (
            O => \N__19938\,
            I => \N__19935\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__19935\,
            I => \N__19932\
        );

    \I__1771\ : Span4Mux_v
    port map (
            O => \N__19932\,
            I => \N__19929\
        );

    \I__1770\ : Odrv4
    port map (
            O => \N__19929\,
            I => \pwm_generator_inst.un2_threshold_acc_2_13\
        );

    \I__1769\ : InMux
    port map (
            O => \N__19926\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\
        );

    \I__1768\ : InMux
    port map (
            O => \N__19923\,
            I => \N__19920\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__19920\,
            I => \N__19917\
        );

    \I__1766\ : Span4Mux_v
    port map (
            O => \N__19917\,
            I => \N__19914\
        );

    \I__1765\ : Odrv4
    port map (
            O => \N__19914\,
            I => \pwm_generator_inst.un2_threshold_acc_2_14\
        );

    \I__1764\ : InMux
    port map (
            O => \N__19911\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\
        );

    \I__1763\ : CascadeMux
    port map (
            O => \N__19908\,
            I => \N__19902\
        );

    \I__1762\ : CascadeMux
    port map (
            O => \N__19907\,
            I => \N__19898\
        );

    \I__1761\ : CascadeMux
    port map (
            O => \N__19906\,
            I => \N__19894\
        );

    \I__1760\ : InMux
    port map (
            O => \N__19905\,
            I => \N__19879\
        );

    \I__1759\ : InMux
    port map (
            O => \N__19902\,
            I => \N__19879\
        );

    \I__1758\ : InMux
    port map (
            O => \N__19901\,
            I => \N__19879\
        );

    \I__1757\ : InMux
    port map (
            O => \N__19898\,
            I => \N__19879\
        );

    \I__1756\ : InMux
    port map (
            O => \N__19897\,
            I => \N__19879\
        );

    \I__1755\ : InMux
    port map (
            O => \N__19894\,
            I => \N__19879\
        );

    \I__1754\ : InMux
    port map (
            O => \N__19893\,
            I => \N__19876\
        );

    \I__1753\ : InMux
    port map (
            O => \N__19892\,
            I => \N__19873\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__19879\,
            I => \N__19870\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__19876\,
            I => \N__19867\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__19873\,
            I => \N__19862\
        );

    \I__1749\ : Span4Mux_v
    port map (
            O => \N__19870\,
            I => \N__19862\
        );

    \I__1748\ : Span4Mux_v
    port map (
            O => \N__19867\,
            I => \N__19857\
        );

    \I__1747\ : Span4Mux_v
    port map (
            O => \N__19862\,
            I => \N__19857\
        );

    \I__1746\ : Odrv4
    port map (
            O => \N__19857\,
            I => \pwm_generator_inst.un2_threshold_acc_1_25\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__19854\,
            I => \N__19851\
        );

    \I__1744\ : InMux
    port map (
            O => \N__19851\,
            I => \N__19848\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__19848\,
            I => \N__19845\
        );

    \I__1742\ : Odrv12
    port map (
            O => \N__19845\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\
        );

    \I__1741\ : InMux
    port map (
            O => \N__19842\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\
        );

    \I__1740\ : InMux
    port map (
            O => \N__19839\,
            I => \N__19836\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__19836\,
            I => \N__19833\
        );

    \I__1738\ : Odrv12
    port map (
            O => \N__19833\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\
        );

    \I__1737\ : InMux
    port map (
            O => \N__19830\,
            I => \N__19827\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__19827\,
            I => \N__19824\
        );

    \I__1735\ : Span4Mux_v
    port map (
            O => \N__19824\,
            I => \N__19821\
        );

    \I__1734\ : Odrv4
    port map (
            O => \N__19821\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1\
        );

    \I__1733\ : CascadeMux
    port map (
            O => \N__19818\,
            I => \N__19815\
        );

    \I__1732\ : InMux
    port map (
            O => \N__19815\,
            I => \N__19812\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__19812\,
            I => \N__19809\
        );

    \I__1730\ : Span4Mux_v
    port map (
            O => \N__19809\,
            I => \N__19806\
        );

    \I__1729\ : Span4Mux_v
    port map (
            O => \N__19806\,
            I => \N__19803\
        );

    \I__1728\ : Odrv4
    port map (
            O => \N__19803\,
            I => \pwm_generator_inst.un2_threshold_acc_1_16\
        );

    \I__1727\ : InMux
    port map (
            O => \N__19800\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\
        );

    \I__1726\ : InMux
    port map (
            O => \N__19797\,
            I => \N__19794\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__19794\,
            I => \N__19791\
        );

    \I__1724\ : Span4Mux_v
    port map (
            O => \N__19791\,
            I => \N__19788\
        );

    \I__1723\ : Odrv4
    port map (
            O => \N__19788\,
            I => \pwm_generator_inst.un2_threshold_acc_2_2\
        );

    \I__1722\ : CascadeMux
    port map (
            O => \N__19785\,
            I => \N__19782\
        );

    \I__1721\ : InMux
    port map (
            O => \N__19782\,
            I => \N__19779\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__19779\,
            I => \N__19776\
        );

    \I__1719\ : Span4Mux_v
    port map (
            O => \N__19776\,
            I => \N__19773\
        );

    \I__1718\ : Span4Mux_v
    port map (
            O => \N__19773\,
            I => \N__19770\
        );

    \I__1717\ : Odrv4
    port map (
            O => \N__19770\,
            I => \pwm_generator_inst.un2_threshold_acc_1_17\
        );

    \I__1716\ : InMux
    port map (
            O => \N__19767\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\
        );

    \I__1715\ : InMux
    port map (
            O => \N__19764\,
            I => \N__19761\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__19761\,
            I => \N__19758\
        );

    \I__1713\ : Span4Mux_v
    port map (
            O => \N__19758\,
            I => \N__19755\
        );

    \I__1712\ : Odrv4
    port map (
            O => \N__19755\,
            I => \pwm_generator_inst.un2_threshold_acc_2_3\
        );

    \I__1711\ : CascadeMux
    port map (
            O => \N__19752\,
            I => \N__19749\
        );

    \I__1710\ : InMux
    port map (
            O => \N__19749\,
            I => \N__19746\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__19746\,
            I => \N__19743\
        );

    \I__1708\ : Span4Mux_v
    port map (
            O => \N__19743\,
            I => \N__19740\
        );

    \I__1707\ : Odrv4
    port map (
            O => \N__19740\,
            I => \pwm_generator_inst.un2_threshold_acc_1_18\
        );

    \I__1706\ : InMux
    port map (
            O => \N__19737\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\
        );

    \I__1705\ : InMux
    port map (
            O => \N__19734\,
            I => \N__19731\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__19731\,
            I => \N__19728\
        );

    \I__1703\ : Span4Mux_v
    port map (
            O => \N__19728\,
            I => \N__19725\
        );

    \I__1702\ : Odrv4
    port map (
            O => \N__19725\,
            I => \pwm_generator_inst.un2_threshold_acc_2_4\
        );

    \I__1701\ : CascadeMux
    port map (
            O => \N__19722\,
            I => \N__19719\
        );

    \I__1700\ : InMux
    port map (
            O => \N__19719\,
            I => \N__19716\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__19716\,
            I => \N__19713\
        );

    \I__1698\ : Span4Mux_h
    port map (
            O => \N__19713\,
            I => \N__19710\
        );

    \I__1697\ : Span4Mux_v
    port map (
            O => \N__19710\,
            I => \N__19707\
        );

    \I__1696\ : Odrv4
    port map (
            O => \N__19707\,
            I => \pwm_generator_inst.un2_threshold_acc_1_19\
        );

    \I__1695\ : InMux
    port map (
            O => \N__19704\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\
        );

    \I__1694\ : InMux
    port map (
            O => \N__19701\,
            I => \N__19698\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__19698\,
            I => \N__19695\
        );

    \I__1692\ : Span4Mux_v
    port map (
            O => \N__19695\,
            I => \N__19692\
        );

    \I__1691\ : Odrv4
    port map (
            O => \N__19692\,
            I => \pwm_generator_inst.un2_threshold_acc_2_5\
        );

    \I__1690\ : CascadeMux
    port map (
            O => \N__19689\,
            I => \N__19686\
        );

    \I__1689\ : InMux
    port map (
            O => \N__19686\,
            I => \N__19683\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__19683\,
            I => \N__19680\
        );

    \I__1687\ : Span4Mux_v
    port map (
            O => \N__19680\,
            I => \N__19677\
        );

    \I__1686\ : Odrv4
    port map (
            O => \N__19677\,
            I => \pwm_generator_inst.un2_threshold_acc_1_20\
        );

    \I__1685\ : InMux
    port map (
            O => \N__19674\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\
        );

    \I__1684\ : InMux
    port map (
            O => \N__19671\,
            I => \N__19668\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__19668\,
            I => \N__19665\
        );

    \I__1682\ : Span4Mux_v
    port map (
            O => \N__19665\,
            I => \N__19662\
        );

    \I__1681\ : Odrv4
    port map (
            O => \N__19662\,
            I => \pwm_generator_inst.un2_threshold_acc_2_6\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__19659\,
            I => \N__19656\
        );

    \I__1679\ : InMux
    port map (
            O => \N__19656\,
            I => \N__19653\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__19653\,
            I => \N__19650\
        );

    \I__1677\ : Span4Mux_v
    port map (
            O => \N__19650\,
            I => \N__19647\
        );

    \I__1676\ : Odrv4
    port map (
            O => \N__19647\,
            I => \pwm_generator_inst.un2_threshold_acc_1_21\
        );

    \I__1675\ : InMux
    port map (
            O => \N__19644\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\
        );

    \I__1674\ : InMux
    port map (
            O => \N__19641\,
            I => \N__19638\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__19638\,
            I => \N__19635\
        );

    \I__1672\ : Span4Mux_v
    port map (
            O => \N__19635\,
            I => \N__19632\
        );

    \I__1671\ : Odrv4
    port map (
            O => \N__19632\,
            I => \pwm_generator_inst.un2_threshold_acc_2_7\
        );

    \I__1670\ : CascadeMux
    port map (
            O => \N__19629\,
            I => \N__19626\
        );

    \I__1669\ : InMux
    port map (
            O => \N__19626\,
            I => \N__19623\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__19623\,
            I => \N__19620\
        );

    \I__1667\ : Span4Mux_v
    port map (
            O => \N__19620\,
            I => \N__19617\
        );

    \I__1666\ : Odrv4
    port map (
            O => \N__19617\,
            I => \pwm_generator_inst.un2_threshold_acc_1_22\
        );

    \I__1665\ : InMux
    port map (
            O => \N__19614\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\
        );

    \I__1664\ : InMux
    port map (
            O => \N__19611\,
            I => \N__19608\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__19608\,
            I => \N__19605\
        );

    \I__1662\ : Odrv12
    port map (
            O => \N__19605\,
            I => \current_shift_inst.PI_CTRL.N_149\
        );

    \I__1661\ : InMux
    port map (
            O => \N__19602\,
            I => \N__19599\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__19599\,
            I => \N__19596\
        );

    \I__1659\ : Odrv4
    port map (
            O => \N__19596\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_16\
        );

    \I__1658\ : InMux
    port map (
            O => \N__19593\,
            I => \N__19589\
        );

    \I__1657\ : InMux
    port map (
            O => \N__19592\,
            I => \N__19586\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__19589\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_15\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__19586\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_15\
        );

    \I__1654\ : InMux
    port map (
            O => \N__19581\,
            I => \N__19578\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__19578\,
            I => \N__19575\
        );

    \I__1652\ : Span4Mux_v
    port map (
            O => \N__19575\,
            I => \N__19572\
        );

    \I__1651\ : Odrv4
    port map (
            O => \N__19572\,
            I => \pwm_generator_inst.un2_threshold_acc_2_0\
        );

    \I__1650\ : CascadeMux
    port map (
            O => \N__19569\,
            I => \N__19566\
        );

    \I__1649\ : InMux
    port map (
            O => \N__19566\,
            I => \N__19563\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__19563\,
            I => \N__19560\
        );

    \I__1647\ : Span4Mux_v
    port map (
            O => \N__19560\,
            I => \N__19557\
        );

    \I__1646\ : Span4Mux_v
    port map (
            O => \N__19557\,
            I => \N__19554\
        );

    \I__1645\ : Odrv4
    port map (
            O => \N__19554\,
            I => \pwm_generator_inst.un2_threshold_acc_1_15\
        );

    \I__1644\ : IoInMux
    port map (
            O => \N__19551\,
            I => \N__19548\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__19548\,
            I => \N__19545\
        );

    \I__1642\ : Span4Mux_s3_v
    port map (
            O => \N__19545\,
            I => \N__19542\
        );

    \I__1641\ : Span4Mux_h
    port map (
            O => \N__19542\,
            I => \N__19539\
        );

    \I__1640\ : Sp12to4
    port map (
            O => \N__19539\,
            I => \N__19536\
        );

    \I__1639\ : Span12Mux_v
    port map (
            O => \N__19536\,
            I => \N__19533\
        );

    \I__1638\ : Span12Mux_v
    port map (
            O => \N__19533\,
            I => \N__19530\
        );

    \I__1637\ : Odrv12
    port map (
            O => \N__19530\,
            I => delay_tr_input_ibuf_gb_io_gb_input
        );

    \I__1636\ : IoInMux
    port map (
            O => \N__19527\,
            I => \N__19524\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__19524\,
            I => \N__19521\
        );

    \I__1634\ : IoSpan4Mux
    port map (
            O => \N__19521\,
            I => \N__19518\
        );

    \I__1633\ : IoSpan4Mux
    port map (
            O => \N__19518\,
            I => \N__19515\
        );

    \I__1632\ : Odrv4
    port map (
            O => \N__19515\,
            I => delay_hc_input_ibuf_gb_io_gb_input
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_6\,
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_14\,
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_9_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_22\,
            carryinitout => \bfn_9_12_0_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_30\,
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_2_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_14_0_\
        );

    \IN_MUX_bfv_2_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_acc_cry_7\,
            carryinitout => \bfn_2_15_0_\
        );

    \IN_MUX_bfv_2_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_acc_cry_15\,
            carryinitout => \bfn_2_16_0_\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_12_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_17_0_\
        );

    \IN_MUX_bfv_12_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_12_18_0_\
        );

    \IN_MUX_bfv_12_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_12_19_0_\
        );

    \IN_MUX_bfv_12_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_12_20_0_\
        );

    \IN_MUX_bfv_14_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_21_0_\
        );

    \IN_MUX_bfv_14_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_14_22_0_\
        );

    \IN_MUX_bfv_14_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_14_23_0_\
        );

    \IN_MUX_bfv_14_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_14_24_0_\
        );

    \IN_MUX_bfv_8_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_23_0_\
        );

    \IN_MUX_bfv_8_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_8_24_0_\
        );

    \IN_MUX_bfv_8_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_8_25_0_\
        );

    \IN_MUX_bfv_8_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_8_26_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_17_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s1\,
            carryinitout => \bfn_17_12_0_\
        );

    \IN_MUX_bfv_17_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s1\,
            carryinitout => \bfn_17_13_0_\
        );

    \IN_MUX_bfv_17_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s1\,
            carryinitout => \bfn_17_14_0_\
        );

    \IN_MUX_bfv_15_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_12_0_\
        );

    \IN_MUX_bfv_15_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s0\,
            carryinitout => \bfn_15_13_0_\
        );

    \IN_MUX_bfv_15_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s0\,
            carryinitout => \bfn_15_14_0_\
        );

    \IN_MUX_bfv_15_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s0\,
            carryinitout => \bfn_15_15_0_\
        );

    \IN_MUX_bfv_15_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_8_0_\
        );

    \IN_MUX_bfv_15_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_7\,
            carryinitout => \bfn_15_9_0_\
        );

    \IN_MUX_bfv_15_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_15\,
            carryinitout => \bfn_15_10_0_\
        );

    \IN_MUX_bfv_15_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_23\,
            carryinitout => \bfn_15_11_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\,
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_1_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\,
            carryinitout => \bfn_1_16_0_\
        );

    \IN_MUX_bfv_3_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_15_0_\
        );

    \IN_MUX_bfv_3_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_acc_1_cry_7\,
            carryinitout => \bfn_3_16_0_\
        );

    \IN_MUX_bfv_3_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_acc_1_cry_15\,
            carryinitout => \bfn_3_17_0_\
        );

    \IN_MUX_bfv_3_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_11_0_\
        );

    \IN_MUX_bfv_3_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_3_12_0_\
        );

    \IN_MUX_bfv_2_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_18_0_\
        );

    \IN_MUX_bfv_2_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un19_threshold_acc_cry_7\,
            carryinitout => \bfn_2_19_0_\
        );

    \IN_MUX_bfv_4_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_12_0_\
        );

    \IN_MUX_bfv_4_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_4_13_0_\
        );

    \IN_MUX_bfv_13_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_16_0_\
        );

    \IN_MUX_bfv_13_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un4_running_cry_8\,
            carryinitout => \bfn_13_17_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un4_running_cry_16\,
            carryinitout => \bfn_13_18_0_\
        );

    \IN_MUX_bfv_12_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_14_0_\
        );

    \IN_MUX_bfv_12_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un4_running_cry_8\,
            carryinitout => \bfn_12_15_0_\
        );

    \IN_MUX_bfv_12_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un4_running_cry_16\,
            carryinitout => \bfn_12_16_0_\
        );

    \IN_MUX_bfv_15_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_20_0_\
        );

    \IN_MUX_bfv_15_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un4_running_cry_8\,
            carryinitout => \bfn_15_21_0_\
        );

    \IN_MUX_bfv_15_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un4_running_cry_16\,
            carryinitout => \bfn_15_22_0_\
        );

    \IN_MUX_bfv_9_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_22_0_\
        );

    \IN_MUX_bfv_9_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un4_running_cry_8\,
            carryinitout => \bfn_9_23_0_\
        );

    \IN_MUX_bfv_9_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un4_running_cry_16\,
            carryinitout => \bfn_9_24_0_\
        );

    \IN_MUX_bfv_17_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_19_0_\
        );

    \IN_MUX_bfv_17_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_17_20_0_\
        );

    \IN_MUX_bfv_17_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_17_21_0_\
        );

    \IN_MUX_bfv_17_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_17_22_0_\
        );

    \IN_MUX_bfv_18_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_18_0_\
        );

    \IN_MUX_bfv_18_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_18_19_0_\
        );

    \IN_MUX_bfv_18_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_18_20_0_\
        );

    \IN_MUX_bfv_18_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_18_21_0_\
        );

    \IN_MUX_bfv_10_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_19_0_\
        );

    \IN_MUX_bfv_10_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_10_20_0_\
        );

    \IN_MUX_bfv_10_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_10_21_0_\
        );

    \IN_MUX_bfv_10_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_10_22_0_\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_15_0_\
        );

    \IN_MUX_bfv_8_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_8_16_0_\
        );

    \IN_MUX_bfv_8_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_8_17_0_\
        );

    \IN_MUX_bfv_8_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_8_18_0_\
        );

    \IN_MUX_bfv_13_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_11_0_\
        );

    \IN_MUX_bfv_13_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_7\,
            carryinitout => \bfn_13_12_0_\
        );

    \IN_MUX_bfv_13_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_7_0_\
        );

    \IN_MUX_bfv_13_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_13_8_0_\
        );

    \IN_MUX_bfv_13_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_13_9_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_17_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_7_0_\
        );

    \IN_MUX_bfv_17_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_8\,
            carryinitout => \bfn_17_8_0_\
        );

    \IN_MUX_bfv_17_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_16\,
            carryinitout => \bfn_17_9_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_24\,
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_14_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_5_0_\
        );

    \IN_MUX_bfv_14_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_14_6_0_\
        );

    \IN_MUX_bfv_14_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_14_7_0_\
        );

    \IN_MUX_bfv_14_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_14_8_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\,
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\,
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\,
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_5_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_9_0_\
        );

    \IN_MUX_bfv_5_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryinitout => \bfn_5_10_0_\
        );

    \IN_MUX_bfv_5_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryinitout => \bfn_5_11_0_\
        );

    \IN_MUX_bfv_5_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryinitout => \bfn_5_12_0_\
        );

    \IN_MUX_bfv_12_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_10_0_\
        );

    \IN_MUX_bfv_12_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            carryinitout => \bfn_12_11_0_\
        );

    \delay_tr_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19551\,
            GLOBALBUFFEROUTPUT => delay_tr_input_c_g
        );

    \delay_hc_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19527\,
            GLOBALBUFFEROUTPUT => delay_hc_input_c_g
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__23451\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_hc_timer.N_393_i_g\
        );

    \current_shift_inst.timer_s1.running_RNII51H_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__35826\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_166_i_g\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__32016\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_tr_timer.N_395_i_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__38270\,
            CLKHFEN => \N__38274\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__38283\,
            RGB2PWM => \N__20142\,
            RGB1 => rgb_g_wire,
            CURREN => \N__38236\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__20148\,
            RGB0PWM => \N__48591\,
            RGB0 => rgb_r_wire
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000110010"
        )
    port map (
            in0 => \N__22203\,
            in1 => \N__23097\,
            in2 => \N__22593\,
            in3 => \N__20979\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49251\,
            ce => 'H',
            sr => \N__48464\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__20175\,
            in1 => \N__22737\,
            in2 => \N__20307\,
            in3 => \N__20094\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49251\,
            ce => 'H',
            sr => \N__48464\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__20174\,
            in1 => \N__22758\,
            in2 => \N__20306\,
            in3 => \N__20093\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49251\,
            ce => 'H',
            sr => \N__48464\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000110010"
        )
    port map (
            in0 => \N__22202\,
            in1 => \N__23096\,
            in2 => \N__22632\,
            in3 => \N__20978\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49251\,
            ce => 'H',
            sr => \N__48464\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111111001101"
        )
    port map (
            in0 => \N__20409\,
            in1 => \N__22707\,
            in2 => \N__20304\,
            in3 => \N__22194\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49250\,
            ce => 'H',
            sr => \N__48470\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010100"
        )
    port map (
            in0 => \N__23090\,
            in1 => \N__22854\,
            in2 => \N__22201\,
            in3 => \N__20968\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49250\,
            ce => 'H',
            sr => \N__48470\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110110000"
        )
    port map (
            in0 => \N__20967\,
            in1 => \N__23089\,
            in2 => \N__22923\,
            in3 => \N__22193\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49250\,
            ce => 'H',
            sr => \N__48470\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__20168\,
            in1 => \N__22722\,
            in2 => \N__20305\,
            in3 => \N__20092\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49250\,
            ce => 'H',
            sr => \N__48470\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011110111"
        )
    port map (
            in0 => \N__20966\,
            in1 => \N__20316\,
            in2 => \N__22671\,
            in3 => \N__19611\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49250\,
            ce => 'H',
            sr => \N__48470\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101110"
        )
    port map (
            in0 => \N__22886\,
            in1 => \N__22185\,
            in2 => \N__20977\,
            in3 => \N__23088\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49249\,
            ce => 'H',
            sr => \N__48476\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010101"
        )
    port map (
            in0 => \N__23086\,
            in1 => \N__22664\,
            in2 => \N__20430\,
            in3 => \N__22186\,
            lcout => \current_shift_inst.PI_CTRL.N_149\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23087\,
            lcout => \N_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49247\,
            ce => 'H',
            sr => \N__48497\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__19593\,
            in1 => \N__19602\,
            in2 => \N__21893\,
            in3 => \N__19892\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__19592\,
            in1 => \N__19893\,
            in2 => \_gnd_net_\,
            in3 => \N__21927\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19581\,
            in2 => \N__19569\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_1_14_0_\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19830\,
            in2 => \N__19818\,
            in3 => \N__19800\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19797\,
            in2 => \N__19785\,
            in3 => \N__19767\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19764\,
            in2 => \N__19752\,
            in3 => \N__19737\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19734\,
            in2 => \N__19722\,
            in3 => \N__19704\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19701\,
            in2 => \N__19689\,
            in3 => \N__19674\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19671\,
            in2 => \N__19659\,
            in3 => \N__19644\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19641\,
            in2 => \N__19629\,
            in3 => \N__19614\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20055\,
            in2 => \N__20043\,
            in3 => \N__20025\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\,
            ltout => OPEN,
            carryin => \bfn_1_15_0_\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20022\,
            in2 => \N__20010\,
            in3 => \N__19992\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19989\,
            in2 => \N__19906\,
            in3 => \N__19977\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19897\,
            in2 => \N__19974\,
            in3 => \N__19959\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19956\,
            in2 => \N__19907\,
            in3 => \N__19944\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19901\,
            in2 => \N__19941\,
            in3 => \N__19926\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19923\,
            in2 => \N__19908\,
            in3 => \N__19911\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19905\,
            in2 => \N__19854\,
            in3 => \N__19842\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20613\,
            in1 => \N__19839\,
            in2 => \_gnd_net_\,
            in3 => \N__20151\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__21669\,
            in1 => \N__21686\,
            in2 => \N__20607\,
            in3 => \N__21293\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__22362\,
            in1 => \N__21351\,
            in2 => \N__22392\,
            in3 => \N__21292\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_7_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110111111101"
        )
    port map (
            in0 => \N__22018\,
            in1 => \N__20790\,
            in2 => \N__21939\,
            in3 => \N__21758\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49211\,
            ce => 'H',
            sr => \N__48542\
        );

    \phase_controller_inst1.un7_start_stop_0_a2_LC_1_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__48589\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23621\,
            lcout => un7_start_stop_0_a2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.N_38_i_i_LC_1_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__48590\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23625\,
            lcout => \N_38_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un1_duty_inputlto2_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__20135\,
            in1 => \N__20120\,
            in2 => \_gnd_net_\,
            in3 => \N__20106\,
            lcout => \pwm_generator_inst.un1_duty_inputlt3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000010"
        )
    port map (
            in0 => \N__20408\,
            in1 => \N__22703\,
            in2 => \N__22200\,
            in3 => \N__20286\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20370\,
            in1 => \N__20355\,
            in2 => \N__20078\,
            in3 => \N__20333\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20071\,
            in2 => \_gnd_net_\,
            in3 => \N__20254\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__20369\,
            in1 => \N__20354\,
            in2 => \N__20340\,
            in3 => \N__20332\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22589\,
            in1 => \N__22919\,
            in2 => \N__20988\,
            in3 => \N__22853\,
            lcout => \current_shift_inst.PI_CTRL.N_27\,
            ltout => \current_shift_inst.PI_CTRL.N_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__23067\,
            in1 => \N__20157\,
            in2 => \N__20310\,
            in3 => \N__20952\,
            lcout => \current_shift_inst.PI_CTRL.N_153\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__20200\,
            in1 => \N__20219\,
            in2 => \N__20265\,
            in3 => \N__20235\,
            lcout => \pwm_generator_inst.N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101011"
        )
    port map (
            in0 => \N__20229\,
            in1 => \N__20220\,
            in2 => \N__20205\,
            in3 => \N__20184\,
            lcout => \pwm_generator_inst.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__23068\,
            in1 => \_gnd_net_\,
            in2 => \N__20429\,
            in3 => \N__22184\,
            lcout => \current_shift_inst.PI_CTRL.N_154\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22656\,
            in2 => \_gnd_net_\,
            in3 => \N__22702\,
            lcout => \current_shift_inst.PI_CTRL.N_155\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22846\,
            in2 => \_gnd_net_\,
            in3 => \N__22625\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__22918\,
            in1 => \N__22585\,
            in2 => \N__20433\,
            in3 => \N__22887\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => \current_shift_inst.PI_CTRL.N_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110101"
        )
    port map (
            in0 => \N__22657\,
            in1 => \_gnd_net_\,
            in2 => \N__20412\,
            in3 => \N__23066\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_2_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__21986\,
            in1 => \N__21852\,
            in2 => \N__20649\,
            in3 => \N__21724\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49245\,
            ce => 'H',
            sr => \N__48498\
        );

    \pwm_generator_inst.threshold_ACC_3_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__21725\,
            in1 => \N__21987\,
            in2 => \N__21911\,
            in3 => \N__20859\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49245\,
            ce => 'H',
            sr => \N__48498\
        );

    \pwm_generator_inst.threshold_ACC_1_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111000111111101"
        )
    port map (
            in0 => \N__21985\,
            in1 => \N__21851\,
            in2 => \N__20670\,
            in3 => \N__21723\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49245\,
            ce => 'H',
            sr => \N__48498\
        );

    \pwm_generator_inst.threshold_7_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20394\,
            lcout => \pwm_generator_inst.thresholdZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49241\,
            ce => 'H',
            sr => \N__48506\
        );

    \pwm_generator_inst.threshold_6_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20382\,
            lcout => \pwm_generator_inst.thresholdZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49237\,
            ce => 'H',
            sr => \N__48516\
        );

    \pwm_generator_inst.threshold_ACC_6_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111000111111101"
        )
    port map (
            in0 => \N__21988\,
            in1 => \N__21943\,
            in2 => \N__20814\,
            in3 => \N__21740\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49237\,
            ce => 'H',
            sr => \N__48516\
        );

    \pwm_generator_inst.threshold_4_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20376\,
            lcout => \pwm_generator_inst.thresholdZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49233\,
            ce => 'H',
            sr => \N__48522\
        );

    \pwm_generator_inst.threshold_ACC_4_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__21741\,
            in1 => \N__21989\,
            in2 => \N__21950\,
            in3 => \N__20841\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49233\,
            ce => 'H',
            sr => \N__48522\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21251\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_14_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20529\,
            in2 => \_gnd_net_\,
            in3 => \N__20514\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20511\,
            in2 => \_gnd_net_\,
            in3 => \N__20496\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20493\,
            in2 => \_gnd_net_\,
            in3 => \N__20481\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20478\,
            in2 => \_gnd_net_\,
            in3 => \N__20472\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38198\,
            in2 => \N__20469\,
            in3 => \N__20460\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38200\,
            in2 => \N__20457\,
            in3 => \N__20448\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38199\,
            in2 => \N__20445\,
            in3 => \N__20436\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20586\,
            in2 => \_gnd_net_\,
            in3 => \N__20580\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_2_15_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20577\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20571\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20565\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20559\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20553\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20547\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20541\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20535\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_16_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20634\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20628\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20622\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20616\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__21527\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20759\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__21687\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20600\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__21653\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20690\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001110010"
        )
    port map (
            in0 => \N__21294\,
            in1 => \N__21600\,
            in2 => \N__21207\,
            in3 => \N__21624\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20735\,
            in1 => \N__21591\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_15\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011110000010"
        )
    port map (
            in0 => \N__21296\,
            in1 => \N__21579\,
            in2 => \N__20739\,
            in3 => \N__20736\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21570\,
            in2 => \_gnd_net_\,
            in3 => \N__20723\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_16\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__20724\,
            in1 => \N__21558\,
            in2 => \N__20712\,
            in3 => \N__21322\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__21549\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20708\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_17\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__20709\,
            in1 => \N__21323\,
            in2 => \N__20697\,
            in3 => \N__21537\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__21654\,
            in1 => \N__21633\,
            in2 => \N__20694\,
            in3 => \N__21295\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20676\,
            in2 => \N__21335\,
            in3 => \N__21331\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_2_18_0_\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21231\,
            in2 => \_gnd_net_\,
            in3 => \N__20658\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_0\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20655\,
            in2 => \_gnd_net_\,
            in3 => \N__20637\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_1\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20865\,
            in2 => \_gnd_net_\,
            in3 => \N__20850\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_2\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20847\,
            in2 => \_gnd_net_\,
            in3 => \N__20832\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_3\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20829\,
            in2 => \_gnd_net_\,
            in3 => \N__20823\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_4\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20820\,
            in2 => \_gnd_net_\,
            in3 => \N__20799\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_5\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20796\,
            in2 => \_gnd_net_\,
            in3 => \N__20784\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_6\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20745\,
            in2 => \_gnd_net_\,
            in3 => \N__20781\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_2_19_0_\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010101101010"
        )
    port map (
            in0 => \N__20778\,
            in1 => \N__21492\,
            in2 => \N__21336\,
            in3 => \N__20769\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100001110100"
        )
    port map (
            in0 => \N__21528\,
            in1 => \N__21327\,
            in2 => \N__20766\,
            in3 => \N__21507\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_3_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22885\,
            in2 => \_gnd_net_\,
            in3 => \N__22624\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22125\,
            in1 => \N__22212\,
            in2 => \N__22326\,
            in3 => \N__22110\,
            lcout => \current_shift_inst.PI_CTRL.N_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_1_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20925\,
            lcout => \pwm_generator_inst.thresholdZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49242\,
            ce => 'H',
            sr => \N__48484\
        );

    \pwm_generator_inst.threshold_3_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20919\,
            lcout => \pwm_generator_inst.thresholdZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49242\,
            ce => 'H',
            sr => \N__48484\
        );

    \pwm_generator_inst.threshold_2_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20913\,
            lcout => \pwm_generator_inst.thresholdZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49242\,
            ce => 'H',
            sr => \N__48484\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22077\,
            in2 => \N__20907\,
            in3 => \N__22298\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_3_11_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20898\,
            in2 => \N__20892\,
            in3 => \N__22276\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20883\,
            in2 => \N__20874\,
            in3 => \N__22256\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21102\,
            in2 => \N__21096\,
            in3 => \N__22234\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21087\,
            in2 => \N__21078\,
            in3 => \N__22555\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22092\,
            in2 => \N__21069\,
            in3 => \N__22534\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21051\,
            in2 => \N__21060\,
            in3 => \N__22513\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22492\,
            in1 => \N__21045\,
            in2 => \N__21036\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22029\,
            in2 => \N__21027\,
            in3 => \N__22472\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_3_12_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21018\,
            in2 => \N__22053\,
            in3 => \N__22408\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21012\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49234\,
            ce => 'H',
            sr => \N__48507\
        );

    \pwm_generator_inst.counter_RNISQD2_0_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22255\,
            in2 => \_gnd_net_\,
            in3 => \N__22297\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIBO26_1_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__22556\,
            in1 => \N__22235\,
            in2 => \N__21219\,
            in3 => \N__22277\,
            lcout => \pwm_generator_inst.un1_counterlt9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIVDL3_9_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__22493\,
            in1 => \N__22471\,
            in2 => \_gnd_net_\,
            in3 => \N__22409\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto9_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_5_LC_3_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__22515\,
            in1 => \N__22536\,
            in2 => \N__21216\,
            in3 => \N__21213\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21197\,
            in2 => \_gnd_net_\,
            in3 => \N__21619\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21168\,
            in2 => \_gnd_net_\,
            in3 => \N__21186\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_3_15_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21147\,
            in2 => \_gnd_net_\,
            in3 => \N__21162\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_0\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21129\,
            in2 => \_gnd_net_\,
            in3 => \N__21141\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_1\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21108\,
            in2 => \_gnd_net_\,
            in3 => \N__21123\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_2\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21468\,
            in2 => \_gnd_net_\,
            in3 => \N__21483\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_3\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21450\,
            in2 => \_gnd_net_\,
            in3 => \N__21462\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_4\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21426\,
            in2 => \_gnd_net_\,
            in3 => \N__21444\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_5\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21402\,
            in2 => \_gnd_net_\,
            in3 => \N__21420\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_6\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21378\,
            in2 => \_gnd_net_\,
            in3 => \N__21396\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_3_16_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21357\,
            in2 => \_gnd_net_\,
            in3 => \N__21372\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_8\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22357\,
            in2 => \_gnd_net_\,
            in3 => \N__21339\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_9\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__21312\,
            in1 => \N__21255\,
            in2 => \_gnd_net_\,
            in3 => \N__21222\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_10\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21685\,
            in2 => \_gnd_net_\,
            in3 => \N__21657\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_11\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21649\,
            in2 => \_gnd_net_\,
            in3 => \N__21627\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_12\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21620\,
            in2 => \_gnd_net_\,
            in3 => \N__21594\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_13\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21590\,
            in2 => \_gnd_net_\,
            in3 => \N__21573\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_14\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21569\,
            in2 => \_gnd_net_\,
            in3 => \N__21552\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_3_17_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21548\,
            in2 => \_gnd_net_\,
            in3 => \N__21531\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_16\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21526\,
            in2 => \_gnd_net_\,
            in3 => \N__21498\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_17\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21495\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_0_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__22008\,
            in1 => \N__22098\,
            in2 => \N__21948\,
            in3 => \N__21761\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49200\,
            ce => 'H',
            sr => \N__48538\
        );

    \pwm_generator_inst.threshold_5_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22059\,
            lcout => \pwm_generator_inst.thresholdZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49200\,
            ce => 'H',
            sr => \N__48538\
        );

    \pwm_generator_inst.threshold_0_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22083\,
            lcout => \pwm_generator_inst.thresholdZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49200\,
            ce => 'H',
            sr => \N__48538\
        );

    \pwm_generator_inst.threshold_ACC_5_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__22009\,
            in1 => \N__22065\,
            in2 => \N__21949\,
            in3 => \N__21762\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49200\,
            ce => 'H',
            sr => \N__48538\
        );

    \pwm_generator_inst.threshold_9_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22035\,
            lcout => \pwm_generator_inst.thresholdZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49196\,
            ce => 'H',
            sr => \N__48540\
        );

    \pwm_generator_inst.threshold_ACC_9_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__21760\,
            in1 => \N__22041\,
            in2 => \N__21951\,
            in3 => \N__22020\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49196\,
            ce => 'H',
            sr => \N__48540\
        );

    \pwm_generator_inst.threshold_8_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21693\,
            lcout => \pwm_generator_inst.thresholdZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49196\,
            ce => 'H',
            sr => \N__48540\
        );

    \pwm_generator_inst.threshold_ACC_8_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111000111111101"
        )
    port map (
            in0 => \N__22019\,
            in1 => \N__21947\,
            in2 => \N__21771\,
            in3 => \N__21759\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49196\,
            ce => 'H',
            sr => \N__48540\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__23033\,
            in1 => \N__23018\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23204\,
            in1 => \N__23184\,
            in2 => \N__22215\,
            in3 => \N__22944\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22812\,
            in1 => \N__22104\,
            in2 => \N__22797\,
            in3 => \N__23385\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22332\,
            in1 => \N__22314\,
            in2 => \N__22206\,
            in3 => \N__22305\,
            lcout => \current_shift_inst.PI_CTRL.N_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22781\,
            in1 => \N__22973\,
            in2 => \N__22992\,
            in3 => \N__22769\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22793\,
            in2 => \_gnd_net_\,
            in3 => \N__22823\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23240\,
            in1 => \N__23126\,
            in2 => \N__23228\,
            in3 => \N__22958\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23151\,
            in1 => \N__22811\,
            in2 => \N__22119\,
            in3 => \N__22116\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22824\,
            in1 => \N__23127\,
            in2 => \N__23019\,
            in3 => \N__23034\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22770\,
            in1 => \N__22782\,
            in2 => \N__23229\,
            in3 => \N__23241\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23165\,
            in1 => \N__23414\,
            in2 => \N__23403\,
            in3 => \N__23112\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22974\,
            in1 => \N__23183\,
            in2 => \N__23205\,
            in3 => \N__22991\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__23166\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23111\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23150\,
            in1 => \N__22943\,
            in2 => \N__22308\,
            in3 => \N__22959\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_0_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22449\,
            in1 => \N__22299\,
            in2 => \_gnd_net_\,
            in3 => \N__22281\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_4_12_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__49228\,
            ce => 'H',
            sr => \N__48499\
        );

    \pwm_generator_inst.counter_1_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22443\,
            in1 => \N__22278\,
            in2 => \_gnd_net_\,
            in3 => \N__22260\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__49228\,
            ce => 'H',
            sr => \N__48499\
        );

    \pwm_generator_inst.counter_2_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22450\,
            in1 => \N__22257\,
            in2 => \_gnd_net_\,
            in3 => \N__22239\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__49228\,
            ce => 'H',
            sr => \N__48499\
        );

    \pwm_generator_inst.counter_3_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22444\,
            in1 => \N__22236\,
            in2 => \_gnd_net_\,
            in3 => \N__22218\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__49228\,
            ce => 'H',
            sr => \N__48499\
        );

    \pwm_generator_inst.counter_4_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22451\,
            in1 => \N__22557\,
            in2 => \_gnd_net_\,
            in3 => \N__22539\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__49228\,
            ce => 'H',
            sr => \N__48499\
        );

    \pwm_generator_inst.counter_5_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22445\,
            in1 => \N__22535\,
            in2 => \_gnd_net_\,
            in3 => \N__22518\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__49228\,
            ce => 'H',
            sr => \N__48499\
        );

    \pwm_generator_inst.counter_6_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22452\,
            in1 => \N__22514\,
            in2 => \_gnd_net_\,
            in3 => \N__22497\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__49228\,
            ce => 'H',
            sr => \N__48499\
        );

    \pwm_generator_inst.counter_7_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22446\,
            in1 => \N__22494\,
            in2 => \_gnd_net_\,
            in3 => \N__22476\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__49228\,
            ce => 'H',
            sr => \N__48499\
        );

    \pwm_generator_inst.counter_8_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22448\,
            in1 => \N__22473\,
            in2 => \_gnd_net_\,
            in3 => \N__22455\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_4_13_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__49222\,
            ce => 'H',
            sr => \N__48508\
        );

    \pwm_generator_inst.counter_9_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__22410\,
            in1 => \N__22447\,
            in2 => \_gnd_net_\,
            in3 => \N__22413\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49222\,
            ce => 'H',
            sr => \N__48508\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__22361\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22385\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_LC_4_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__33234\,
            in1 => \N__30126\,
            in2 => \_gnd_net_\,
            in3 => \N__33035\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49201\,
            ce => \N__32889\,
            sr => \N__48533\
        );

    \SB_DFF_inst_PH2_MAX_D1_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22341\,
            lcout => \il_max_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49248\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_1_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32460\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49246\,
            ce => 'H',
            sr => \N__48436\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI967M_0_13_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23941\,
            in1 => \N__28999\,
            in2 => \N__31907\,
            in3 => \N__29813\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23337\,
            in2 => \N__26214\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_5_9_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            clk => \N__49238\,
            ce => 'H',
            sr => \N__48465\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22746\,
            in2 => \N__32112\,
            in3 => \N__22725\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            clk => \N__49238\,
            ce => 'H',
            sr => \N__48465\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28938\,
            in2 => \N__23328\,
            in3 => \N__22710\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            clk => \N__49238\,
            ce => 'H',
            sr => \N__48465\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23316\,
            in2 => \N__26028\,
            in3 => \N__22674\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            clk => \N__49238\,
            ce => 'H',
            sr => \N__48465\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26510\,
            in2 => \N__23307\,
            in3 => \N__22635\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__49238\,
            ce => 'H',
            sr => \N__48465\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23358\,
            in2 => \N__23805\,
            in3 => \N__22596\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__49238\,
            ce => 'H',
            sr => \N__48465\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23346\,
            in2 => \N__26760\,
            in3 => \N__22926\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__49238\,
            ce => 'H',
            sr => \N__48465\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23430\,
            in2 => \N__23733\,
            in3 => \N__22890\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__49238\,
            ce => 'H',
            sr => \N__48465\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33366\,
            in2 => \N__26172\,
            in3 => \N__22857\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_5_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__49235\,
            ce => 'H',
            sr => \N__48471\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23286\,
            in2 => \N__26301\,
            in3 => \N__22827\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__49235\,
            ce => 'H',
            sr => \N__48471\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27027\,
            in2 => \N__23277\,
            in3 => \N__22815\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__49235\,
            ce => 'H',
            sr => \N__48471\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23295\,
            in2 => \N__37899\,
            in3 => \N__22800\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__49235\,
            ce => 'H',
            sr => \N__48471\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24462\,
            in2 => \N__32175\,
            in3 => \N__22785\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__49235\,
            ce => 'H',
            sr => \N__48471\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31908\,
            in2 => \N__23958\,
            in3 => \N__22773\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__49235\,
            ce => 'H',
            sr => \N__48471\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23823\,
            in2 => \N__29004\,
            in3 => \N__22761\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__49235\,
            ce => 'H',
            sr => \N__48471\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26357\,
            in2 => \N__23861\,
            in3 => \N__23022\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__49235\,
            ce => 'H',
            sr => \N__48471\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23862\,
            in2 => \N__23946\,
            in3 => \N__23001\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_5_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__49229\,
            ce => 'H',
            sr => \N__48477\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32328\,
            in2 => \N__23892\,
            in3 => \N__22998\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__49229\,
            ce => 'H',
            sr => \N__48477\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23866\,
            in2 => \N__32271\,
            in3 => \N__22995\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__49229\,
            ce => 'H',
            sr => \N__48477\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26421\,
            in2 => \N__23893\,
            in3 => \N__22977\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__49229\,
            ce => 'H',
            sr => \N__48477\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23870\,
            in2 => \N__26850\,
            in3 => \N__22962\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__49229\,
            ce => 'H',
            sr => \N__48477\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26898\,
            in2 => \N__23894\,
            in3 => \N__22947\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__49229\,
            ce => 'H',
            sr => \N__48477\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23874\,
            in2 => \N__31848\,
            in3 => \N__22929\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__49229\,
            ce => 'H',
            sr => \N__48477\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29814\,
            in2 => \N__23895\,
            in3 => \N__23232\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__49229\,
            ce => 'H',
            sr => \N__48477\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23878\,
            in2 => \N__26567\,
            in3 => \N__23208\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_5_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__49223\,
            ce => 'H',
            sr => \N__48485\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44741\,
            in2 => \N__23896\,
            in3 => \N__23187\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__49223\,
            ce => 'H',
            sr => \N__48485\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23882\,
            in2 => \N__40073\,
            in3 => \N__23169\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__49223\,
            ce => 'H',
            sr => \N__48485\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31970\,
            in2 => \N__23897\,
            in3 => \N__23154\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__49223\,
            ce => 'H',
            sr => \N__48485\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23886\,
            in2 => \N__29223\,
            in3 => \N__23130\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__49223\,
            ce => 'H',
            sr => \N__48485\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40314\,
            in2 => \N__23898\,
            in3 => \N__23115\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__49223\,
            ce => 'H',
            sr => \N__48485\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23890\,
            in2 => \N__26691\,
            in3 => \N__23103\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__49223\,
            ce => 'H',
            sr => \N__48485\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__23891\,
            in1 => \_gnd_net_\,
            in2 => \N__27357\,
            in3 => \N__23100\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49223\,
            ce => 'H',
            sr => \N__48485\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29651\,
            in2 => \_gnd_net_\,
            in3 => \N__44594\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44595\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29597\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D2_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23265\,
            lcout => \il_max_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49213\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_hc_RNO_1_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24560\,
            in2 => \_gnd_net_\,
            in3 => \N__23503\,
            lcout => \phase_controller_inst2.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D1_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23253\,
            lcout => \il_min_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49239\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29805\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26166\,
            in1 => \N__23725\,
            in2 => \N__26755\,
            in3 => \N__26291\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__26509\,
            in1 => \N__26024\,
            in2 => \N__23244\,
            in3 => \N__23801\,
            lcout => \current_shift_inst.PI_CTRL.N_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI654B_29_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40318\,
            in2 => \_gnd_net_\,
            in3 => \N__27022\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32358\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49230\,
            ce => 'H',
            sr => \N__48448\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32685\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49230\,
            ce => 'H',
            sr => \N__48448\
        );

    \current_shift_inst.PI_CTRL.prop_term_0_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36840\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49230\,
            ce => 'H',
            sr => \N__48448\
        );

    \current_shift_inst.PI_CTRL.prop_term_2_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32436\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49230\,
            ce => 'H',
            sr => \N__48448\
        );

    \current_shift_inst.PI_CTRL.prop_term_3_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32412\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49230\,
            ce => 'H',
            sr => \N__48448\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32388\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49230\,
            ce => 'H',
            sr => \N__48448\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32612\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49224\,
            ce => 'H',
            sr => \N__48458\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33351\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49224\,
            ce => 'H',
            sr => \N__48458\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33447\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49224\,
            ce => 'H',
            sr => \N__48458\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110011111110"
        )
    port map (
            in0 => \N__27515\,
            in1 => \N__27355\,
            in2 => \N__27198\,
            in3 => \N__24747\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49224\,
            ce => 'H',
            sr => \N__48458\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32654\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49224\,
            ce => 'H',
            sr => \N__48458\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26416\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26338\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23418\,
            in2 => \_gnd_net_\,
            in3 => \N__23399\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23921\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D2_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23373\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_min_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26546\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_tr_RNO_0_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23558\,
            in2 => \_gnd_net_\,
            in3 => \N__23477\,
            lcout => \phase_controller_inst2.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_tr_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__35407\,
            in1 => \N__23987\,
            in2 => \N__34958\,
            in3 => \N__23364\,
            lcout => \phase_controller_inst2.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49206\,
            ce => 'H',
            sr => \N__48478\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__24029\,
            in1 => \N__24052\,
            in2 => \_gnd_net_\,
            in3 => \N__24507\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49206\,
            ce => 'H',
            sr => \N__48478\
        );

    \phase_controller_inst2.state_1_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__23483\,
            in1 => \N__23466\,
            in2 => \N__29961\,
            in3 => \N__23553\,
            lcout => \phase_controller_inst2.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49202\,
            ce => 'H',
            sr => \N__48486\
        );

    \phase_controller_inst2.state_2_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010001000100"
        )
    port map (
            in0 => \N__29960\,
            in1 => \N__23465\,
            in2 => \N__24559\,
            in3 => \N__23504\,
            lcout => \phase_controller_inst2.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49202\,
            ce => 'H',
            sr => \N__48486\
        );

    \phase_controller_inst2.state_3_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__23988\,
            in1 => \N__23505\,
            in2 => \N__24558\,
            in3 => \N__31683\,
            lcout => \phase_controller_inst2.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49202\,
            ce => 'H',
            sr => \N__48486\
        );

    \phase_controller_inst2.state_0_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__23554\,
            in1 => \N__34986\,
            in2 => \N__24003\,
            in3 => \N__23484\,
            lcout => \phase_controller_inst2.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49202\,
            ce => 'H',
            sr => \N__48486\
        );

    \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__23643\,
            in1 => \N__30432\,
            in2 => \_gnd_net_\,
            in3 => \N__29982\,
            lcout => \phase_controller_inst2.stoper_hc.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24054\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34929\,
            in2 => \_gnd_net_\,
            in3 => \N__34957\,
            lcout => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_hc_RNO_0_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__29951\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23464\,
            lcout => \phase_controller_inst2.start_timer_hc_RNO_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24053\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24030\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_393_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_hc_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__35400\,
            in1 => \N__23664\,
            in2 => \N__23649\,
            in3 => \N__23658\,
            lcout => \phase_controller_inst2.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49189\,
            ce => 'H',
            sr => \N__48509\
        );

    \phase_controller_inst2.stoper_hc.start_latched_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23645\,
            lcout => \phase_controller_inst2.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49189\,
            ce => 'H',
            sr => \N__48509\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30433\,
            in2 => \_gnd_net_\,
            in3 => \N__23644\,
            lcout => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_4_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__23608\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35396\,
            lcout => phase_controller_inst1_state_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49153\,
            ce => 'H',
            sr => \N__48537\
        );

    \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31717\,
            in2 => \_gnd_net_\,
            in3 => \N__31649\,
            lcout => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_ns_i_a2_1_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23609\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35383\,
            lcout => state_ns_i_a2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.S2_LC_7_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23562\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49131\,
            ce => 'H',
            sr => \N__48544\
        );

    \SB_DFF_inst_PH1_MAX_D1_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23520\,
            lcout => \il_max_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49243\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D2_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23511\,
            lcout => \il_max_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49243\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_hc_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24496\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24473\,
            ce => 'H',
            sr => \N__48416\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFE9M_18_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32258\,
            in1 => \N__31836\,
            in2 => \N__26420\,
            in3 => \N__27316\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__23797\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23729\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI967M_13_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23942\,
            in1 => \N__31886\,
            in2 => \N__29003\,
            in3 => \N__29806\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIMJHC1_28_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29222\,
            in1 => \N__23676\,
            in2 => \N__23697\,
            in3 => \N__31961\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIHF8M_18_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26553\,
            in1 => \N__31835\,
            in2 => \N__32266\,
            in3 => \N__26411\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNID8UD2_11_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23682\,
            in1 => \N__23670\,
            in2 => \N__23694\,
            in3 => \N__23691\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__40049\,
            in1 => \N__44732\,
            in2 => \N__29221\,
            in3 => \N__26891\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI005B_30_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26690\,
            in2 => \_gnd_net_\,
            in3 => \N__32153\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26831\,
            in1 => \N__26349\,
            in2 => \N__32322\,
            in3 => \N__37881\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26554\,
            in1 => \N__44733\,
            in2 => \N__40062\,
            in3 => \N__26892\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI24CN6_18_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23763\,
            in1 => \N__23757\,
            in2 => \N__23751\,
            in3 => \N__23739\,
            lcout => \current_shift_inst.PI_CTRL.N_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26350\,
            in1 => \N__26832\,
            in2 => \N__37891\,
            in3 => \N__32312\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIHL6U3_29_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27026\,
            in1 => \N__40319\,
            in2 => \N__23748\,
            in3 => \N__23745\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIISQ01_11_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__23721\,
            in1 => \N__44575\,
            in2 => \N__32613\,
            in3 => \N__29292\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIISQ01Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23720\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000111110101"
        )
    port map (
            in0 => \N__27317\,
            in1 => \N__27502\,
            in2 => \N__27176\,
            in3 => \N__24603\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49225\,
            ce => 'H',
            sr => \N__48437\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__27501\,
            in1 => \N__27318\,
            in2 => \N__24951\,
            in3 => \N__27132\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49225\,
            ce => 'H',
            sr => \N__48437\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110100011101"
        )
    port map (
            in0 => \N__27369\,
            in1 => \N__27169\,
            in2 => \N__24855\,
            in3 => \N__27514\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49220\,
            ce => 'H',
            sr => \N__48449\
        );

    \current_shift_inst.PI_CTRL.error_control_RNICIJ3_13_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32539\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_13_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32540\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49220\,
            ce => 'H',
            sr => \N__48449\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__29459\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44515\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\,
            ltout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6I_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111110101"
        )
    port map (
            in0 => \N__44516\,
            in1 => \N__23931\,
            in2 => \N__23901\,
            in3 => \N__29445\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_14_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44517\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49220\,
            ce => 'H',
            sr => \N__48449\
        );

    \current_shift_inst.PI_CTRL.error_control_RNILF8U_9_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__23787\,
            in1 => \N__33347\,
            in2 => \N__44590\,
            in3 => \N__29322\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNILF8UZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23786\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000110111011"
        )
    port map (
            in0 => \N__27165\,
            in1 => \N__27314\,
            in2 => \N__27524\,
            in3 => \N__24633\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49214\,
            ce => 'H',
            sr => \N__48459\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010111100101110"
        )
    port map (
            in0 => \N__27311\,
            in1 => \N__27167\,
            in2 => \N__24867\,
            in3 => \N__27512\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49214\,
            ce => 'H',
            sr => \N__48459\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011111110"
        )
    port map (
            in0 => \N__27164\,
            in1 => \N__27313\,
            in2 => \N__27523\,
            in3 => \N__25038\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49214\,
            ce => 'H',
            sr => \N__48459\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010111100101110"
        )
    port map (
            in0 => \N__27312\,
            in1 => \N__27168\,
            in2 => \N__25029\,
            in3 => \N__27513\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49214\,
            ce => 'H',
            sr => \N__48459\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000110111"
        )
    port map (
            in0 => \N__27166\,
            in1 => \N__24588\,
            in2 => \N__27525\,
            in3 => \N__27315\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49214\,
            ce => 'H',
            sr => \N__48459\
        );

    \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26142\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__27516\,
            in1 => \N__27351\,
            in2 => \N__24777\,
            in3 => \N__27160\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49207\,
            ce => 'H',
            sr => \N__48466\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011111110"
        )
    port map (
            in0 => \N__27350\,
            in1 => \N__27522\,
            in2 => \N__27191\,
            in3 => \N__24900\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49207\,
            ce => 'H',
            sr => \N__48466\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__27518\,
            in1 => \N__27353\,
            in2 => \N__24879\,
            in3 => \N__27162\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49207\,
            ce => 'H',
            sr => \N__48466\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011111110"
        )
    port map (
            in0 => \N__27349\,
            in1 => \N__27521\,
            in2 => \N__27190\,
            in3 => \N__24924\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49207\,
            ce => 'H',
            sr => \N__48466\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__27517\,
            in1 => \N__27352\,
            in2 => \N__24936\,
            in3 => \N__27161\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49207\,
            ce => 'H',
            sr => \N__48466\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011111110"
        )
    port map (
            in0 => \N__27348\,
            in1 => \N__27520\,
            in2 => \N__27189\,
            in3 => \N__24984\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49207\,
            ce => 'H',
            sr => \N__48466\
        );

    \current_shift_inst.PI_CTRL.integrator_31_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__27519\,
            in1 => \N__27354\,
            in2 => \N__25002\,
            in3 => \N__27163\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49207\,
            ce => 'H',
            sr => \N__48466\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__24503\,
            in1 => \N__24051\,
            in2 => \_gnd_net_\,
            in3 => \N__24028\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_394_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9A0221_17_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011000"
        )
    port map (
            in0 => \N__31128\,
            in1 => \N__30786\,
            in2 => \N__29091\,
            in3 => \N__47699\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_RNI9M3O_0_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34985\,
            in2 => \_gnd_net_\,
            in3 => \N__23999\,
            lcout => \phase_controller_inst2.state_RNI9M3OZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24267\,
            in1 => \N__28042\,
            in2 => \_gnd_net_\,
            in3 => \N__23976\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_15_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__49190\,
            ce => \N__24145\,
            sr => \N__48487\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24241\,
            in1 => \N__27989\,
            in2 => \_gnd_net_\,
            in3 => \N__23973\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__49190\,
            ce => \N__24145\,
            sr => \N__48487\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24268\,
            in1 => \N__27937\,
            in2 => \_gnd_net_\,
            in3 => \N__23970\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__49190\,
            ce => \N__24145\,
            sr => \N__48487\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24242\,
            in1 => \N__27878\,
            in2 => \_gnd_net_\,
            in3 => \N__23967\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__49190\,
            ce => \N__24145\,
            sr => \N__48487\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24269\,
            in1 => \N__27824\,
            in2 => \_gnd_net_\,
            in3 => \N__23964\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__49190\,
            ce => \N__24145\,
            sr => \N__48487\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24243\,
            in1 => \N__28336\,
            in2 => \_gnd_net_\,
            in3 => \N__23961\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__49190\,
            ce => \N__24145\,
            sr => \N__48487\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24270\,
            in1 => \N__28310\,
            in2 => \_gnd_net_\,
            in3 => \N__24081\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__49190\,
            ce => \N__24145\,
            sr => \N__48487\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24244\,
            in1 => \N__28291\,
            in2 => \_gnd_net_\,
            in3 => \N__24078\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__49190\,
            ce => \N__24145\,
            sr => \N__48487\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24248\,
            in1 => \N__28255\,
            in2 => \_gnd_net_\,
            in3 => \N__24075\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_16_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__49182\,
            ce => \N__24144\,
            sr => \N__48500\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24252\,
            in1 => \N__28225\,
            in2 => \_gnd_net_\,
            in3 => \N__24072\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__49182\,
            ce => \N__24144\,
            sr => \N__48500\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24245\,
            in1 => \N__28189\,
            in2 => \_gnd_net_\,
            in3 => \N__24069\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__49182\,
            ce => \N__24144\,
            sr => \N__48500\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24249\,
            in1 => \N__28154\,
            in2 => \_gnd_net_\,
            in3 => \N__24066\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__49182\,
            ce => \N__24144\,
            sr => \N__48500\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24246\,
            in1 => \N__28130\,
            in2 => \_gnd_net_\,
            in3 => \N__24063\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__49182\,
            ce => \N__24144\,
            sr => \N__48500\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24250\,
            in1 => \N__28100\,
            in2 => \_gnd_net_\,
            in3 => \N__24060\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__49182\,
            ce => \N__24144\,
            sr => \N__48500\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24247\,
            in1 => \N__28571\,
            in2 => \_gnd_net_\,
            in3 => \N__24057\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__49182\,
            ce => \N__24144\,
            sr => \N__48500\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24251\,
            in1 => \N__28537\,
            in2 => \_gnd_net_\,
            in3 => \N__24108\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__49182\,
            ce => \N__24144\,
            sr => \N__48500\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24263\,
            in1 => \N__28507\,
            in2 => \_gnd_net_\,
            in3 => \N__24105\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_8_17_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__49174\,
            ce => \N__24146\,
            sr => \N__48510\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24253\,
            in1 => \N__28480\,
            in2 => \_gnd_net_\,
            in3 => \N__24102\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__49174\,
            ce => \N__24146\,
            sr => \N__48510\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24264\,
            in1 => \N__28459\,
            in2 => \_gnd_net_\,
            in3 => \N__24099\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__49174\,
            ce => \N__24146\,
            sr => \N__48510\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24254\,
            in1 => \N__28429\,
            in2 => \_gnd_net_\,
            in3 => \N__24096\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__49174\,
            ce => \N__24146\,
            sr => \N__48510\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24265\,
            in1 => \N__28394\,
            in2 => \_gnd_net_\,
            in3 => \N__24093\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__49174\,
            ce => \N__24146\,
            sr => \N__48510\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24255\,
            in1 => \N__28366\,
            in2 => \_gnd_net_\,
            in3 => \N__24090\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__49174\,
            ce => \N__24146\,
            sr => \N__48510\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24266\,
            in1 => \N__28883\,
            in2 => \_gnd_net_\,
            in3 => \N__24087\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__49174\,
            ce => \N__24146\,
            sr => \N__48510\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24256\,
            in1 => \N__28859\,
            in2 => \_gnd_net_\,
            in3 => \N__24084\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__49174\,
            ce => \N__24146\,
            sr => \N__48510\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24257\,
            in1 => \N__28828\,
            in2 => \_gnd_net_\,
            in3 => \N__24285\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_8_18_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__49167\,
            ce => \N__24150\,
            sr => \N__48517\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24261\,
            in1 => \N__28775\,
            in2 => \_gnd_net_\,
            in3 => \N__24282\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__49167\,
            ce => \N__24150\,
            sr => \N__48517\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24258\,
            in1 => \N__28735\,
            in2 => \_gnd_net_\,
            in3 => \N__24279\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__49167\,
            ce => \N__24150\,
            sr => \N__48517\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24262\,
            in1 => \N__28658\,
            in2 => \_gnd_net_\,
            in3 => \N__24276\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__49167\,
            ce => \N__24150\,
            sr => \N__48517\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24259\,
            in1 => \N__28709\,
            in2 => \_gnd_net_\,
            in3 => \N__24273\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__49167\,
            ce => \N__24150\,
            sr => \N__48517\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__28688\,
            in1 => \N__24260\,
            in2 => \_gnd_net_\,
            in3 => \N__24153\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49167\,
            ce => \N__24150\,
            sr => \N__48517\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28053\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49159\,
            ce => \N__28620\,
            sr => \N__48523\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101000011001100"
        )
    port map (
            in0 => \N__25689\,
            in1 => \N__31558\,
            in2 => \N__31722\,
            in3 => \N__24339\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49154\,
            ce => 'H',
            sr => \N__48528\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__24334\,
            in1 => \N__24351\,
            in2 => \N__25203\,
            in3 => \N__32765\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49148\,
            ce => 'H',
            sr => \N__48534\
        );

    \phase_controller_inst1.stoper_hc.running_LC_8_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111110000"
        )
    port map (
            in0 => \N__31718\,
            in1 => \N__25688\,
            in2 => \N__24366\,
            in3 => \N__24335\,
            lcout => \phase_controller_inst1.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49148\,
            ce => 'H',
            sr => \N__48534\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_8_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24332\,
            in2 => \_gnd_net_\,
            in3 => \N__24350\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_8_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__31706\,
            in1 => \N__24362\,
            in2 => \_gnd_net_\,
            in3 => \N__31648\,
            lcout => \phase_controller_inst1.stoper_hc.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI1LP11_28_LC_8_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100111011"
        )
    port map (
            in0 => \N__25704\,
            in1 => \N__31707\,
            in2 => \N__25635\,
            in3 => \N__25664\,
            lcout => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIM9HS1_28_LC_8_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__24333\,
            in1 => \_gnd_net_\,
            in2 => \N__24312\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIM9HS1Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_8_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25202\,
            in2 => \N__24309\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_23_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32758\,
            in1 => \N__25155\,
            in2 => \_gnd_net_\,
            in3 => \N__24300\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__49137\,
            ce => 'H',
            sr => \N__48539\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__32762\,
            in1 => \N__24297\,
            in2 => \N__25425\,
            in3 => \N__24291\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__49137\,
            ce => 'H',
            sr => \N__48539\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32759\,
            in1 => \N__25389\,
            in2 => \_gnd_net_\,
            in3 => \N__24288\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__49137\,
            ce => 'H',
            sr => \N__48539\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32763\,
            in1 => \N__25368\,
            in2 => \_gnd_net_\,
            in3 => \N__24393\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__49137\,
            ce => 'H',
            sr => \N__48539\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32760\,
            in1 => \N__25320\,
            in2 => \_gnd_net_\,
            in3 => \N__24390\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__49137\,
            ce => 'H',
            sr => \N__48539\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32764\,
            in1 => \N__25284\,
            in2 => \_gnd_net_\,
            in3 => \N__24387\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__49137\,
            ce => 'H',
            sr => \N__48539\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32761\,
            in1 => \N__25263\,
            in2 => \_gnd_net_\,
            in3 => \N__24384\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__49137\,
            ce => 'H',
            sr => \N__48539\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32866\,
            in1 => \N__25233\,
            in2 => \_gnd_net_\,
            in3 => \N__24381\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_8_24_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__49132\,
            ce => 'H',
            sr => \N__48541\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32851\,
            in1 => \N__25605\,
            in2 => \_gnd_net_\,
            in3 => \N__24378\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__49132\,
            ce => 'H',
            sr => \N__48541\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32863\,
            in1 => \N__25572\,
            in2 => \_gnd_net_\,
            in3 => \N__24375\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__49132\,
            ce => 'H',
            sr => \N__48541\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32852\,
            in1 => \N__25542\,
            in2 => \_gnd_net_\,
            in3 => \N__24372\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__49132\,
            ce => 'H',
            sr => \N__48541\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32864\,
            in1 => \N__25515\,
            in2 => \_gnd_net_\,
            in3 => \N__24369\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__49132\,
            ce => 'H',
            sr => \N__48541\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32853\,
            in1 => \N__25485\,
            in2 => \_gnd_net_\,
            in3 => \N__24420\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__49132\,
            ce => 'H',
            sr => \N__48541\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32865\,
            in1 => \N__25452\,
            in2 => \_gnd_net_\,
            in3 => \N__24417\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__49132\,
            ce => 'H',
            sr => \N__48541\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32854\,
            in1 => \N__25791\,
            in2 => \_gnd_net_\,
            in3 => \N__24414\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__49132\,
            ce => 'H',
            sr => \N__48541\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32855\,
            in1 => \N__25824\,
            in2 => \_gnd_net_\,
            in3 => \N__24411\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_8_25_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__49125\,
            ce => 'H',
            sr => \N__48543\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32859\,
            in1 => \N__25896\,
            in2 => \_gnd_net_\,
            in3 => \N__24408\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__49125\,
            ce => 'H',
            sr => \N__48543\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32856\,
            in1 => \N__25880\,
            in2 => \_gnd_net_\,
            in3 => \N__24405\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \N__49125\,
            ce => 'H',
            sr => \N__48543\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_8_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32860\,
            in1 => \N__25842\,
            in2 => \_gnd_net_\,
            in3 => \N__24402\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \N__49125\,
            ce => 'H',
            sr => \N__48543\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_8_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32857\,
            in1 => \N__25854\,
            in2 => \_gnd_net_\,
            in3 => \N__24399\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\,
            clk => \N__49125\,
            ce => 'H',
            sr => \N__48543\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_8_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32861\,
            in1 => \N__25755\,
            in2 => \_gnd_net_\,
            in3 => \N__24396\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\,
            clk => \N__49125\,
            ce => 'H',
            sr => \N__48543\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_8_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32858\,
            in1 => \N__25767\,
            in2 => \_gnd_net_\,
            in3 => \N__24447\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\,
            clk => \N__49125\,
            ce => 'H',
            sr => \N__48543\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_8_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32862\,
            in1 => \N__25929\,
            in2 => \_gnd_net_\,
            in3 => \N__24444\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\,
            clk => \N__49125\,
            ce => 'H',
            sr => \N__48543\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_8_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32844\,
            in1 => \N__25941\,
            in2 => \_gnd_net_\,
            in3 => \N__24441\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_8_26_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\,
            clk => \N__49121\,
            ce => 'H',
            sr => \N__48545\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_8_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32848\,
            in1 => \N__25737\,
            in2 => \_gnd_net_\,
            in3 => \N__24438\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\,
            clk => \N__49121\,
            ce => 'H',
            sr => \N__48545\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_8_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32845\,
            in1 => \N__25725\,
            in2 => \_gnd_net_\,
            in3 => \N__24435\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\,
            clk => \N__49121\,
            ce => 'H',
            sr => \N__48545\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_8_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32849\,
            in1 => \N__26094\,
            in2 => \_gnd_net_\,
            in3 => \N__24432\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\,
            clk => \N__49121\,
            ce => 'H',
            sr => \N__48545\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_8_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32846\,
            in1 => \N__26106\,
            in2 => \_gnd_net_\,
            in3 => \N__24429\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\,
            clk => \N__49121\,
            ce => 'H',
            sr => \N__48545\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_8_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32850\,
            in1 => \N__25631\,
            in2 => \_gnd_net_\,
            in3 => \N__24426\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\,
            clk => \N__49121\,
            ce => 'H',
            sr => \N__48545\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_8_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32847\,
            in1 => \N__25663\,
            in2 => \_gnd_net_\,
            in3 => \N__24423\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49121\,
            ce => 'H',
            sr => \N__48545\
        );

    \phase_controller_inst2.S1_LC_8_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24567\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49112\,
            ce => 'H',
            sr => \N__48546\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26499\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D1_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24516\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_min_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49240\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_hc_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24495\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24474\,
            ce => 'H',
            sr => \N__48408\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011111110"
        )
    port map (
            in0 => \N__27370\,
            in1 => \N__27477\,
            in2 => \N__27177\,
            in3 => \N__24669\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49231\,
            ce => 'H',
            sr => \N__48417\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32573\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49231\,
            ce => 'H',
            sr => \N__48417\
        );

    \current_shift_inst.PI_CTRL.integrator_0_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__27473\,
            in1 => \N__27137\,
            in2 => \_gnd_net_\,
            in3 => \N__24579\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49231\,
            ce => 'H',
            sr => \N__48417\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__27133\,
            in1 => \N__27476\,
            in2 => \_gnd_net_\,
            in3 => \N__24714\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49231\,
            ce => 'H',
            sr => \N__48417\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__27474\,
            in1 => \N__27371\,
            in2 => \N__24732\,
            in3 => \N__27138\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49231\,
            ce => 'H',
            sr => \N__48417\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__27475\,
            in1 => \N__27372\,
            in2 => \N__24966\,
            in3 => \N__27139\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49231\,
            ce => 'H',
            sr => \N__48417\
        );

    \current_shift_inst.PI_CTRL.error_control_RNID56U_7_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__26013\,
            in1 => \N__32655\,
            in2 => \N__44598\,
            in3 => \N__29103\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNID56UZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26012\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__27126\,
            in1 => \N__27438\,
            in2 => \_gnd_net_\,
            in3 => \N__24687\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49226\,
            ce => 'H',
            sr => \N__48422\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__27434\,
            in1 => \N__27360\,
            in2 => \N__24840\,
            in3 => \N__27127\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49226\,
            ce => 'H',
            sr => \N__48422\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011111110"
        )
    port map (
            in0 => \N__27358\,
            in1 => \N__27436\,
            in2 => \N__27174\,
            in3 => \N__24825\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49226\,
            ce => 'H',
            sr => \N__48422\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__27435\,
            in1 => \N__27361\,
            in2 => \N__24813\,
            in3 => \N__27128\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49226\,
            ce => 'H',
            sr => \N__48422\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011111110"
        )
    port map (
            in0 => \N__27359\,
            in1 => \N__27437\,
            in2 => \N__27175\,
            in3 => \N__24798\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49226\,
            ce => 'H',
            sr => \N__48422\
        );

    \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26636\,
            in2 => \N__26640\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26244\,
            in2 => \N__26235\,
            in3 => \N__24570\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26220\,
            in2 => \N__32067\,
            in3 => \N__24717\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28902\,
            in2 => \N__26442\,
            in3 => \N__24705\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24702\,
            in2 => \N__24696\,
            in3 => \N__24681\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24678\,
            in2 => \N__26466\,
            in3 => \N__24660\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24657\,
            in2 => \N__24645\,
            in3 => \N__24624\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26781\,
            in2 => \N__26796\,
            in3 => \N__24621\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24618\,
            in2 => \N__24612\,
            in3 => \N__24597\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \bfn_9_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24594\,
            in2 => \N__26121\,
            in3 => \N__24582\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26073\,
            in2 => \N__26253\,
            in3 => \N__24846\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26112\,
            in2 => \N__26181\,
            in3 => \N__24843\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37848\,
            in2 => \N__26430\,
            in3 => \N__24828\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32124\,
            in2 => \N__26625\,
            in3 => \N__24816\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31860\,
            in2 => \N__26313\,
            in3 => \N__24801\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28950\,
            in2 => \N__26649\,
            in3 => \N__24789\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24786\,
            in2 => \N__26322\,
            in3 => \N__24768\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \bfn_9_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24765\,
            in2 => \N__24756\,
            in3 => \N__24735\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32283\,
            in2 => \N__26616\,
            in3 => \N__24987\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32220\,
            in2 => \N__26586\,
            in3 => \N__24978\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24975\,
            in2 => \N__26373\,
            in3 => \N__24954\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25959\,
            in2 => \N__26805\,
            in3 => \N__24939\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26859\,
            in2 => \N__26595\,
            in3 => \N__24927\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31800\,
            in2 => \N__26607\,
            in3 => \N__24918\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24915\,
            in2 => \N__29754\,
            in3 => \N__24891\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \bfn_9_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24888\,
            in2 => \N__26520\,
            in3 => \N__24870\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44694\,
            in2 => \N__29838\,
            in3 => \N__24858\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40017\,
            in2 => \N__26577\,
            in3 => \N__25032\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31923\,
            in2 => \N__29547\,
            in3 => \N__25017\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29884\,
            in2 => \N__29169\,
            in3 => \N__25014\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29886\,
            in2 => \N__40278\,
            in3 => \N__25011\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29885\,
            in2 => \N__26457\,
            in3 => \N__25008\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__27277\,
            in1 => \N__44565\,
            in2 => \_gnd_net_\,
            in3 => \N__25005\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRB3CP1_3_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24993\,
            in2 => \_gnd_net_\,
            in3 => \N__47691\,
            lcout => \elapsed_time_ns_1_RNIRB3CP1_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFKEE1_3_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__31105\,
            in1 => \N__28026\,
            in2 => \N__30255\,
            in3 => \N__30155\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_3_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__33293\,
            in1 => \N__30154\,
            in2 => \N__29676\,
            in3 => \N__32997\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49191\,
            ce => \N__32900\,
            sr => \N__48472\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8N721_6_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100010"
        )
    port map (
            in0 => \N__30001\,
            in1 => \N__31106\,
            in2 => \N__27864\,
            in3 => \N__47703\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUE3CP1_6_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__30251\,
            in1 => \_gnd_net_\,
            in2 => \N__25047\,
            in3 => \_gnd_net_\,
            lcout => \elapsed_time_ns_1_RNIUE3CP1_0_6\,
            ltout => \elapsed_time_ns_1_RNIUE3CP1_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__32996\,
            in1 => \N__33229\,
            in2 => \N__25044\,
            in3 => \N__33294\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49191\,
            ce => \N__32900\,
            sr => \N__48472\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__32995\,
            in1 => \N__27569\,
            in2 => \N__33309\,
            in3 => \N__33230\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49191\,
            ce => \N__32900\,
            sr => \N__48472\
        );

    \phase_controller_inst1.stoper_hc.target_time_15_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33202\,
            in1 => \N__30057\,
            in2 => \N__31400\,
            in3 => \N__27628\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49183\,
            ce => \N__32901\,
            sr => \N__48479\
        );

    \phase_controller_inst1.stoper_hc.target_time_1_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__27585\,
            in1 => \N__30195\,
            in2 => \N__27597\,
            in3 => \N__33314\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49183\,
            ce => \N__32901\,
            sr => \N__48479\
        );

    \phase_controller_inst1.stoper_hc.target_time_5_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__33203\,
            in1 => \N__28083\,
            in2 => \N__33315\,
            in3 => \N__33003\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49183\,
            ce => \N__32901\,
            sr => \N__48479\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI890221_16_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111000"
        )
    port map (
            in0 => \N__30762\,
            in1 => \N__31093\,
            in2 => \N__25106\,
            in3 => \N__47702\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIFFC6P1_16_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25041\,
            in3 => \N__30231\,
            lcout => \elapsed_time_ns_1_RNIFFC6P1_0_16\,
            ltout => \elapsed_time_ns_1_RNIFFC6P1_0_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_16_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010000"
        )
    port map (
            in0 => \N__33240\,
            in1 => \_gnd_net_\,
            in2 => \N__25074\,
            in3 => \N__31371\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49175\,
            ce => \N__34507\,
            sr => \N__48488\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111010101111"
        )
    port map (
            in0 => \N__25061\,
            in1 => \N__25070\,
            in2 => \N__34038\,
            in3 => \N__34064\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011001110"
        )
    port map (
            in0 => \N__25071\,
            in1 => \N__25062\,
            in2 => \N__34065\,
            in3 => \N__34037\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_17_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__31370\,
            in1 => \N__33242\,
            in2 => \_gnd_net_\,
            in3 => \N__29090\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49175\,
            ce => \N__34507\,
            sr => \N__48488\
        );

    \phase_controller_inst2.stoper_hc.target_time_19_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__33241\,
            in1 => \N__30945\,
            in2 => \_gnd_net_\,
            in3 => \N__31372\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49175\,
            ce => \N__34507\,
            sr => \N__48488\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__31272\,
            in1 => \N__34253\,
            in2 => \N__34224\,
            in3 => \N__31247\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILGKEE1_4_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__31043\,
            in1 => \N__30655\,
            in2 => \N__27565\,
            in3 => \N__27977\,
            lcout => \elapsed_time_ns_1_RNILGKEE1_0_4\,
            ltout => \elapsed_time_ns_1_RNILGKEE1_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3_2_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30938\,
            in1 => \N__28077\,
            in2 => \N__25053\,
            in3 => \N__31290\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4_2_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__29064\,
            in1 => \_gnd_net_\,
            in2 => \N__25050\,
            in3 => \N__25104\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_9_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__25105\,
            in1 => \N__29065\,
            in2 => \N__30949\,
            in3 => \N__31291\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9\,
            ltout => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_a2_10_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27734\,
            in2 => \N__25134\,
            in3 => \N__30051\,
            lcout => \phase_controller_inst1.stoper_hc.N_316\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4N_0_31_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__48588\,
            in1 => \N__27778\,
            in2 => \_gnd_net_\,
            in3 => \N__47633\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_342_i\,
            ltout => \delay_measurement_inst.delay_hc_timer.N_342_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHHC6P1_18_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25131\,
            in3 => \N__25125\,
            lcout => \elapsed_time_ns_1_RNIHHC6P1_0_18\,
            ltout => \elapsed_time_ns_1_RNIHHC6P1_0_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAB0221_18_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111000"
        )
    port map (
            in0 => \N__30743\,
            in1 => \N__31042\,
            in2 => \N__25128\,
            in3 => \N__47634\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGGC6P1_17_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25119\,
            in2 => \_gnd_net_\,
            in3 => \N__30238\,
            lcout => \elapsed_time_ns_1_RNIGGC6P1_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_16_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__31429\,
            in1 => \N__33121\,
            in2 => \_gnd_net_\,
            in3 => \N__25107\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49160\,
            ce => \N__32896\,
            sr => \N__48511\
        );

    \phase_controller_inst1.stoper_hc.N_267_i_1_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000010"
        )
    port map (
            in0 => \N__27754\,
            in1 => \N__27629\,
            in2 => \N__30330\,
            in3 => \N__30064\,
            lcout => \phase_controller_inst1.stoper_hc.N_267_iZ0Z_1\,
            ltout => \phase_controller_inst1.stoper_hc.N_267_iZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_9_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__26922\,
            in1 => \N__33120\,
            in2 => \N__25077\,
            in3 => \N__31425\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49155\,
            ce => \N__34575\,
            sr => \N__48518\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQBN721_9_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100100"
        )
    port map (
            in0 => \N__31124\,
            in1 => \N__26923\,
            in2 => \N__29741\,
            in3 => \N__47698\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1I3CP1_9_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25212\,
            in3 => \N__30252\,
            lcout => \elapsed_time_ns_1_RNI1I3CP1_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_15_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33119\,
            in1 => \N__30065\,
            in2 => \N__31441\,
            in3 => \N__27630\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49155\,
            ce => \N__34575\,
            sr => \N__48518\
        );

    \phase_controller_inst2.stoper_hc.target_time_14_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__33118\,
            in1 => \N__27758\,
            in2 => \N__31440\,
            in3 => \N__31479\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49155\,
            ce => \N__34575\,
            sr => \N__48518\
        );

    \phase_controller_inst1.stoper_hc.target_time_9_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__33239\,
            in1 => \N__25209\,
            in2 => \N__31442\,
            in3 => \N__26921\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49149\,
            ce => \N__32897\,
            sr => \N__48524\
        );

    \phase_controller_inst1.stoper_hc.target_time_12_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__31437\,
            in1 => \N__33237\,
            in2 => \N__30501\,
            in3 => \N__31494\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49142\,
            ce => \N__32898\,
            sr => \N__48529\
        );

    \phase_controller_inst1.stoper_hc.target_time_13_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__33235\,
            in1 => \N__31541\,
            in2 => \N__31504\,
            in3 => \N__31439\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49142\,
            ce => \N__32898\,
            sr => \N__48529\
        );

    \phase_controller_inst1.stoper_hc.target_time_14_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__31438\,
            in1 => \N__33238\,
            in2 => \N__27762\,
            in3 => \N__31495\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49142\,
            ce => \N__32898\,
            sr => \N__48529\
        );

    \phase_controller_inst1.stoper_hc.target_time_11_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__30539\,
            in1 => \N__33236\,
            in2 => \N__31443\,
            in3 => \N__31493\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49142\,
            ce => \N__32898\,
            sr => \N__48529\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25201\,
            in1 => \N__25176\,
            in2 => \N__25164\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_9_22_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32919\,
            in2 => \N__25143\,
            in3 => \N__25154\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25434\,
            in2 => \N__25410\,
            in3 => \N__25421\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25401\,
            in2 => \N__25377\,
            in3 => \N__25388\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25367\,
            in1 => \N__25356\,
            in2 => \N__25347\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25335\,
            in2 => \N__25308\,
            in3 => \N__25319\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25299\,
            in2 => \N__25272\,
            in3 => \N__25283\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25262\,
            in1 => \N__29010\,
            in2 => \N__25251\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25242\,
            in2 => \N__25221\,
            in3 => \N__25232\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_9_23_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29031\,
            in2 => \N__25593\,
            in3 => \N__25604\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25560\,
            in2 => \N__25584\,
            in3 => \N__25571\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25530\,
            in2 => \N__25554\,
            in3 => \N__25541\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25524\,
            in2 => \N__25503\,
            in3 => \N__25514\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25494\,
            in2 => \N__25473\,
            in3 => \N__25484\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25440\,
            in2 => \N__25464\,
            in3 => \N__25451\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_9_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25776\,
            in2 => \N__25911\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25947\,
            in2 => \N__25863\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_24_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25830\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25743\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25917\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25713\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26082\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25611\,
            in2 => \N__25668\,
            in3 => \N__25695\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_9_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25692\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25659\,
            in2 => \_gnd_net_\,
            in3 => \N__25630\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__25894\,
            in1 => \N__25876\,
            in2 => \N__29025\,
            in3 => \N__28599\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25940\,
            in2 => \_gnd_net_\,
            in3 => \N__25928\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_df24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_9_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001100010000"
        )
    port map (
            in0 => \N__25790\,
            in1 => \N__25823\,
            in2 => \N__25809\,
            in3 => \N__29045\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_9_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__28598\,
            in1 => \N__25895\,
            in2 => \N__25881\,
            in3 => \N__29024\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_9_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25853\,
            in2 => \_gnd_net_\,
            in3 => \N__25841\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_df20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_9_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010011110101"
        )
    port map (
            in0 => \N__25822\,
            in1 => \N__25808\,
            in2 => \N__29046\,
            in3 => \N__25789\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_9_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25766\,
            in2 => \_gnd_net_\,
            in3 => \N__25754\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_df22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_9_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25736\,
            in2 => \_gnd_net_\,
            in3 => \N__25724\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_df26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_9_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26105\,
            in2 => \_gnd_net_\,
            in3 => \N__26093\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_df28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26299\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29389\,
            in2 => \_gnd_net_\,
            in3 => \N__44586\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI78BM_30_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26683\,
            in1 => \N__31969\,
            in2 => \N__32167\,
            in3 => \N__27356\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIC35V7_13_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26061\,
            in1 => \N__26052\,
            in2 => \N__26043\,
            in3 => \N__25989\,
            lcout => \current_shift_inst.PI_CTRL.N_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__26167\,
            in1 => \N__26040\,
            in2 => \N__26759\,
            in3 => \N__26300\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110011"
        )
    port map (
            in0 => \N__26187\,
            in1 => \N__26492\,
            in2 => \N__26031\,
            in3 => \N__26020\,
            lcout => \current_shift_inst.PI_CTRL.N_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__48583\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pll_inst.red_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26845\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32383\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26200\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_0\,
            ltout => \current_shift_inst.PI_CTRL.integrator_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI1M2U_4_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__32384\,
            in1 => \N__44535\,
            in2 => \N__26238\,
            in3 => \N__29124\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI1M2UZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__27170\,
            in1 => \N__27439\,
            in2 => \_gnd_net_\,
            in3 => \N__26226\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49215\,
            ce => 'H',
            sr => \N__48412\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32091\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__32092\,
            in1 => \N__28929\,
            in2 => \_gnd_net_\,
            in3 => \N__26201\,
            lcout => \current_shift_inst.PI_CTRL.un1_enablelt3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVH_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110101111"
        )
    port map (
            in0 => \N__32508\,
            in1 => \N__27009\,
            in2 => \N__44597\,
            in3 => \N__29244\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIM1S01_12_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110011"
        )
    port map (
            in0 => \N__26168\,
            in1 => \N__32574\,
            in2 => \N__29280\,
            in3 => \N__44570\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIM1S01Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27008\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIHA7U_8_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__26511\,
            in1 => \N__44569\,
            in2 => \N__33390\,
            in3 => \N__29331\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIHA7UZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44199\,
            lcout => \current_shift_inst.un4_control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26682\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI905U_6_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__28937\,
            in1 => \N__32681\,
            in2 => \N__44596\,
            in3 => \N__29112\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI905UZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11I_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011111111"
        )
    port map (
            in0 => \N__32486\,
            in1 => \N__37877\,
            in2 => \N__29235\,
            in3 => \N__44574\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82J_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011111111"
        )
    port map (
            in0 => \N__29364\,
            in1 => \N__26415\,
            in2 => \N__29343\,
            in3 => \N__44531\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5I_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110101111"
        )
    port map (
            in0 => \N__31995\,
            in1 => \N__26361\,
            in2 => \N__44584\,
            in3 => \N__29469\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73I_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011111111"
        )
    port map (
            in0 => \N__29520\,
            in1 => \N__31899\,
            in2 => \N__29496\,
            in3 => \N__44522\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIQ6T01_13_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__26298\,
            in1 => \N__32541\,
            in2 => \N__44583\,
            in3 => \N__29253\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIQ6T01Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4I_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011111111"
        )
    port map (
            in0 => \N__37926\,
            in1 => \N__28997\,
            in2 => \N__29481\,
            in3 => \N__44524\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_0_14_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44518\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_i_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42I_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011111111"
        )
    port map (
            in0 => \N__29868\,
            in1 => \N__32168\,
            in2 => \N__29532\,
            in3 => \N__44523\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20J_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__32326\,
            in1 => \N__29433\,
            in2 => \N__44585\,
            in3 => \N__29406\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96J_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__31847\,
            in1 => \N__29610\,
            in2 => \N__44592\,
            in3 => \N__29583\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65J_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111110011"
        )
    port map (
            in0 => \N__26897\,
            in1 => \N__44555\,
            in2 => \N__32208\,
            in3 => \N__29619\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51J_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110101111"
        )
    port map (
            in0 => \N__29397\,
            in1 => \N__32270\,
            in2 => \N__44591\,
            in3 => \N__29373\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJ_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110111011"
        )
    port map (
            in0 => \N__44928\,
            in1 => \N__44559\,
            in2 => \N__40074\,
            in3 => \N__29559\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8J_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110101111"
        )
    port map (
            in0 => \N__40446\,
            in1 => \N__26568\,
            in2 => \N__44593\,
            in3 => \N__29571\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41697\,
            lcout => \current_shift_inst.un4_control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26896\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34J_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011111111"
        )
    port map (
            in0 => \N__26846\,
            in1 => \N__29664\,
            in2 => \N__29637\,
            in3 => \N__44554\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI7T941_10_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__26728\,
            in1 => \N__44587\,
            in2 => \N__29307\,
            in3 => \N__33443\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI7T941Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26727\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000111110101"
        )
    port map (
            in0 => \N__27345\,
            in1 => \N__27500\,
            in2 => \N__27197\,
            in3 => \N__26769\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49193\,
            ce => 'H',
            sr => \N__48441\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__27497\,
            in1 => \N__27347\,
            in2 => \N__26712\,
            in3 => \N__27188\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49193\,
            ce => 'H',
            sr => \N__48441\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011111110"
        )
    port map (
            in0 => \N__27343\,
            in1 => \N__27498\,
            in2 => \N__27195\,
            in3 => \N__26703\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49193\,
            ce => 'H',
            sr => \N__48441\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011111110"
        )
    port map (
            in0 => \N__27344\,
            in1 => \N__27499\,
            in2 => \N__27196\,
            in3 => \N__26697\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49193\,
            ce => 'H',
            sr => \N__48441\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__27496\,
            in1 => \N__27346\,
            in2 => \N__27213\,
            in3 => \N__27187\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49193\,
            ce => 'H',
            sr => \N__48441\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI63452_2_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000000"
        )
    port map (
            in0 => \N__28025\,
            in1 => \N__26939\,
            in2 => \N__27978\,
            in3 => \N__27687\,
            lcout => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_2_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__27743\,
            in1 => \N__26930\,
            in2 => \N__30066\,
            in3 => \N__26976\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2\,
            ltout => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_0_a5_1_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__26958\,
            in1 => \N__30082\,
            in2 => \N__26964\,
            in3 => \N__31376\,
            lcout => \phase_controller_inst1.stoper_hc.N_308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJEKEE1_2_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__26948\,
            in1 => \N__26940\,
            in2 => \N__30690\,
            in3 => \N__31112\,
            lcout => \elapsed_time_ns_1_RNIJEKEE1_0_2\,
            ltout => \elapsed_time_ns_1_RNIJEKEE1_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_0_o2_1_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26961\,
            in3 => \N__30149\,
            lcout => \phase_controller_inst1.stoper_hc.N_284\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_0_2_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100001111"
        )
    port map (
            in0 => \N__30150\,
            in1 => \N__30083\,
            in2 => \N__26952\,
            in3 => \N__29687\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28005\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49185\,
            ce => \N__28623\,
            sr => \N__48453\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0_6_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110111011"
        )
    port map (
            in0 => \N__30323\,
            in1 => \N__27744\,
            in2 => \_gnd_net_\,
            in3 => \N__26931\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0_6_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011100"
        )
    port map (
            in0 => \N__30062\,
            in1 => \N__27627\,
            in2 => \N__27603\,
            in3 => \N__31346\,
            lcout => \phase_controller_inst1.stoper_hc.N_326\,
            ltout => \phase_controller_inst1.stoper_hc.N_326_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_1_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30189\,
            in2 => \N__27600\,
            in3 => \N__33183\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1\,
            ltout => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_1_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__30190\,
            in1 => \N__33306\,
            in2 => \N__27588\,
            in3 => \N__27581\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49177\,
            ce => \N__34502\,
            sr => \N__48460\
        );

    \phase_controller_inst2.stoper_hc.target_time_4_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__33184\,
            in1 => \N__33307\,
            in2 => \N__33034\,
            in3 => \N__27570\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49177\,
            ce => \N__34502\,
            sr => \N__48460\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29924\,
            in1 => \N__28760\,
            in2 => \N__28812\,
            in3 => \N__30296\,
            lcout => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAMU8E1_27_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__31099\,
            in1 => \N__27540\,
            in2 => \N__30685\,
            in3 => \N__28811\,
            lcout => \elapsed_time_ns_1_RNIAMU8E1_0_27\,
            ltout => \elapsed_time_ns_1_RNIAMU8E1_0_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6_15_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30362\,
            in1 => \N__27794\,
            in2 => \N__27534\,
            in3 => \N__27674\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJKEE1_7_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__30677\,
            in1 => \N__30114\,
            in2 => \N__31122\,
            in3 => \N__29721\,
            lcout => \elapsed_time_ns_1_RNIOJKEE1_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI6IU8E1_23_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__31103\,
            in1 => \N__27531\,
            in2 => \N__30686\,
            in3 => \N__30870\,
            lcout => \elapsed_time_ns_1_RNI6IU8E1_0_23\,
            ltout => \elapsed_time_ns_1_RNI6IU8E1_0_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0_15_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27699\,
            in3 => \N__27806\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_o5_15_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27641\,
            in1 => \N__30453\,
            in2 => \N__27696\,
            in3 => \N__27693\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__27860\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27917\,
            lcout => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9LU8E1_26_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__30852\,
            in1 => \N__30663\,
            in2 => \N__27678\,
            in3 => \N__31066\,
            lcout => \elapsed_time_ns_1_RNI9LU8E1_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDDC6P1_14_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__27705\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30253\,
            lcout => \elapsed_time_ns_1_RNIDDC6P1_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPR8P8_10_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29700\,
            in1 => \N__30696\,
            in2 => \N__27663\,
            in3 => \N__27651\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlt31_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP0VUB_31_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111011"
        )
    port map (
            in0 => \N__28637\,
            in1 => \N__49968\,
            in2 => \N__27645\,
            in3 => \N__42450\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_367\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5HU8E1_22_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__27642\,
            in1 => \N__30665\,
            in2 => \N__31749\,
            in3 => \N__31068\,
            lcout => \elapsed_time_ns_1_RNI5HU8E1_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7IT8E1_15_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__30666\,
            in1 => \N__30058\,
            in2 => \N__31108\,
            in3 => \N__30720\,
            lcout => \elapsed_time_ns_1_RNI7IT8E1_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7JU8E1_24_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__27807\,
            in1 => \N__30664\,
            in2 => \N__30888\,
            in3 => \N__31067\,
            lcout => \elapsed_time_ns_1_RNI7JU8E1_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBNU8E1_28_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__30662\,
            in1 => \N__28761\,
            in2 => \N__31107\,
            in3 => \N__27795\,
            lcout => \elapsed_time_ns_1_RNIBNU8E1_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMHKEE1_5_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__28082\,
            in1 => \N__30667\,
            in2 => \N__27918\,
            in3 => \N__31072\,
            lcout => \elapsed_time_ns_1_RNIMHKEE1_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5GT8E1_13_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__30668\,
            in1 => \N__31537\,
            in2 => \N__31109\,
            in3 => \N__31203\,
            lcout => \elapsed_time_ns_1_RNI5GT8E1_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIIC6P1_19_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__30915\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30232\,
            lcout => \elapsed_time_ns_1_RNIIIC6P1_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0TDSM_31_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47630\,
            in2 => \_gnd_net_\,
            in3 => \N__27779\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_365_clk\,
            ltout => \delay_measurement_inst.delay_hc_timer.N_365_clk_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4FT8E1_12_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__30494\,
            in1 => \N__31173\,
            in2 => \N__27783\,
            in3 => \N__30669\,
            lcout => \elapsed_time_ns_1_RNI4FT8E1_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4N_31_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__48587\,
            in1 => \N__47631\,
            in2 => \_gnd_net_\,
            in3 => \N__27780\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31\,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4GU8E1_21_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__30468\,
            in1 => \N__30825\,
            in2 => \N__27765\,
            in3 => \N__31073\,
            lcout => \elapsed_time_ns_1_RNI4GU8E1_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI670221_14_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001110"
        )
    port map (
            in0 => \N__27742\,
            in1 => \N__47632\,
            in2 => \N__31110\,
            in3 => \N__31188\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_5_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__28078\,
            in1 => \N__33310\,
            in2 => \N__33042\,
            in3 => \N__33117\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49150\,
            ce => \N__34506\,
            sr => \N__48492\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5IV8E1_31_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__28638\,
            in1 => \N__30673\,
            in2 => \N__33180\,
            in3 => \N__31092\,
            lcout => \elapsed_time_ns_1_RNI5IV8E1_0_31\,
            ltout => \elapsed_time_ns_1_RNI5IV8E1_0_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_7_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__33040\,
            in1 => \_gnd_net_\,
            in2 => \N__28056\,
            in3 => \N__30118\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49150\,
            ce => \N__34506\,
            sr => \N__48492\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28049\,
            in2 => \N__27948\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_10_19_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__49144\,
            ce => \N__28622\,
            sr => \N__48504\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28001\,
            in2 => \N__27893\,
            in3 => \N__27951\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__49144\,
            ce => \N__28622\,
            sr => \N__48504\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27947\,
            in2 => \N__27839\,
            in3 => \N__27897\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__49144\,
            ce => \N__28622\,
            sr => \N__48504\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28343\,
            in2 => \N__27894\,
            in3 => \N__27843\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__49144\,
            ce => \N__28622\,
            sr => \N__48504\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28316\,
            in2 => \N__27840\,
            in3 => \N__27810\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__49144\,
            ce => \N__28622\,
            sr => \N__48504\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28292\,
            in2 => \N__28347\,
            in3 => \N__28320\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__49144\,
            ce => \N__28622\,
            sr => \N__48504\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28317\,
            in2 => \N__28268\,
            in3 => \N__28296\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__49144\,
            ce => \N__28622\,
            sr => \N__48504\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28293\,
            in2 => \N__28232\,
            in3 => \N__28272\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__49144\,
            ce => \N__28622\,
            sr => \N__48504\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28196\,
            in2 => \N__28269\,
            in3 => \N__28239\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_10_20_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__49139\,
            ce => \N__28621\,
            sr => \N__48512\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28163\,
            in2 => \N__28236\,
            in3 => \N__28203\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__49139\,
            ce => \N__28621\,
            sr => \N__48512\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28136\,
            in2 => \N__28200\,
            in3 => \N__28167\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__49139\,
            ce => \N__28621\,
            sr => \N__48512\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28164\,
            in2 => \N__28112\,
            in3 => \N__28140\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__49139\,
            ce => \N__28621\,
            sr => \N__48512\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28137\,
            in2 => \N__28586\,
            in3 => \N__28116\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__49139\,
            ce => \N__28621\,
            sr => \N__48512\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28550\,
            in2 => \N__28113\,
            in3 => \N__28086\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__49139\,
            ce => \N__28621\,
            sr => \N__48512\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28514\,
            in2 => \N__28587\,
            in3 => \N__28557\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__49139\,
            ce => \N__28621\,
            sr => \N__48512\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28487\,
            in2 => \N__28554\,
            in3 => \N__28521\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__49139\,
            ce => \N__28621\,
            sr => \N__48512\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28460\,
            in2 => \N__28518\,
            in3 => \N__28491\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_10_21_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__49134\,
            ce => \N__28619\,
            sr => \N__48519\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28488\,
            in2 => \N__28436\,
            in3 => \N__28464\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__49134\,
            ce => \N__28619\,
            sr => \N__48519\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28461\,
            in2 => \N__28406\,
            in3 => \N__28440\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__49134\,
            ce => \N__28619\,
            sr => \N__48519\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28373\,
            in2 => \N__28437\,
            in3 => \N__28410\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__49134\,
            ce => \N__28619\,
            sr => \N__48519\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28889\,
            in2 => \N__28407\,
            in3 => \N__28380\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__49134\,
            ce => \N__28619\,
            sr => \N__48519\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28865\,
            in2 => \N__28377\,
            in3 => \N__28350\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__49134\,
            ce => \N__28619\,
            sr => \N__48519\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28890\,
            in2 => \N__28841\,
            in3 => \N__28869\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__49134\,
            ce => \N__28619\,
            sr => \N__48519\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28866\,
            in2 => \N__28793\,
            in3 => \N__28845\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__49134\,
            ce => \N__28619\,
            sr => \N__48519\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28736\,
            in2 => \N__28842\,
            in3 => \N__28797\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_10_22_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__49127\,
            ce => \N__28618\,
            sr => \N__48525\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28670\,
            in2 => \N__28794\,
            in3 => \N__28740\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__49127\,
            ce => \N__28618\,
            sr => \N__48525\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28737\,
            in2 => \N__28716\,
            in3 => \N__28695\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__49127\,
            ce => \N__28618\,
            sr => \N__48525\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28692\,
            in2 => \N__28674\,
            in3 => \N__28644\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__49127\,
            ce => \N__28618\,
            sr => \N__48525\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28641\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49127\,
            ce => \N__28618\,
            sr => \N__48525\
        );

    \phase_controller_inst1.stoper_hc.target_time_18_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__33187\,
            in1 => \N__31431\,
            in2 => \_gnd_net_\,
            in3 => \N__31305\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49122\,
            ce => \N__32879\,
            sr => \N__48530\
        );

    \phase_controller_inst1.stoper_hc.target_time_17_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__33186\,
            in1 => \N__29083\,
            in2 => \_gnd_net_\,
            in3 => \N__31432\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49122\,
            ce => \N__32879\,
            sr => \N__48530\
        );

    \phase_controller_inst1.stoper_hc.target_time_10_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__33188\,
            in1 => \N__31489\,
            in2 => \N__30570\,
            in3 => \N__31433\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49122\,
            ce => \N__32879\,
            sr => \N__48530\
        );

    \phase_controller_inst1.stoper_hc.target_time_19_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__31430\,
            in1 => \N__33189\,
            in2 => \_gnd_net_\,
            in3 => \N__30950\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49122\,
            ce => \N__32879\,
            sr => \N__48530\
        );

    \phase_controller_inst1.stoper_hc.target_time_8_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__31236\,
            in1 => \N__33190\,
            in2 => \_gnd_net_\,
            in3 => \N__33018\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49122\,
            ce => \N__32879\,
            sr => \N__48530\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__29515\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44581\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__29428\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44582\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44514\,
            in2 => \_gnd_net_\,
            in3 => \N__29362\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28998\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28933\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29214\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29154\,
            in2 => \_gnd_net_\,
            in3 => \N__36836\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29148\,
            in2 => \_gnd_net_\,
            in3 => \N__32453\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29142\,
            in2 => \_gnd_net_\,
            in3 => \N__32429\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29136\,
            in2 => \_gnd_net_\,
            in3 => \N__32408\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29130\,
            in2 => \_gnd_net_\,
            in3 => \N__29118\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32040\,
            in2 => \_gnd_net_\,
            in3 => \N__29115\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32514\,
            in2 => \_gnd_net_\,
            in3 => \N__29106\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31788\,
            in2 => \_gnd_net_\,
            in3 => \N__29094\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33402\,
            in3 => \N__29325\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_8\,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33327\,
            in2 => \_gnd_net_\,
            in3 => \N__29310\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33420\,
            in2 => \_gnd_net_\,
            in3 => \N__29295\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32046\,
            in2 => \_gnd_net_\,
            in3 => \N__29283\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNI9BCC_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32052\,
            in2 => \_gnd_net_\,
            in3 => \N__29268\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNIBEDC_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29265\,
            in2 => \_gnd_net_\,
            in3 => \N__29247\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32503\,
            in2 => \_gnd_net_\,
            in3 => \N__29238\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32479\,
            in2 => \_gnd_net_\,
            in3 => \N__29226\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29867\,
            in2 => \_gnd_net_\,
            in3 => \N__29523\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29516\,
            in2 => \_gnd_net_\,
            in3 => \N__29484\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37922\,
            in2 => \_gnd_net_\,
            in3 => \N__29472\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31994\,
            in2 => \_gnd_net_\,
            in3 => \N__29463\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29460\,
            in2 => \_gnd_net_\,
            in3 => \N__29436\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29429\,
            in2 => \_gnd_net_\,
            in3 => \N__29400\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29396\,
            in2 => \_gnd_net_\,
            in3 => \N__29367\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29363\,
            in2 => \_gnd_net_\,
            in3 => \N__29334\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29663\,
            in2 => \_gnd_net_\,
            in3 => \N__29622\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32204\,
            in3 => \N__29613\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29609\,
            in2 => \_gnd_net_\,
            in3 => \N__29577\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29825\,
            in2 => \_gnd_net_\,
            in3 => \N__29574\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40445\,
            in2 => \_gnd_net_\,
            in3 => \N__29565\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44282\,
            in2 => \_gnd_net_\,
            in3 => \N__29562\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44924\,
            in2 => \_gnd_net_\,
            in3 => \N__29553\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74K_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \N__31971\,
            in1 => \N__44400\,
            in2 => \_gnd_net_\,
            in3 => \N__29550\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74KZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D2_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29901\,
            lcout => \il_min_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49186\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_14_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44380\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_i_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__29866\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44374\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9J_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__44740\,
            in1 => \N__44283\,
            in2 => \N__44474\,
            in3 => \N__29844\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44375\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29826\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\,
            ltout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7J_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111110011"
        )
    port map (
            in0 => \N__29804\,
            in1 => \N__44376\,
            in2 => \N__29763\,
            in3 => \N__29760\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_2_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000110010"
        )
    port map (
            in0 => \N__33291\,
            in1 => \N__33185\,
            in2 => \N__33019\,
            in3 => \N__32930\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49178\,
            ce => \N__34574\,
            sr => \N__48442\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_10_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29742\,
            in1 => \N__29720\,
            in2 => \N__30810\,
            in3 => \N__30350\,
            lcout => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_3_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__31345\,
            in1 => \N__33181\,
            in2 => \N__30087\,
            in3 => \N__29688\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3\,
            ltout => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_3_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__30162\,
            in1 => \N__32999\,
            in2 => \N__30129\,
            in3 => \N__33308\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49169\,
            ce => \N__34558\,
            sr => \N__48454\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0_2_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__31231\,
            in1 => \N__30122\,
            in2 => \N__30006\,
            in3 => \N__30322\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2\,
            ltout => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_6_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__30063\,
            in1 => \_gnd_net_\,
            in2 => \N__30009\,
            in3 => \N__31344\,
            lcout => \phase_controller_inst1.stoper_hc.N_328\,
            ltout => \phase_controller_inst1.stoper_hc.N_328_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_6_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__30005\,
            in1 => \N__32998\,
            in2 => \N__29985\,
            in3 => \N__33182\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49169\,
            ce => \N__34558\,
            sr => \N__48454\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30389\,
            in2 => \_gnd_net_\,
            in3 => \N__30407\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__34441\,
            in1 => \N__30408\,
            in2 => \N__33792\,
            in3 => \N__30390\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49161\,
            ce => 'H',
            sr => \N__48461\
        );

    \phase_controller_inst2.stoper_hc.running_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111110000"
        )
    port map (
            in0 => \N__30443\,
            in1 => \N__33800\,
            in2 => \N__29981\,
            in3 => \N__30391\,
            lcout => \phase_controller_inst2.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49161\,
            ce => 'H',
            sr => \N__48461\
        );

    \phase_controller_inst2.stoper_hc.time_passed_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011000010101010"
        )
    port map (
            in0 => \N__29950\,
            in1 => \N__33801\,
            in2 => \N__30447\,
            in3 => \N__30392\,
            lcout => \phase_controller_inst2.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49161\,
            ce => 'H',
            sr => \N__48461\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICOU8E1_29_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__29928\,
            in1 => \N__30657\,
            in2 => \N__31104\,
            in3 => \N__29907\,
            lcout => \elapsed_time_ns_1_RNICOU8E1_0_29\,
            ltout => \elapsed_time_ns_1_RNICOU8E1_0_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7_15_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30278\,
            in1 => \N__30467\,
            in2 => \N__30456\,
            in3 => \N__30581\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI5B3T_28_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110101"
        )
    port map (
            in0 => \N__30442\,
            in1 => \N__35142\,
            in2 => \N__33819\,
            in3 => \N__35171\,
            lcout => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNITOIN1_28_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30399\,
            in3 => \N__30396\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNITOIN1Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8KU8E1_25_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__31056\,
            in1 => \N__30906\,
            in2 => \N__30366\,
            in3 => \N__30661\,
            lcout => \elapsed_time_ns_1_RNI8KU8E1_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2DT8E1_10_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__30656\,
            in1 => \N__31055\,
            in2 => \N__30562\,
            in3 => \N__30351\,
            lcout => \elapsed_time_ns_1_RNI2DT8E1_0_10\,
            ltout => \elapsed_time_ns_1_RNI2DT8E1_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2_2_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30489\,
            in1 => \N__31524\,
            in2 => \N__30333\,
            in3 => \N__30522\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4HV8E1_30_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__30279\,
            in1 => \N__30300\,
            in2 => \N__30684\,
            in3 => \N__31057\,
            lcout => \elapsed_time_ns_1_RNI4HV8E1_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII3N721_1_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111010"
        )
    port map (
            in0 => \N__47677\,
            in1 => \N__30270\,
            in2 => \N__30194\,
            in3 => \N__31085\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP93CP1_1_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30258\,
            in3 => \N__30254\,
            lcout => \elapsed_time_ns_1_RNIP93CP1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3ET8E1_11_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__31155\,
            in1 => \N__30671\,
            in2 => \N__30538\,
            in3 => \N__31081\,
            lcout => \elapsed_time_ns_1_RNI3ET8E1_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPKKEE1_8_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__30672\,
            in1 => \N__31235\,
            in2 => \N__31111\,
            in3 => \N__30806\,
            lcout => \elapsed_time_ns_1_RNIPKKEE1_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30785\,
            in1 => \N__30758\,
            in2 => \N__30744\,
            in3 => \N__30716\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPFU14_11_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__31731\,
            in1 => \N__30834\,
            in2 => \N__30699\,
            in3 => \N__31140\,
            lcout => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3FU8E1_20_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__30582\,
            in1 => \N__30670\,
            in2 => \N__31782\,
            in3 => \N__31080\,
            lcout => \elapsed_time_ns_1_RNI3FU8E1_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_10_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__33225\,
            in1 => \N__30566\,
            in2 => \N__31505\,
            in3 => \N__31398\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49145\,
            ce => \N__34559\,
            sr => \N__48480\
        );

    \phase_controller_inst2.stoper_hc.target_time_11_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__31395\,
            in1 => \N__31502\,
            in2 => \N__30540\,
            in3 => \N__33228\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49145\,
            ce => \N__34559\,
            sr => \N__48480\
        );

    \phase_controller_inst2.stoper_hc.target_time_12_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__33226\,
            in1 => \N__30493\,
            in2 => \N__31506\,
            in3 => \N__31399\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49145\,
            ce => \N__34559\,
            sr => \N__48480\
        );

    \phase_controller_inst2.stoper_hc.target_time_13_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__31396\,
            in1 => \N__33227\,
            in2 => \N__31542\,
            in3 => \N__31503\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49145\,
            ce => \N__34559\,
            sr => \N__48480\
        );

    \phase_controller_inst2.stoper_hc.target_time_18_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__33223\,
            in1 => \N__31397\,
            in2 => \_gnd_net_\,
            in3 => \N__31304\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49145\,
            ce => \N__34559\,
            sr => \N__48480\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000100"
        )
    port map (
            in0 => \N__34216\,
            in1 => \N__31268\,
            in2 => \N__34254\,
            in3 => \N__31254\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_8_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__33224\,
            in1 => \N__33036\,
            in2 => \_gnd_net_\,
            in3 => \N__31230\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49145\,
            ce => \N__34559\,
            sr => \N__48480\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMHD01_11_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31199\,
            in1 => \N__31184\,
            in2 => \N__31172\,
            in3 => \N__31151\,
            lcout => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0_9_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__46885\,
            in1 => \N__42129\,
            in2 => \_gnd_net_\,
            in3 => \N__46320\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC0221_19_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111000"
        )
    port map (
            in0 => \N__31760\,
            in1 => \N__31123\,
            in2 => \N__30954\,
            in3 => \N__47700\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30899\,
            in1 => \N__30881\,
            in2 => \N__30869\,
            in3 => \N__30845\,
            lcout => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30821\,
            in1 => \N__31772\,
            in2 => \N__31761\,
            in3 => \N__31742\,
            lcout => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_tr_RNO_0_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__35557\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34357\,
            lcout => \phase_controller_inst1.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_1_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35615\,
            in2 => \_gnd_net_\,
            in3 => \N__31613\,
            lcout => \phase_controller_inst1.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_0_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34309\,
            in2 => \_gnd_net_\,
            in3 => \N__31567\,
            lcout => \phase_controller_inst1.start_timer_hc_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.start_latched_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31644\,
            lcout => \phase_controller_inst1.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49123\,
            ce => 'H',
            sr => \N__48520\
        );

    \phase_controller_inst1.state_3_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__35628\,
            in1 => \N__35424\,
            in2 => \N__31620\,
            in3 => \N__31682\,
            lcout => state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49123\,
            ce => 'H',
            sr => \N__48520\
        );

    \phase_controller_inst1.start_timer_hc_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__35408\,
            in1 => \N__31662\,
            in2 => \N__31650\,
            in3 => \N__31656\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49123\,
            ce => 'H',
            sr => \N__48520\
        );

    \phase_controller_inst1.state_2_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001100"
        )
    port map (
            in0 => \N__31612\,
            in1 => \N__34302\,
            in2 => \N__31578\,
            in3 => \N__35629\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49118\,
            ce => 'H',
            sr => \N__48526\
        );

    \phase_controller_inst1.state_1_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__31577\,
            in1 => \N__34308\,
            in2 => \N__35568\,
            in3 => \N__34361\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49115\,
            ce => 'H',
            sr => \N__48531\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_11_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32034\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40922\,
            in2 => \_gnd_net_\,
            in3 => \N__37507\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_395_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_tr_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37545\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32004\,
            ce => 'H',
            sr => \N__48396\
        );

    \delay_measurement_inst.stop_timer_tr_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37546\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32004\,
            ce => 'H',
            sr => \N__48396\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44513\,
            in2 => \_gnd_net_\,
            in3 => \N__31987\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31968\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31900\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31843\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32650\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32327\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32265\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43579\,
            lcout => \current_shift_inst.un4_control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__32197\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44495\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32163\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI5R3U_5_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44512\,
            in1 => \N__32108\,
            in2 => \N__32351\,
            in3 => \N__32073\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI5R3UZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32566\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32599\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32344\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32669\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__32507\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44510\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44511\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32487\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34686\,
            in1 => \N__32466\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axb_0\,
            ltout => OPEN,
            carryin => \bfn_12_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_1_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34680\,
            in2 => \_gnd_net_\,
            in3 => \N__32439\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            clk => \N__49192\,
            ce => 'H',
            sr => \N__48413\
        );

    \current_shift_inst.PI_CTRL.error_control_2_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34671\,
            in2 => \_gnd_net_\,
            in3 => \N__32415\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            clk => \N__49192\,
            ce => 'H',
            sr => \N__48413\
        );

    \current_shift_inst.PI_CTRL.error_control_3_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34767\,
            in2 => \_gnd_net_\,
            in3 => \N__32391\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            clk => \N__49192\,
            ce => 'H',
            sr => \N__48413\
        );

    \current_shift_inst.PI_CTRL.error_control_4_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34758\,
            in2 => \_gnd_net_\,
            in3 => \N__32361\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            clk => \N__49192\,
            ce => 'H',
            sr => \N__48413\
        );

    \current_shift_inst.PI_CTRL.error_control_5_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34749\,
            in2 => \_gnd_net_\,
            in3 => \N__32331\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            clk => \N__49192\,
            ce => 'H',
            sr => \N__48413\
        );

    \current_shift_inst.PI_CTRL.error_control_6_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34740\,
            in2 => \_gnd_net_\,
            in3 => \N__32658\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            clk => \N__49192\,
            ce => 'H',
            sr => \N__48413\
        );

    \current_shift_inst.PI_CTRL.error_control_7_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34731\,
            in2 => \_gnd_net_\,
            in3 => \N__32625\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            clk => \N__49192\,
            ce => 'H',
            sr => \N__48413\
        );

    \current_shift_inst.PI_CTRL.error_control_8_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34722\,
            in2 => \_gnd_net_\,
            in3 => \N__32622\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_8\,
            ltout => OPEN,
            carryin => \bfn_12_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            clk => \N__49184\,
            ce => 'H',
            sr => \N__48418\
        );

    \current_shift_inst.PI_CTRL.error_control_9_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34713\,
            in2 => \_gnd_net_\,
            in3 => \N__32619\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            clk => \N__49184\,
            ce => 'H',
            sr => \N__48418\
        );

    \current_shift_inst.PI_CTRL.error_control_10_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34704\,
            in2 => \_gnd_net_\,
            in3 => \N__32616\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            clk => \N__49184\,
            ce => 'H',
            sr => \N__48418\
        );

    \current_shift_inst.PI_CTRL.error_control_11_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34812\,
            in2 => \_gnd_net_\,
            in3 => \N__32577\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            clk => \N__49184\,
            ce => 'H',
            sr => \N__48418\
        );

    \current_shift_inst.PI_CTRL.error_control_12_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34803\,
            in2 => \_gnd_net_\,
            in3 => \N__32544\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            clk => \N__49184\,
            ce => 'H',
            sr => \N__48418\
        );

    \current_shift_inst.PI_CTRL.error_control_13_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33408\,
            in2 => \_gnd_net_\,
            in3 => \N__32520\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            clk => \N__49184\,
            ce => 'H',
            sr => \N__48418\
        );

    \current_shift_inst.PI_CTRL.error_control_14_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34791\,
            in2 => \_gnd_net_\,
            in3 => \N__32517\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49184\,
            ce => 'H',
            sr => \N__48418\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33431\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37290\,
            in2 => \_gnd_net_\,
            in3 => \N__37314\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_df26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37242\,
            in2 => \_gnd_net_\,
            in3 => \N__37266\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_df28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34790\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33379\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33380\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49176\,
            ce => 'H',
            sr => \N__48426\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33340\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_2_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000110010"
        )
    port map (
            in0 => \N__33292\,
            in1 => \N__33243\,
            in2 => \N__33041\,
            in3 => \N__32934\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49168\,
            ce => \N__32899\,
            sr => \N__48431\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33603\,
            in2 => \N__33594\,
            in3 => \N__33784\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_12_14_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33585\,
            in2 => \N__33579\,
            in3 => \N__33999\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33570\,
            in2 => \N__33564\,
            in3 => \N__33974\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33555\,
            in2 => \N__33546\,
            in3 => \N__33954\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33537\,
            in2 => \N__33522\,
            in3 => \N__33936\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33918\,
            in1 => \N__33504\,
            in2 => \N__33513\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33498\,
            in2 => \N__33483\,
            in3 => \N__33900\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33471\,
            in2 => \N__33459\,
            in3 => \N__33882\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33768\,
            in2 => \N__33756\,
            in3 => \N__33861\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_12_15_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33747\,
            in2 => \N__33738\,
            in3 => \N__34173\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33717\,
            in2 => \N__33729\,
            in3 => \N__34155\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33711\,
            in2 => \N__33702\,
            in3 => \N__34137\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33681\,
            in2 => \N__33693\,
            in3 => \N__34119\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34101\,
            in1 => \N__33675\,
            in2 => \N__33660\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33651\,
            in2 => \N__33639\,
            in3 => \N__34083\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33630\,
            in2 => \N__33618\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33840\,
            in2 => \N__33831\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_16_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35463\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35286\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35253\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35217\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35181\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35172\,
            in2 => \N__35118\,
            in3 => \N__33807\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33804\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33791\,
            in2 => \N__34011\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_17_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34551\,
            in1 => \N__33998\,
            in2 => \_gnd_net_\,
            in3 => \N__33984\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__49143\,
            ce => 'H',
            sr => \N__48467\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__34555\,
            in1 => \N__33981\,
            in2 => \N__33975\,
            in3 => \N__33957\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__49143\,
            ce => 'H',
            sr => \N__48467\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34552\,
            in1 => \N__33953\,
            in2 => \_gnd_net_\,
            in3 => \N__33939\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__49143\,
            ce => 'H',
            sr => \N__48467\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34556\,
            in1 => \N__33935\,
            in2 => \_gnd_net_\,
            in3 => \N__33921\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__49143\,
            ce => 'H',
            sr => \N__48467\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34553\,
            in1 => \N__33917\,
            in2 => \_gnd_net_\,
            in3 => \N__33903\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__49143\,
            ce => 'H',
            sr => \N__48467\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34557\,
            in1 => \N__33899\,
            in2 => \_gnd_net_\,
            in3 => \N__33885\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__49143\,
            ce => 'H',
            sr => \N__48467\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34554\,
            in1 => \N__33878\,
            in2 => \_gnd_net_\,
            in3 => \N__33864\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__49143\,
            ce => 'H',
            sr => \N__48467\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34531\,
            in1 => \N__33857\,
            in2 => \_gnd_net_\,
            in3 => \N__33843\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_12_18_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__49138\,
            ce => 'H',
            sr => \N__48473\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34508\,
            in1 => \N__34172\,
            in2 => \_gnd_net_\,
            in3 => \N__34158\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__49138\,
            ce => 'H',
            sr => \N__48473\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34528\,
            in1 => \N__34154\,
            in2 => \_gnd_net_\,
            in3 => \N__34140\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__49138\,
            ce => 'H',
            sr => \N__48473\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34509\,
            in1 => \N__34136\,
            in2 => \_gnd_net_\,
            in3 => \N__34122\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__49138\,
            ce => 'H',
            sr => \N__48473\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34529\,
            in1 => \N__34118\,
            in2 => \_gnd_net_\,
            in3 => \N__34104\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__49138\,
            ce => 'H',
            sr => \N__48473\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34510\,
            in1 => \N__34100\,
            in2 => \_gnd_net_\,
            in3 => \N__34086\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__49138\,
            ce => 'H',
            sr => \N__48473\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34530\,
            in1 => \N__34082\,
            in2 => \_gnd_net_\,
            in3 => \N__34068\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__49138\,
            ce => 'H',
            sr => \N__48473\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34511\,
            in1 => \N__34055\,
            in2 => \_gnd_net_\,
            in3 => \N__34041\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__49138\,
            ce => 'H',
            sr => \N__48473\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34512\,
            in1 => \N__34028\,
            in2 => \_gnd_net_\,
            in3 => \N__34014\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_12_19_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__49133\,
            ce => 'H',
            sr => \N__48481\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34567\,
            in1 => \N__34246\,
            in2 => \_gnd_net_\,
            in3 => \N__34227\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__49133\,
            ce => 'H',
            sr => \N__48481\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34513\,
            in1 => \N__34217\,
            in2 => \_gnd_net_\,
            in3 => \N__34197\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \N__49133\,
            ce => 'H',
            sr => \N__48481\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34568\,
            in1 => \N__35475\,
            in2 => \_gnd_net_\,
            in3 => \N__34194\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \N__49133\,
            ce => 'H',
            sr => \N__48481\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34514\,
            in1 => \N__35487\,
            in2 => \_gnd_net_\,
            in3 => \N__34191\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\,
            clk => \N__49133\,
            ce => 'H',
            sr => \N__48481\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34569\,
            in1 => \N__35298\,
            in2 => \_gnd_net_\,
            in3 => \N__34188\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\,
            clk => \N__49133\,
            ce => 'H',
            sr => \N__48481\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34515\,
            in1 => \N__35310\,
            in2 => \_gnd_net_\,
            in3 => \N__34185\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\,
            clk => \N__49133\,
            ce => 'H',
            sr => \N__48481\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34570\,
            in1 => \N__35277\,
            in2 => \_gnd_net_\,
            in3 => \N__34182\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\,
            clk => \N__49133\,
            ce => 'H',
            sr => \N__48481\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34560\,
            in1 => \N__35265\,
            in2 => \_gnd_net_\,
            in3 => \N__34179\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_12_20_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\,
            clk => \N__49126\,
            ce => 'H',
            sr => \N__48493\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34571\,
            in1 => \N__35241\,
            in2 => \_gnd_net_\,
            in3 => \N__34176\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\,
            clk => \N__49126\,
            ce => 'H',
            sr => \N__48493\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34561\,
            in1 => \N__35229\,
            in2 => \_gnd_net_\,
            in3 => \N__34587\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\,
            clk => \N__49126\,
            ce => 'H',
            sr => \N__48493\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34572\,
            in1 => \N__35193\,
            in2 => \_gnd_net_\,
            in3 => \N__34584\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\,
            clk => \N__49126\,
            ce => 'H',
            sr => \N__48493\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34562\,
            in1 => \N__35205\,
            in2 => \_gnd_net_\,
            in3 => \N__34581\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\,
            clk => \N__49126\,
            ce => 'H',
            sr => \N__48493\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34573\,
            in1 => \N__35138\,
            in2 => \_gnd_net_\,
            in3 => \N__34578\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\,
            clk => \N__49126\,
            ce => 'H',
            sr => \N__48493\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34563\,
            in1 => \N__35164\,
            in2 => \_gnd_net_\,
            in3 => \N__34368\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49126\,
            ce => 'H',
            sr => \N__48493\
        );

    \phase_controller_inst1.stoper_tr.time_passed_RNI7NN7_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35668\,
            in2 => \_gnd_net_\,
            in3 => \N__35449\,
            lcout => \phase_controller_inst1.time_passed_RNI7NN7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_0_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__35450\,
            in1 => \N__34365\,
            in2 => \N__35571\,
            in3 => \N__35669\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49117\,
            ce => 'H',
            sr => \N__48513\
        );

    \phase_controller_inst1.T12_LC_12_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__34322\,
            in1 => \N__34311\,
            in2 => \_gnd_net_\,
            in3 => \N__35564\,
            lcout => \T12_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49110\,
            ce => 'H',
            sr => \N__48535\
        );

    \phase_controller_inst1.T01_LC_12_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__35645\,
            in1 => \N__34310\,
            in2 => \_gnd_net_\,
            in3 => \N__34265\,
            lcout => \T01_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49110\,
            ce => 'H',
            sr => \N__48535\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35813\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__35757\,
            in1 => \N__35814\,
            in2 => \_gnd_net_\,
            in3 => \N__35784\,
            lcout => \current_shift_inst.timer_s1.N_167_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40734\,
            in2 => \N__36020\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_13_7_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__49216\,
            ce => \N__44133\,
            sr => \N__48397\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44159\,
            in2 => \N__35994\,
            in3 => \N__34605\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__49216\,
            ce => \N__44133\,
            sr => \N__48397\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35960\,
            in2 => \N__36021\,
            in3 => \N__34602\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__49216\,
            ce => \N__44133\,
            sr => \N__48397\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35990\,
            in2 => \N__35939\,
            in3 => \N__34599\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__49216\,
            ce => \N__44133\,
            sr => \N__48397\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35961\,
            in2 => \N__35912\,
            in3 => \N__34596\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__49216\,
            ce => \N__44133\,
            sr => \N__48397\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35882\,
            in2 => \N__35940\,
            in3 => \N__34593\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__49216\,
            ce => \N__44133\,
            sr => \N__48397\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35845\,
            in2 => \N__35913\,
            in3 => \N__34590\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__49216\,
            ce => \N__44133\,
            sr => \N__48397\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36226\,
            in2 => \N__35883\,
            in3 => \N__34632\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__49216\,
            ce => \N__44133\,
            sr => \N__48397\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36206\,
            in2 => \N__35853\,
            in3 => \N__34629\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_13_8_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__49208\,
            ce => \N__44131\,
            sr => \N__48400\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36182\,
            in2 => \N__36237\,
            in3 => \N__34626\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__49208\,
            ce => \N__44131\,
            sr => \N__48400\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36207\,
            in2 => \N__36161\,
            in3 => \N__34623\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__49208\,
            ce => \N__44131\,
            sr => \N__48400\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36183\,
            in2 => \N__36131\,
            in3 => \N__34620\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__49208\,
            ce => \N__44131\,
            sr => \N__48400\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36104\,
            in2 => \N__36162\,
            in3 => \N__34617\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__49208\,
            ce => \N__44131\,
            sr => \N__48400\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36080\,
            in2 => \N__36132\,
            in3 => \N__34614\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__49208\,
            ce => \N__44131\,
            sr => \N__48400\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36105\,
            in2 => \N__36050\,
            in3 => \N__34611\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__49208\,
            ce => \N__44131\,
            sr => \N__48400\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36469\,
            in2 => \N__36084\,
            in3 => \N__34608\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__49208\,
            ce => \N__44131\,
            sr => \N__48400\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36449\,
            in2 => \N__36054\,
            in3 => \N__34662\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_13_9_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__49203\,
            ce => \N__44130\,
            sr => \N__48403\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36425\,
            in2 => \N__36480\,
            in3 => \N__34659\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__49203\,
            ce => \N__44130\,
            sr => \N__48403\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36450\,
            in2 => \N__36404\,
            in3 => \N__34656\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__49203\,
            ce => \N__44130\,
            sr => \N__48403\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36426\,
            in2 => \N__36374\,
            in3 => \N__34653\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__49203\,
            ce => \N__44130\,
            sr => \N__48403\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36347\,
            in2 => \N__36405\,
            in3 => \N__34650\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__49203\,
            ce => \N__44130\,
            sr => \N__48403\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36326\,
            in2 => \N__36375\,
            in3 => \N__34647\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__49203\,
            ce => \N__44130\,
            sr => \N__48403\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36348\,
            in2 => \N__36293\,
            in3 => \N__34644\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__49203\,
            ce => \N__44130\,
            sr => \N__48403\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36256\,
            in2 => \N__36327\,
            in3 => \N__34641\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__49203\,
            ce => \N__44130\,
            sr => \N__48403\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36297\,
            in2 => \N__36737\,
            in3 => \N__34638\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_13_10_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__49197\,
            ce => \N__44128\,
            sr => \N__48405\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36710\,
            in2 => \N__36267\,
            in3 => \N__34635\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__49197\,
            ce => \N__44128\,
            sr => \N__48405\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36690\,
            in2 => \N__36738\,
            in3 => \N__34695\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__49197\,
            ce => \N__44128\,
            sr => \N__48405\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36711\,
            in2 => \N__36546\,
            in3 => \N__34692\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__49197\,
            ce => \N__44128\,
            sr => \N__48405\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34689\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40204\,
            lcout => \current_shift_inst.un4_control_input_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40397\,
            lcout => \current_shift_inst.un4_control_input_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39851\,
            lcout => \current_shift_inst.un4_control_input_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36744\,
            in2 => \N__36791\,
            in3 => \N__36787\,
            lcout => \current_shift_inst.control_input_18\,
            ltout => OPEN,
            carryin => \bfn_13_11_0_\,
            carryout => \current_shift_inst.control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36804\,
            in2 => \_gnd_net_\,
            in3 => \N__34674\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_0\,
            carryout => \current_shift_inst.control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36768\,
            in2 => \_gnd_net_\,
            in3 => \N__34665\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_1\,
            carryout => \current_shift_inst.control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36762\,
            in2 => \_gnd_net_\,
            in3 => \N__34761\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_2\,
            carryout => \current_shift_inst.control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36756\,
            in2 => \_gnd_net_\,
            in3 => \N__34752\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_3\,
            carryout => \current_shift_inst.control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36750\,
            in2 => \_gnd_net_\,
            in3 => \N__34743\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_4\,
            carryout => \current_shift_inst.control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36954\,
            in2 => \_gnd_net_\,
            in3 => \N__34734\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_5\,
            carryout => \current_shift_inst.control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36948\,
            in2 => \_gnd_net_\,
            in3 => \N__34725\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_6\,
            carryout => \current_shift_inst.control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36939\,
            in2 => \_gnd_net_\,
            in3 => \N__34716\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_13_12_0_\,
            carryout => \current_shift_inst.control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36930\,
            in2 => \_gnd_net_\,
            in3 => \N__34707\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_8\,
            carryout => \current_shift_inst.control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36924\,
            in2 => \_gnd_net_\,
            in3 => \N__34698\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_9\,
            carryout => \current_shift_inst.control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38451\,
            in2 => \_gnd_net_\,
            in3 => \N__34806\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_10\,
            carryout => \current_shift_inst.control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36798\,
            in2 => \_gnd_net_\,
            in3 => \N__34797\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_11\,
            carryout => \current_shift_inst.control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38529\,
            in2 => \_gnd_net_\,
            in3 => \N__34794\,
            lcout => \current_shift_inst.control_input_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_11_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__40868\,
            in1 => \N__49596\,
            in2 => \N__42339\,
            in3 => \N__46823\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49179\,
            ce => \N__48802\,
            sr => \N__48427\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34889\,
            in2 => \_gnd_net_\,
            in3 => \N__34868\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIHOGI1_28_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110101"
        )
    port map (
            in0 => \N__34917\,
            in1 => \N__37458\,
            in2 => \N__37491\,
            in3 => \N__35337\,
            lcout => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIQU8A2_28_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34779\,
            in3 => \N__34890\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIQU8A2Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.running_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000101011111010"
        )
    port map (
            in0 => \N__34776\,
            in1 => \N__35322\,
            in2 => \N__34898\,
            in3 => \N__34919\,
            lcout => \phase_controller_inst2.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49170\,
            ce => 'H',
            sr => \N__48432\
        );

    \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__34916\,
            in1 => \N__34775\,
            in2 => \_gnd_net_\,
            in3 => \N__34964\,
            lcout => \phase_controller_inst2.stoper_tr.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.time_passed_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101000001010"
        )
    port map (
            in0 => \N__34984\,
            in1 => \N__35321\,
            in2 => \N__34899\,
            in3 => \N__34918\,
            lcout => \phase_controller_inst2.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49170\,
            ce => 'H',
            sr => \N__48432\
        );

    \phase_controller_inst2.stoper_tr.start_latched_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34965\,
            lcout => \phase_controller_inst2.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49170\,
            ce => 'H',
            sr => \N__48432\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__34891\,
            in1 => \N__34869\,
            in2 => \N__36918\,
            in3 => \N__50170\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49162\,
            ce => 'H',
            sr => \N__48443\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__40914\,
            in1 => \N__37563\,
            in2 => \_gnd_net_\,
            in3 => \N__37523\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49162\,
            ce => 'H',
            sr => \N__48443\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47490\,
            in2 => \N__34857\,
            in3 => \N__36913\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_13_16_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50436\,
            in2 => \N__34848\,
            in3 => \N__36888\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36861\,
            in1 => \N__46503\,
            in2 => \N__34839\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50295\,
            in2 => \N__34830\,
            in3 => \N__37119\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46518\,
            in2 => \N__34821\,
            in3 => \N__37101\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37083\,
            in1 => \N__35061\,
            in2 => \N__46668\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47502\,
            in2 => \N__35055\,
            in3 => \N__37065\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37047\,
            in1 => \N__45021\,
            in2 => \N__35046\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37029\,
            in1 => \N__38700\,
            in2 => \N__35037\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_13_17_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37380\,
            in2 => \N__35028\,
            in3 => \N__37011\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36990\,
            in1 => \N__38745\,
            in2 => \N__35019\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38733\,
            in2 => \N__35010\,
            in3 => \N__36972\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38439\,
            in2 => \N__34998\,
            in3 => \N__37218\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37200\,
            in1 => \N__37371\,
            in2 => \N__35100\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35091\,
            in2 => \N__37395\,
            in3 => \N__37182\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38829\,
            in2 => \N__38769\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38688\,
            in2 => \N__38625\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_18_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35106\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35496\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37401\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35085\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35073\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37483\,
            in2 => \N__37437\,
            in3 => \N__35328\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35325\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35309\,
            in2 => \_gnd_net_\,
            in3 => \N__35297\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_df22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__35276\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35264\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_df24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__35240\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35228\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_df26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35204\,
            in2 => \_gnd_net_\,
            in3 => \N__35192\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_df28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35163\,
            in2 => \_gnd_net_\,
            in3 => \N__35137\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37134\,
            in2 => \_gnd_net_\,
            in3 => \N__37152\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_df20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__37356\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37338\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_df22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__37652\,
            in1 => \N__37607\,
            in2 => \_gnd_net_\,
            in3 => \N__35352\,
            lcout => \phase_controller_inst1.stoper_tr.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__35353\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37653\,
            lcout => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__37737\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37719\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_df22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35486\,
            in2 => \_gnd_net_\,
            in3 => \N__35474\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_df20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101000011001100"
        )
    port map (
            in0 => \N__39456\,
            in1 => \N__35451\,
            in2 => \N__37659\,
            in3 => \N__37631\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49128\,
            ce => 'H',
            sr => \N__48494\
        );

    \phase_controller_inst1.stoper_tr.start_latched_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35355\,
            lcout => \phase_controller_inst1.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49128\,
            ce => 'H',
            sr => \N__48494\
        );

    \phase_controller_inst1.start_timer_tr_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101110101010"
        )
    port map (
            in0 => \N__35433\,
            in1 => \N__35423\,
            in2 => \N__35412\,
            in3 => \N__35354\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49128\,
            ce => 'H',
            sr => \N__48494\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37751\,
            in2 => \_gnd_net_\,
            in3 => \N__37766\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_df20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37818\,
            in2 => \_gnd_net_\,
            in3 => \N__37832\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_df24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNII51H_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__35800\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35775\,
            lcout => \current_shift_inst.timer_s1.N_166_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__35779\,
            in1 => \N__35750\,
            in2 => \_gnd_net_\,
            in3 => \N__35806\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49119\,
            ce => 'H',
            sr => \N__48514\
        );

    \current_shift_inst.stop_timer_s1_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101100"
        )
    port map (
            in0 => \N__35749\,
            in1 => \N__35780\,
            in2 => \N__35652\,
            in3 => \N__35723\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49119\,
            ce => 'H',
            sr => \N__48514\
        );

    \current_shift_inst.start_timer_s1_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__35716\,
            in1 => \N__35748\,
            in2 => \_gnd_net_\,
            in3 => \N__35651\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49116\,
            ce => 'H',
            sr => \N__48521\
        );

    \phase_controller_inst1.S1_LC_13_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35650\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49114\,
            ce => 'H',
            sr => \N__48527\
        );

    \phase_controller_inst1.T23_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__35690\,
            in1 => \N__35569\,
            in2 => \_gnd_net_\,
            in3 => \N__35678\,
            lcout => \T23_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49113\,
            ce => 'H',
            sr => \N__48532\
        );

    \phase_controller_inst1.T45_LC_13_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__35679\,
            in1 => \N__35582\,
            in2 => \_gnd_net_\,
            in3 => \N__35649\,
            lcout => \T45_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49113\,
            ce => 'H',
            sr => \N__48532\
        );

    \phase_controller_inst1.S2_LC_13_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35570\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49111\,
            ce => 'H',
            sr => \N__48536\
        );

    \current_shift_inst.timer_s1.counter_0_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36667\,
            in1 => \N__40726\,
            in2 => \_gnd_net_\,
            in3 => \N__35499\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_14_5_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__49232\,
            ce => \N__36523\,
            sr => \N__48393\
        );

    \current_shift_inst.timer_s1.counter_1_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36629\,
            in1 => \N__44155\,
            in2 => \_gnd_net_\,
            in3 => \N__36024\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__49232\,
            ce => \N__36523\,
            sr => \N__48393\
        );

    \current_shift_inst.timer_s1.counter_2_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36668\,
            in1 => \N__36013\,
            in2 => \_gnd_net_\,
            in3 => \N__35997\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__49232\,
            ce => \N__36523\,
            sr => \N__48393\
        );

    \current_shift_inst.timer_s1.counter_3_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36630\,
            in1 => \N__35986\,
            in2 => \_gnd_net_\,
            in3 => \N__35964\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__49232\,
            ce => \N__36523\,
            sr => \N__48393\
        );

    \current_shift_inst.timer_s1.counter_4_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36669\,
            in1 => \N__35959\,
            in2 => \_gnd_net_\,
            in3 => \N__35943\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__49232\,
            ce => \N__36523\,
            sr => \N__48393\
        );

    \current_shift_inst.timer_s1.counter_5_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36631\,
            in1 => \N__35932\,
            in2 => \_gnd_net_\,
            in3 => \N__35916\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__49232\,
            ce => \N__36523\,
            sr => \N__48393\
        );

    \current_shift_inst.timer_s1.counter_6_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36670\,
            in1 => \N__35900\,
            in2 => \_gnd_net_\,
            in3 => \N__35886\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__49232\,
            ce => \N__36523\,
            sr => \N__48393\
        );

    \current_shift_inst.timer_s1.counter_7_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36632\,
            in1 => \N__35875\,
            in2 => \_gnd_net_\,
            in3 => \N__35856\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__49232\,
            ce => \N__36523\,
            sr => \N__48393\
        );

    \current_shift_inst.timer_s1.counter_8_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36666\,
            in1 => \N__35849\,
            in2 => \_gnd_net_\,
            in3 => \N__35829\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_14_6_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__49227\,
            ce => \N__36524\,
            sr => \N__48394\
        );

    \current_shift_inst.timer_s1.counter_9_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36636\,
            in1 => \N__36230\,
            in2 => \_gnd_net_\,
            in3 => \N__36210\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__49227\,
            ce => \N__36524\,
            sr => \N__48394\
        );

    \current_shift_inst.timer_s1.counter_10_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36663\,
            in1 => \N__36200\,
            in2 => \_gnd_net_\,
            in3 => \N__36186\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__49227\,
            ce => \N__36524\,
            sr => \N__48394\
        );

    \current_shift_inst.timer_s1.counter_11_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36633\,
            in1 => \N__36181\,
            in2 => \_gnd_net_\,
            in3 => \N__36165\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__49227\,
            ce => \N__36524\,
            sr => \N__48394\
        );

    \current_shift_inst.timer_s1.counter_12_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36664\,
            in1 => \N__36149\,
            in2 => \_gnd_net_\,
            in3 => \N__36135\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__49227\,
            ce => \N__36524\,
            sr => \N__48394\
        );

    \current_shift_inst.timer_s1.counter_13_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36634\,
            in1 => \N__36124\,
            in2 => \_gnd_net_\,
            in3 => \N__36108\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__49227\,
            ce => \N__36524\,
            sr => \N__48394\
        );

    \current_shift_inst.timer_s1.counter_14_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36665\,
            in1 => \N__36103\,
            in2 => \_gnd_net_\,
            in3 => \N__36087\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__49227\,
            ce => \N__36524\,
            sr => \N__48394\
        );

    \current_shift_inst.timer_s1.counter_15_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36635\,
            in1 => \N__36073\,
            in2 => \_gnd_net_\,
            in3 => \N__36057\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__49227\,
            ce => \N__36524\,
            sr => \N__48394\
        );

    \current_shift_inst.timer_s1.counter_16_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36646\,
            in1 => \N__36049\,
            in2 => \_gnd_net_\,
            in3 => \N__36027\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_14_7_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__49221\,
            ce => \N__36516\,
            sr => \N__48395\
        );

    \current_shift_inst.timer_s1.counter_17_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36654\,
            in1 => \N__36473\,
            in2 => \_gnd_net_\,
            in3 => \N__36453\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__49221\,
            ce => \N__36516\,
            sr => \N__48395\
        );

    \current_shift_inst.timer_s1.counter_18_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36647\,
            in1 => \N__36443\,
            in2 => \_gnd_net_\,
            in3 => \N__36429\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__49221\,
            ce => \N__36516\,
            sr => \N__48395\
        );

    \current_shift_inst.timer_s1.counter_19_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36655\,
            in1 => \N__36424\,
            in2 => \_gnd_net_\,
            in3 => \N__36408\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__49221\,
            ce => \N__36516\,
            sr => \N__48395\
        );

    \current_shift_inst.timer_s1.counter_20_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36648\,
            in1 => \N__36392\,
            in2 => \_gnd_net_\,
            in3 => \N__36378\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__49221\,
            ce => \N__36516\,
            sr => \N__48395\
        );

    \current_shift_inst.timer_s1.counter_21_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36656\,
            in1 => \N__36367\,
            in2 => \_gnd_net_\,
            in3 => \N__36351\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__49221\,
            ce => \N__36516\,
            sr => \N__48395\
        );

    \current_shift_inst.timer_s1.counter_22_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36649\,
            in1 => \N__36346\,
            in2 => \_gnd_net_\,
            in3 => \N__36330\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__49221\,
            ce => \N__36516\,
            sr => \N__48395\
        );

    \current_shift_inst.timer_s1.counter_23_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36657\,
            in1 => \N__36319\,
            in2 => \_gnd_net_\,
            in3 => \N__36300\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__49221\,
            ce => \N__36516\,
            sr => \N__48395\
        );

    \current_shift_inst.timer_s1.counter_24_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36650\,
            in1 => \N__36292\,
            in2 => \_gnd_net_\,
            in3 => \N__36270\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_14_8_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__49217\,
            ce => \N__36528\,
            sr => \N__48398\
        );

    \current_shift_inst.timer_s1.counter_25_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36671\,
            in1 => \N__36260\,
            in2 => \_gnd_net_\,
            in3 => \N__36240\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__49217\,
            ce => \N__36528\,
            sr => \N__48398\
        );

    \current_shift_inst.timer_s1.counter_26_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36651\,
            in1 => \N__36730\,
            in2 => \_gnd_net_\,
            in3 => \N__36714\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__49217\,
            ce => \N__36528\,
            sr => \N__48398\
        );

    \current_shift_inst.timer_s1.counter_27_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36672\,
            in1 => \N__36709\,
            in2 => \_gnd_net_\,
            in3 => \N__36693\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__49217\,
            ce => \N__36528\,
            sr => \N__48398\
        );

    \current_shift_inst.timer_s1.counter_28_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36652\,
            in1 => \N__36689\,
            in2 => \_gnd_net_\,
            in3 => \N__36675\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__49217\,
            ce => \N__36528\,
            sr => \N__48398\
        );

    \current_shift_inst.timer_s1.counter_29_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__36542\,
            in1 => \N__36653\,
            in2 => \_gnd_net_\,
            in3 => \N__36549\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49217\,
            ce => \N__36528\,
            sr => \N__48398\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39791\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44652\,
            lcout => \current_shift_inst.un4_control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__44052\,
            in1 => \N__41064\,
            in2 => \_gnd_net_\,
            in3 => \N__40666\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\,
            ltout => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_inv_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__38162\,
            in1 => \_gnd_net_\,
            in2 => \N__36486\,
            in3 => \N__36813\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_31\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38163\,
            in2 => \N__36483\,
            in3 => \N__41616\,
            lcout => \current_shift_inst.un38_control_input_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46162\,
            lcout => \current_shift_inst.un4_control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44053\,
            in1 => \_gnd_net_\,
            in2 => \N__41761\,
            in3 => \N__41735\,
            lcout => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41752\,
            lcout => \current_shift_inst.un4_control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__40244\,
            in1 => \N__45443\,
            in2 => \_gnd_net_\,
            in3 => \N__41473\,
            lcout => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40243\,
            lcout => \current_shift_inst.un4_control_input_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__43414\,
            in1 => \N__44036\,
            in2 => \_gnd_net_\,
            in3 => \N__43385\,
            lcout => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43413\,
            lcout => \current_shift_inst.un4_control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__39683\,
            in1 => \N__44037\,
            in2 => \_gnd_net_\,
            in3 => \N__41157\,
            lcout => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39682\,
            lcout => \current_shift_inst.un4_control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__41886\,
            in1 => \N__38418\,
            in2 => \_gnd_net_\,
            in3 => \N__38494\,
            lcout => \current_shift_inst.control_input_axb_0\,
            ltout => \current_shift_inst.control_input_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_0_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36843\,
            in3 => \N__36792\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49204\,
            ce => 'H',
            sr => \N__48404\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39973\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49198\,
            ce => \N__44129\,
            sr => \N__48406\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__38403\,
            in1 => \N__41862\,
            in2 => \_gnd_net_\,
            in3 => \N__38496\,
            lcout => \current_shift_inst.control_input_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38514\,
            lcout => \current_shift_inst.control_input_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38495\,
            lcout => \current_shift_inst.N_1460_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__38497\,
            in1 => \N__38391\,
            in2 => \_gnd_net_\,
            in3 => \N__42063\,
            lcout => \current_shift_inst.control_input_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__38379\,
            in1 => \N__42048\,
            in2 => \_gnd_net_\,
            in3 => \N__38498\,
            lcout => \current_shift_inst.control_input_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__38367\,
            in1 => \N__38512\,
            in2 => \_gnd_net_\,
            in3 => \N__42021\,
            lcout => \current_shift_inst.control_input_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__38513\,
            in1 => \N__42000\,
            in2 => \_gnd_net_\,
            in3 => \N__38601\,
            lcout => \current_shift_inst.control_input_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100100111"
        )
    port map (
            in0 => \N__38499\,
            in1 => \N__38589\,
            in2 => \N__41976\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.control_input_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__41946\,
            in1 => \N__38577\,
            in2 => \_gnd_net_\,
            in3 => \N__38518\,
            lcout => \current_shift_inst.control_input_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__38519\,
            in1 => \N__41916\,
            in2 => \_gnd_net_\,
            in3 => \N__38565\,
            lcout => \current_shift_inst.control_input_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__41901\,
            in1 => \N__38553\,
            in2 => \_gnd_net_\,
            in3 => \N__38520\,
            lcout => \current_shift_inst.control_input_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__38521\,
            in1 => \N__42300\,
            in2 => \_gnd_net_\,
            in3 => \N__38541\,
            lcout => \current_shift_inst.control_input_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36914\,
            in2 => \N__36897\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50260\,
            in1 => \N__36887\,
            in2 => \_gnd_net_\,
            in3 => \N__36873\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__49180\,
            ce => 'H',
            sr => \N__48428\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__50277\,
            in1 => \N__36860\,
            in2 => \N__36870\,
            in3 => \N__36846\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__49180\,
            ce => 'H',
            sr => \N__48428\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50261\,
            in1 => \N__37118\,
            in2 => \_gnd_net_\,
            in3 => \N__37104\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__49180\,
            ce => 'H',
            sr => \N__48428\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50278\,
            in1 => \N__37100\,
            in2 => \_gnd_net_\,
            in3 => \N__37086\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__49180\,
            ce => 'H',
            sr => \N__48428\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50262\,
            in1 => \N__37082\,
            in2 => \_gnd_net_\,
            in3 => \N__37068\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__49180\,
            ce => 'H',
            sr => \N__48428\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50279\,
            in1 => \N__37064\,
            in2 => \_gnd_net_\,
            in3 => \N__37050\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__49180\,
            ce => 'H',
            sr => \N__48428\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50263\,
            in1 => \N__37046\,
            in2 => \_gnd_net_\,
            in3 => \N__37032\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__49180\,
            ce => 'H',
            sr => \N__48428\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50163\,
            in1 => \N__37028\,
            in2 => \_gnd_net_\,
            in3 => \N__37014\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__49171\,
            ce => 'H',
            sr => \N__48433\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50156\,
            in1 => \N__37007\,
            in2 => \_gnd_net_\,
            in3 => \N__36993\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__49171\,
            ce => 'H',
            sr => \N__48433\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50160\,
            in1 => \N__36989\,
            in2 => \_gnd_net_\,
            in3 => \N__36975\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__49171\,
            ce => 'H',
            sr => \N__48433\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50157\,
            in1 => \N__36971\,
            in2 => \_gnd_net_\,
            in3 => \N__36957\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__49171\,
            ce => 'H',
            sr => \N__48433\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50161\,
            in1 => \N__37217\,
            in2 => \_gnd_net_\,
            in3 => \N__37203\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__49171\,
            ce => 'H',
            sr => \N__48433\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50158\,
            in1 => \N__37199\,
            in2 => \_gnd_net_\,
            in3 => \N__37185\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__49171\,
            ce => 'H',
            sr => \N__48433\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50162\,
            in1 => \N__37181\,
            in2 => \_gnd_net_\,
            in3 => \N__37167\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__49171\,
            ce => 'H',
            sr => \N__48433\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50159\,
            in1 => \N__38812\,
            in2 => \_gnd_net_\,
            in3 => \N__37164\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__49171\,
            ce => 'H',
            sr => \N__48433\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50237\,
            in1 => \N__38784\,
            in2 => \_gnd_net_\,
            in3 => \N__37161\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__49163\,
            ce => 'H',
            sr => \N__48444\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50245\,
            in1 => \N__38660\,
            in2 => \_gnd_net_\,
            in3 => \N__37158\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__49163\,
            ce => 'H',
            sr => \N__48444\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50238\,
            in1 => \N__38643\,
            in2 => \_gnd_net_\,
            in3 => \N__37155\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \N__49163\,
            ce => 'H',
            sr => \N__48444\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50246\,
            in1 => \N__37151\,
            in2 => \_gnd_net_\,
            in3 => \N__37137\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \N__49163\,
            ce => 'H',
            sr => \N__48444\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50239\,
            in1 => \N__37133\,
            in2 => \_gnd_net_\,
            in3 => \N__37359\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\,
            clk => \N__49163\,
            ce => 'H',
            sr => \N__48444\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50247\,
            in1 => \N__37355\,
            in2 => \_gnd_net_\,
            in3 => \N__37341\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\,
            clk => \N__49163\,
            ce => 'H',
            sr => \N__48444\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50240\,
            in1 => \N__37337\,
            in2 => \_gnd_net_\,
            in3 => \N__37323\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\,
            clk => \N__49163\,
            ce => 'H',
            sr => \N__48444\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50248\,
            in1 => \N__37427\,
            in2 => \_gnd_net_\,
            in3 => \N__37320\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\,
            clk => \N__49163\,
            ce => 'H',
            sr => \N__48444\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50241\,
            in1 => \N__37413\,
            in2 => \_gnd_net_\,
            in3 => \N__37317\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\,
            clk => \N__49156\,
            ce => 'H',
            sr => \N__48455\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50249\,
            in1 => \N__37307\,
            in2 => \_gnd_net_\,
            in3 => \N__37293\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\,
            clk => \N__49156\,
            ce => 'H',
            sr => \N__48455\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50242\,
            in1 => \N__37283\,
            in2 => \_gnd_net_\,
            in3 => \N__37269\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\,
            clk => \N__49156\,
            ce => 'H',
            sr => \N__48455\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50250\,
            in1 => \N__37259\,
            in2 => \_gnd_net_\,
            in3 => \N__37245\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\,
            clk => \N__49156\,
            ce => 'H',
            sr => \N__48455\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50243\,
            in1 => \N__37235\,
            in2 => \_gnd_net_\,
            in3 => \N__37221\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\,
            clk => \N__49156\,
            ce => 'H',
            sr => \N__48455\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50251\,
            in1 => \N__37457\,
            in2 => \_gnd_net_\,
            in3 => \N__37569\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\,
            clk => \N__49156\,
            ce => 'H',
            sr => \N__48455\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50244\,
            in1 => \N__37484\,
            in2 => \_gnd_net_\,
            in3 => \N__37566\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49156\,
            ce => 'H',
            sr => \N__48455\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__37559\,
            in1 => \N__40921\,
            in2 => \_gnd_net_\,
            in3 => \N__37527\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_396_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__37482\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37456\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__37428\,
            in1 => \N__37412\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_df24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_15_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__42404\,
            in1 => \N__49566\,
            in2 => \N__46890\,
            in3 => \N__46817\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49146\,
            ce => \N__50259\,
            sr => \N__48468\
        );

    \phase_controller_inst2.stoper_tr.target_time_10_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__40866\,
            in1 => \N__49564\,
            in2 => \N__42266\,
            in3 => \N__46815\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49146\,
            ce => \N__50259\,
            sr => \N__48468\
        );

    \phase_controller_inst2.stoper_tr.target_time_14_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__40867\,
            in1 => \N__49565\,
            in2 => \N__42180\,
            in3 => \N__46816\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49146\,
            ce => \N__50259\,
            sr => \N__48468\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNID27N1_28_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011111111"
        )
    port map (
            in0 => \N__39471\,
            in1 => \N__39359\,
            in2 => \N__39330\,
            in3 => \N__37654\,
            lcout => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37625\,
            in2 => \N__37671\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIJF7V2_28_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__37626\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37667\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIJF7V2Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__37668\,
            in1 => \N__37630\,
            in2 => \N__38957\,
            in3 => \N__48666\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49140\,
            ce => 'H',
            sr => \N__48474\
        );

    \phase_controller_inst1.stoper_tr.running_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011111100110000"
        )
    port map (
            in0 => \N__39455\,
            in1 => \N__37655\,
            in2 => \N__37632\,
            in3 => \N__37608\,
            lcout => \phase_controller_inst1.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49140\,
            ce => 'H',
            sr => \N__48474\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37596\,
            in2 => \N__38958\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_21_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48667\,
            in1 => \N__38922\,
            in2 => \_gnd_net_\,
            in3 => \N__37590\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__49135\,
            ce => 'H',
            sr => \N__48482\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__48753\,
            in1 => \N__38901\,
            in2 => \N__37587\,
            in3 => \N__37578\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__49135\,
            ce => 'H',
            sr => \N__48482\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48668\,
            in1 => \N__38880\,
            in2 => \_gnd_net_\,
            in3 => \N__37575\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__49135\,
            ce => 'H',
            sr => \N__48482\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48754\,
            in1 => \N__38859\,
            in2 => \_gnd_net_\,
            in3 => \N__37572\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__49135\,
            ce => 'H',
            sr => \N__48482\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48669\,
            in1 => \N__39167\,
            in2 => \_gnd_net_\,
            in3 => \N__37698\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__49135\,
            ce => 'H',
            sr => \N__48482\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48755\,
            in1 => \N__39135\,
            in2 => \_gnd_net_\,
            in3 => \N__37695\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__49135\,
            ce => 'H',
            sr => \N__48482\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48670\,
            in1 => \N__39117\,
            in2 => \_gnd_net_\,
            in3 => \N__37692\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__49135\,
            ce => 'H',
            sr => \N__48482\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48763\,
            in1 => \N__39090\,
            in2 => \_gnd_net_\,
            in3 => \N__37689\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_14_22_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__49129\,
            ce => 'H',
            sr => \N__48495\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48749\,
            in1 => \N__39069\,
            in2 => \_gnd_net_\,
            in3 => \N__37686\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__49129\,
            ce => 'H',
            sr => \N__48495\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48760\,
            in1 => \N__39021\,
            in2 => \_gnd_net_\,
            in3 => \N__37683\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__49129\,
            ce => 'H',
            sr => \N__48495\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48750\,
            in1 => \N__39000\,
            in2 => \_gnd_net_\,
            in3 => \N__37680\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__49129\,
            ce => 'H',
            sr => \N__48495\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48761\,
            in1 => \N__38979\,
            in2 => \_gnd_net_\,
            in3 => \N__37677\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__49129\,
            ce => 'H',
            sr => \N__48495\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48751\,
            in1 => \N__39249\,
            in2 => \_gnd_net_\,
            in3 => \N__37674\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__49129\,
            ce => 'H',
            sr => \N__48495\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48762\,
            in1 => \N__39216\,
            in2 => \_gnd_net_\,
            in3 => \N__37782\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__49129\,
            ce => 'H',
            sr => \N__48495\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48752\,
            in1 => \N__39424\,
            in2 => \_gnd_net_\,
            in3 => \N__37779\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__49129\,
            ce => 'H',
            sr => \N__48495\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48745\,
            in1 => \N__39408\,
            in2 => \_gnd_net_\,
            in3 => \N__37776\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_14_23_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__49124\,
            ce => 'H',
            sr => \N__48505\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48812\,
            in1 => \N__39561\,
            in2 => \_gnd_net_\,
            in3 => \N__37773\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__49124\,
            ce => 'H',
            sr => \N__48505\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48746\,
            in1 => \N__39579\,
            in2 => \_gnd_net_\,
            in3 => \N__37770\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \N__49124\,
            ce => 'H',
            sr => \N__48505\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48813\,
            in1 => \N__37767\,
            in2 => \_gnd_net_\,
            in3 => \N__37755\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \N__49124\,
            ce => 'H',
            sr => \N__48505\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48747\,
            in1 => \N__37752\,
            in2 => \_gnd_net_\,
            in3 => \N__37740\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\,
            clk => \N__49124\,
            ce => 'H',
            sr => \N__48505\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48814\,
            in1 => \N__37736\,
            in2 => \_gnd_net_\,
            in3 => \N__37722\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\,
            clk => \N__49124\,
            ce => 'H',
            sr => \N__48505\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48748\,
            in1 => \N__37715\,
            in2 => \_gnd_net_\,
            in3 => \N__37701\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\,
            clk => \N__49124\,
            ce => 'H',
            sr => \N__48505\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48815\,
            in1 => \N__37833\,
            in2 => \_gnd_net_\,
            in3 => \N__37821\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\,
            clk => \N__49124\,
            ce => 'H',
            sr => \N__48505\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_14_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48756\,
            in1 => \N__37817\,
            in2 => \_gnd_net_\,
            in3 => \N__37803\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_14_24_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\,
            clk => \N__49120\,
            ce => 'H',
            sr => \N__48515\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48805\,
            in1 => \N__39612\,
            in2 => \_gnd_net_\,
            in3 => \N__37800\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\,
            clk => \N__49120\,
            ce => 'H',
            sr => \N__48515\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_14_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48757\,
            in1 => \N__39600\,
            in2 => \_gnd_net_\,
            in3 => \N__37797\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\,
            clk => \N__49120\,
            ce => 'H',
            sr => \N__48515\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48806\,
            in1 => \N__39279\,
            in2 => \_gnd_net_\,
            in3 => \N__37794\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\,
            clk => \N__49120\,
            ce => 'H',
            sr => \N__48515\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48758\,
            in1 => \N__39291\,
            in2 => \_gnd_net_\,
            in3 => \N__37791\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\,
            clk => \N__49120\,
            ce => 'H',
            sr => \N__48515\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_14_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48807\,
            in1 => \N__39323\,
            in2 => \_gnd_net_\,
            in3 => \N__37788\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\,
            clk => \N__49120\,
            ce => 'H',
            sr => \N__48515\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_14_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48759\,
            in1 => \N__39358\,
            in2 => \_gnd_net_\,
            in3 => \N__37785\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49120\,
            ce => 'H',
            sr => \N__48515\
        );

    \CONSTANT_ONE_LUT4_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37915\,
            in2 => \_gnd_net_\,
            in3 => \N__44580\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37895\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__45885\,
            in1 => \N__45421\,
            in2 => \N__44676\,
            in3 => \N__44634\,
            lcout => \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__45418\,
            in1 => \N__45886\,
            in2 => \N__40950\,
            in3 => \N__39525\,
            lcout => \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__45884\,
            in1 => \N__45420\,
            in2 => \N__43740\,
            in3 => \N__43775\,
            lcout => \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45419\,
            in1 => \N__45887\,
            in2 => \N__41103\,
            in3 => \N__41208\,
            lcout => \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43774\,
            lcout => \current_shift_inst.un4_control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__43302\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__41088\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40692\,
            lcout => \current_shift_inst.un4_control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110001101"
        )
    port map (
            in0 => \N__45422\,
            in1 => \N__41256\,
            in2 => \N__40702\,
            in3 => \N__45882\,
            lcout => \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__45883\,
            in1 => \N__45423\,
            in2 => \N__43312\,
            in3 => \N__43334\,
            lcout => \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40113\,
            lcout => \current_shift_inst.un4_control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39514\,
            lcout => \current_shift_inst.un4_control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__41089\,
            in1 => \N__44055\,
            in2 => \_gnd_net_\,
            in3 => \N__41204\,
            lcout => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43841\,
            in2 => \N__37935\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_8_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38057\,
            in2 => \N__43899\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_0\,
            carryout => \current_shift_inst.un10_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39531\,
            in2 => \N__38138\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_1\,
            carryout => \current_shift_inst.un10_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38061\,
            in2 => \N__39480\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_2\,
            carryout => \current_shift_inst.un10_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39495\,
            in2 => \N__38139\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_3\,
            carryout => \current_shift_inst.un10_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38065\,
            in2 => \N__39489\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_4\,
            carryout => \current_shift_inst.un10_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37965\,
            in2 => \N__38140\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_5\,
            carryout => \current_shift_inst.un10_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38069\,
            in2 => \N__37956\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_6\,
            carryout => \current_shift_inst.un10_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38082\,
            in2 => \N__39624\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_9_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37947\,
            in2 => \N__38144\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_8\,
            carryout => \current_shift_inst.un10_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38070\,
            in2 => \N__39774\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_9\,
            carryout => \current_shift_inst.un10_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37941\,
            in2 => \N__38141\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_10\,
            carryout => \current_shift_inst.un10_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38074\,
            in2 => \N__39654\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_11\,
            carryout => \current_shift_inst.un10_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39636\,
            in2 => \N__38142\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_12\,
            carryout => \current_shift_inst.un10_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38078\,
            in2 => \N__39645\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_13\,
            carryout => \current_shift_inst.un10_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39630\,
            in2 => \N__38143\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_14\,
            carryout => \current_shift_inst.un10_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38086\,
            in2 => \N__39723\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_10_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39714\,
            in2 => \N__38145\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_16\,
            carryout => \current_shift_inst.un10_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38090\,
            in2 => \N__39756\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_17\,
            carryout => \current_shift_inst.un10_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39702\,
            in2 => \N__38146\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_18\,
            carryout => \current_shift_inst.un10_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38094\,
            in2 => \N__39732\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_19\,
            carryout => \current_shift_inst.un10_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39780\,
            in2 => \N__38147\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_20\,
            carryout => \current_shift_inst.un10_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38098\,
            in2 => \N__39765\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_21\,
            carryout => \current_shift_inst.un10_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39708\,
            in2 => \N__38148\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_22\,
            carryout => \current_shift_inst.un10_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38149\,
            in2 => \N__40143\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_11_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38289\,
            in2 => \N__38192\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_24\,
            carryout => \current_shift_inst.un10_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38153\,
            in2 => \N__40083\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_25\,
            carryout => \current_shift_inst.un10_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39993\,
            in2 => \N__38193\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_26\,
            carryout => \current_shift_inst.un10_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38157\,
            in2 => \N__39840\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_27\,
            carryout => \current_shift_inst.un10_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39888\,
            in2 => \N__38194\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_28\,
            carryout => \current_shift_inst.un10_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38161\,
            in2 => \N__43884\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_29\,
            carryout => \current_shift_inst.un10_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45393\,
            in2 => \_gnd_net_\,
            in3 => \N__38328\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41633\,
            in2 => \N__39924\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_12_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44086\,
            in2 => \N__43266\,
            in3 => \N__43842\,
            lcout => \current_shift_inst.un38_control_input_5_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__43843\,
            in1 => \N__45583\,
            in2 => \N__39960\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un38_control_input_5_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40089\,
            in2 => \N__45748\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45587\,
            in2 => \N__38325\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38313\,
            in2 => \N__45749\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45591\,
            in2 => \N__39906\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38301\,
            in2 => \N__45750\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45637\,
            in2 => \N__38355\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_13_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39696\,
            in2 => \N__45840\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45641\,
            in2 => \N__40329\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40335\,
            in2 => \N__45841\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45645\,
            in2 => \N__43626\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40149\,
            in2 => \N__45842\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45649\,
            in2 => \N__39897\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38340\,
            in2 => \N__45843\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45719\,
            in2 => \N__40170\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_14_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40347\,
            in2 => \N__45900\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45723\,
            in2 => \N__40002\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38427\,
            in2 => \N__45901\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45727\,
            in2 => \N__39747\,
            in3 => \N__38406\,
            lcout => \current_shift_inst.un38_control_input_0_s0_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39819\,
            in2 => \N__45902\,
            in3 => \N__38394\,
            lcout => \current_shift_inst.un38_control_input_0_s0_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45731\,
            in2 => \N__46215\,
            in3 => \N__38382\,
            lcout => \current_shift_inst.un38_control_input_0_s0_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40341\,
            in2 => \N__45903\,
            in3 => \N__38370\,
            lcout => \current_shift_inst.un38_control_input_0_s0_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45735\,
            in2 => \N__40179\,
            in3 => \N__38358\,
            lcout => \current_shift_inst.un38_control_input_0_s0_24\,
            ltout => OPEN,
            carryin => \bfn_15_15_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40230\,
            in2 => \N__45904\,
            in3 => \N__38592\,
            lcout => \current_shift_inst.un38_control_input_0_s0_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45739\,
            in2 => \N__40188\,
            in3 => \N__38580\,
            lcout => \current_shift_inst.un38_control_input_0_s0_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40386\,
            in2 => \N__45905\,
            in3 => \N__38568\,
            lcout => \current_shift_inst.un38_control_input_0_s0_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45743\,
            in2 => \N__39882\,
            in3 => \N__38556\,
            lcout => \current_shift_inst.un38_control_input_0_s0_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40161\,
            in2 => \N__45906\,
            in3 => \N__38544\,
            lcout => \current_shift_inst.un38_control_input_0_s0_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45747\,
            in2 => \N__43800\,
            in3 => \N__38532\,
            lcout => \current_shift_inst.un38_control_input_0_s0_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101101000111"
        )
    port map (
            in0 => \N__39831\,
            in1 => \N__38528\,
            in2 => \N__42282\,
            in3 => \N__38454\,
            lcout => \current_shift_inst.control_input_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_13_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__49468\,
            in1 => \N__42203\,
            in2 => \N__40860\,
            in3 => \N__46752\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49172\,
            ce => \N__50285\,
            sr => \N__48434\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_a2_10_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__46878\,
            in1 => \N__42397\,
            in2 => \_gnd_net_\,
            in3 => \N__42170\,
            lcout => \phase_controller_inst1.stoper_tr.N_242\,
            ltout => \phase_controller_inst1.stoper_tr.N_242_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_11_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__49467\,
            in1 => \N__42334\,
            in2 => \N__38748\,
            in3 => \N__46751\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49172\,
            ce => \N__50285\,
            sr => \N__48434\
        );

    \phase_controller_inst2.stoper_tr.target_time_12_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__46749\,
            in1 => \N__42229\,
            in2 => \N__40859\,
            in3 => \N__49469\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49172\,
            ce => \N__50285\,
            sr => \N__48434\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1_9_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111110"
        )
    port map (
            in0 => \N__49466\,
            in1 => \N__38715\,
            in2 => \N__42489\,
            in3 => \N__46748\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_9_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__46750\,
            in1 => \N__40838\,
            in2 => \N__38703\,
            in3 => \N__42123\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49172\,
            ce => \N__50285\,
            sr => \N__48434\
        );

    \phase_controller_inst2.stoper_tr.target_time_19_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111100001010"
        )
    port map (
            in0 => \N__47784\,
            in1 => \_gnd_net_\,
            in2 => \N__49598\,
            in3 => \N__46765\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49164\,
            ce => \N__50276\,
            sr => \N__48445\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__38609\,
            in1 => \N__38641\,
            in2 => \N__38676\,
            in3 => \N__38659\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__38672\,
            in1 => \N__38610\,
            in2 => \N__38661\,
            in3 => \N__38642\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_18_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49567\,
            in2 => \N__46807\,
            in3 => \N__42556\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49164\,
            ce => \N__50276\,
            sr => \N__48445\
        );

    \phase_controller_inst2.stoper_tr.target_time_17_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111100001010"
        )
    port map (
            in0 => \N__42517\,
            in1 => \_gnd_net_\,
            in2 => \N__49597\,
            in3 => \N__46764\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49164\,
            ce => \N__50276\,
            sr => \N__48445\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011101010001"
        )
    port map (
            in0 => \N__38782\,
            in1 => \N__38814\,
            in2 => \N__46446\,
            in3 => \N__38792\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__38813\,
            in1 => \N__46445\,
            in2 => \N__38796\,
            in3 => \N__38783\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110010"
        )
    port map (
            in0 => \N__42560\,
            in1 => \N__49860\,
            in2 => \N__47644\,
            in3 => \N__42948\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101100"
        )
    port map (
            in0 => \N__42978\,
            in1 => \N__42521\,
            in2 => \N__49887\,
            in3 => \N__47611\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQENQL1_9_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47822\,
            in2 => \_gnd_net_\,
            in3 => \N__38754\,
            lcout => \elapsed_time_ns_1_RNIQENQL1_0_9\,
            ltout => \elapsed_time_ns_1_RNIQENQL1_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111000"
        )
    port map (
            in0 => \N__42834\,
            in1 => \N__49817\,
            in2 => \N__38757\,
            in3 => \N__47610\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_10_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__40864\,
            in1 => \N__49584\,
            in2 => \N__42267\,
            in3 => \N__46813\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49151\,
            ce => \N__48803\,
            sr => \N__48462\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50386\,
            in2 => \N__47538\,
            in3 => \N__49583\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49151\,
            ce => \N__48803\,
            sr => \N__48462\
        );

    \phase_controller_inst1.stoper_tr.target_time_5_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__49582\,
            in1 => \N__49382\,
            in2 => \N__46551\,
            in3 => \N__50392\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49151\,
            ce => \N__48803\,
            sr => \N__48462\
        );

    \phase_controller_inst1.stoper_tr.target_time_15_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__46886\,
            in1 => \N__49585\,
            in2 => \N__42408\,
            in3 => \N__46814\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49151\,
            ce => \N__48803\,
            sr => \N__48462\
        );

    \phase_controller_inst1.stoper_tr.target_time_8_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__49581\,
            in1 => \N__47886\,
            in2 => \_gnd_net_\,
            in3 => \N__50393\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49151\,
            ce => \N__48803\,
            sr => \N__48462\
        );

    \phase_controller_inst1.stoper_tr.target_time_14_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__42168\,
            in1 => \N__46812\,
            in2 => \N__49599\,
            in3 => \N__40865\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49151\,
            ce => \N__48803\,
            sr => \N__48462\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38947\,
            in1 => \N__49266\,
            in2 => \N__38931\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_15_20_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46644\,
            in2 => \N__38910\,
            in3 => \N__38921\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45057\,
            in2 => \N__38889\,
            in3 => \N__38900\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46656\,
            in2 => \N__38868\,
            in3 => \N__38879\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38858\,
            in1 => \N__38847\,
            in2 => \N__38841\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46617\,
            in2 => \N__39153\,
            in3 => \N__39168\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39123\,
            in2 => \N__39144\,
            in3 => \N__39134\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39116\,
            in1 => \N__39096\,
            in2 => \N__39105\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39089\,
            in1 => \N__40359\,
            in2 => \N__39078\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_15_21_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39068\,
            in1 => \N__39057\,
            in2 => \N__39045\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39036\,
            in2 => \N__39009\,
            in3 => \N__39020\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40785\,
            in2 => \N__38988\,
            in3 => \N__38999\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40377\,
            in2 => \N__38967\,
            in3 => \N__38978\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39258\,
            in2 => \N__39237\,
            in3 => \N__39248\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39204\,
            in2 => \N__39228\,
            in3 => \N__39215\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39435\,
            in2 => \N__39393\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39366\,
            in2 => \N__39543\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_22_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39198\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39189\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39177\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39588\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39267\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39360\,
            in2 => \N__39303\,
            in3 => \N__39462\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39459\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011010100"
        )
    port map (
            in0 => \N__39406\,
            in1 => \N__40775\,
            in2 => \N__39378\,
            in3 => \N__39426\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100110001"
        )
    port map (
            in0 => \N__39425\,
            in1 => \N__39407\,
            in2 => \N__40779\,
            in3 => \N__39374\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_17_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__49580\,
            in1 => \N__42525\,
            in2 => \_gnd_net_\,
            in3 => \N__46824\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49130\,
            ce => \N__48804\,
            sr => \N__48496\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__40745\,
            in1 => \N__39577\,
            in2 => \N__40766\,
            in3 => \N__39559\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39354\,
            in2 => \_gnd_net_\,
            in3 => \N__39322\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39290\,
            in2 => \_gnd_net_\,
            in3 => \N__39278\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_df28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__39611\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39599\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_df26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_15_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__40746\,
            in1 => \N__39578\,
            in2 => \N__40767\,
            in3 => \N__39560\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45409\,
            in1 => \N__45988\,
            in2 => \N__40130\,
            in3 => \N__40979\,
            lcout => \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__40943\,
            in1 => \N__45410\,
            in2 => \N__46013\,
            in3 => \N__39524\,
            lcout => \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__39941\,
            in1 => \N__44038\,
            in2 => \_gnd_net_\,
            in3 => \N__41009\,
            lcout => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39940\,
            lcout => \current_shift_inst.un4_control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__39523\,
            in1 => \N__44040\,
            in2 => \_gnd_net_\,
            in3 => \N__40942\,
            lcout => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44041\,
            in1 => \N__40703\,
            in2 => \_gnd_net_\,
            in3 => \N__41251\,
            lcout => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__40123\,
            in1 => \N__44039\,
            in2 => \_gnd_net_\,
            in3 => \N__40978\,
            lcout => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \N__45986\,
            in1 => \N__41149\,
            in2 => \N__39684\,
            in3 => \N__45411\,
            lcout => \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__45412\,
            in1 => \N__39681\,
            in2 => \N__41156\,
            in3 => \N__45987\,
            lcout => \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43488\,
            lcout => \current_shift_inst.un4_control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44802\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__43683\,
            in1 => \N__44047\,
            in2 => \_gnd_net_\,
            in3 => \N__43642\,
            lcout => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44049\,
            in1 => \N__46095\,
            in2 => \_gnd_net_\,
            in3 => \N__46045\,
            lcout => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__43456\,
            in1 => \N__44048\,
            in2 => \_gnd_net_\,
            in3 => \N__43489\,
            lcout => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44050\,
            in1 => \N__43773\,
            in2 => \_gnd_net_\,
            in3 => \N__43736\,
            lcout => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__43313\,
            in1 => \N__44045\,
            in2 => \_gnd_net_\,
            in3 => \N__43327\,
            lcout => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44046\,
            in1 => \_gnd_net_\,
            in2 => \N__44812\,
            in3 => \N__44773\,
            lcout => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44022\,
            in1 => \_gnd_net_\,
            in2 => \N__46273\,
            in3 => \N__46231\,
            lcout => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__44212\,
            in1 => \N__44019\,
            in2 => \_gnd_net_\,
            in3 => \N__44236\,
            lcout => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__45345\,
            in1 => \N__45876\,
            in2 => \N__45122\,
            in3 => \N__45095\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__45094\,
            in1 => \N__44021\,
            in2 => \_gnd_net_\,
            in3 => \N__45115\,
            lcout => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44017\,
            in1 => \N__43607\,
            in2 => \_gnd_net_\,
            in3 => \N__43553\,
            lcout => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__46189\,
            in1 => \N__44018\,
            in2 => \_gnd_net_\,
            in3 => \N__46138\,
            lcout => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44023\,
            in1 => \N__44994\,
            in2 => \_gnd_net_\,
            in3 => \N__44956\,
            lcout => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__44671\,
            in1 => \N__44020\,
            in2 => \_gnd_net_\,
            in3 => \N__44626\,
            lcout => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45301\,
            in1 => \N__39863\,
            in2 => \N__45974\,
            in3 => \N__41357\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__41358\,
            in1 => \N__45300\,
            in2 => \N__39864\,
            in3 => \N__45848\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45299\,
            in1 => \N__39859\,
            in2 => \_gnd_net_\,
            in3 => \N__41356\,
            lcout => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45302\,
            in2 => \_gnd_net_\,
            in3 => \N__45844\,
            lcout => \current_shift_inst.un38_control_input_axb_31_s0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45297\,
            in1 => \N__39806\,
            in2 => \N__45975\,
            in3 => \N__41549\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__41550\,
            in1 => \N__45298\,
            in2 => \N__39807\,
            in3 => \N__45852\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44024\,
            in1 => \N__39802\,
            in2 => \_gnd_net_\,
            in3 => \N__41548\,
            lcout => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__39980\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49218\,
            ce => \N__44134\,
            sr => \N__48399\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__45251\,
            in1 => \N__45672\,
            in2 => \N__41390\,
            in3 => \N__40415\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45392\,
            in1 => \N__40414\,
            in2 => \_gnd_net_\,
            in3 => \N__41383\,
            lcout => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39987\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49209\,
            ce => \N__44132\,
            sr => \N__48401\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__45673\,
            in1 => \N__45250\,
            in2 => \N__39951\,
            in3 => \N__41018\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110100011"
        )
    port map (
            in0 => \N__41019\,
            in1 => \N__39947\,
            in2 => \N__45364\,
            in3 => \N__45674\,
            lcout => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__39915\,
            in1 => \N__40668\,
            in2 => \_gnd_net_\,
            in3 => \N__45249\,
            lcout => \current_shift_inst.un38_control_input_cry_0_s0_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41063\,
            lcout => \current_shift_inst.un4_control_input1_1\,
            ltout => \current_shift_inst.un4_control_input1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45245\,
            in2 => \N__39909\,
            in3 => \N__40667\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__45805\,
            in1 => \N__45339\,
            in2 => \N__43428\,
            in3 => \N__43386\,
            lcout => \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45341\,
            in1 => \N__45803\,
            in2 => \N__46112\,
            in3 => \N__46056\,
            lcout => \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__44900\,
            in1 => \N__45343\,
            in2 => \_gnd_net_\,
            in3 => \N__44858\,
            lcout => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__45344\,
            in1 => \N__45801\,
            in2 => \N__44862\,
            in3 => \N__44901\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__45802\,
            in1 => \N__45340\,
            in2 => \N__43503\,
            in3 => \N__43464\,
            lcout => \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__41657\,
            in1 => \N__44051\,
            in2 => \_gnd_net_\,
            in3 => \N__41701\,
            lcout => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__45804\,
            in1 => \N__45338\,
            in2 => \N__40134\,
            in3 => \N__40986\,
            lcout => \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__45342\,
            in1 => \N__40222\,
            in2 => \_gnd_net_\,
            in3 => \N__41431\,
            lcout => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40072\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000101"
        )
    port map (
            in0 => \N__40223\,
            in1 => \N__45679\,
            in2 => \N__45444\,
            in3 => \N__41438\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__40256\,
            in1 => \N__45399\,
            in2 => \N__45874\,
            in3 => \N__41480\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45397\,
            in1 => \N__45685\,
            in2 => \N__44220\,
            in3 => \N__44247\,
            lcout => \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__46193\,
            in1 => \N__45396\,
            in2 => \N__45875\,
            in3 => \N__46146\,
            lcout => \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45398\,
            in1 => \N__45675\,
            in2 => \N__45006\,
            in3 => \N__44964\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__45681\,
            in1 => \N__45395\,
            in2 => \N__41781\,
            in3 => \N__41739\,
            lcout => \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45394\,
            in1 => \N__45680\,
            in2 => \N__44829\,
            in3 => \N__44781\,
            lcout => \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40320\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110011"
        )
    port map (
            in0 => \N__45980\,
            in1 => \N__40260\,
            in2 => \N__41484\,
            in3 => \N__45406\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__45407\,
            in1 => \N__45981\,
            in2 => \N__41442\,
            in3 => \N__40224\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__41708\,
            in1 => \N__45405\,
            in2 => \N__46012\,
            in3 => \N__41661\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__45982\,
            in1 => \N__45404\,
            in2 => \N__43563\,
            in3 => \N__43603\,
            lcout => \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__40433\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44576\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110011"
        )
    port map (
            in0 => \N__45976\,
            in1 => \N__40419\,
            in2 => \N__41397\,
            in3 => \N__45408\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__49874\,
            in1 => \N__42735\,
            in2 => \N__42204\,
            in3 => \N__49700\,
            lcout => \elapsed_time_ns_1_RNISAHF91_0_13\,
            ltout => \elapsed_time_ns_1_RNISAHF91_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_13_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__40831\,
            in1 => \N__49574\,
            in2 => \N__40380\,
            in3 => \N__46766\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49187\,
            ce => \N__48819\,
            sr => \N__48419\
        );

    \phase_controller_inst1.stoper_tr.target_time_9_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__42128\,
            in1 => \N__40365\,
            in2 => \N__40858\,
            in3 => \N__46767\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49187\,
            ce => \N__48819\,
            sr => \N__48419\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__40506\,
            in1 => \N__43155\,
            in2 => \N__49876\,
            in3 => \N__49696\,
            lcout => \elapsed_time_ns_1_RNI1HIF91_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__42870\,
            in1 => \N__40494\,
            in2 => \N__49711\,
            in3 => \N__49845\,
            lcout => \elapsed_time_ns_1_RNISBIF91_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__42579\,
            in1 => \N__49839\,
            in2 => \N__43227\,
            in3 => \N__49691\,
            lcout => \elapsed_time_ns_1_RNIUDIF91_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__49690\,
            in1 => \N__42230\,
            in2 => \N__49875\,
            in3 => \N__42759\,
            lcout => \elapsed_time_ns_1_RNIR9HF91_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__49840\,
            in1 => \N__40512\,
            in2 => \N__43203\,
            in3 => \N__49692\,
            lcout => \elapsed_time_ns_1_RNIVEIF91_0_25\,
            ltout => \elapsed_time_ns_1_RNIVEIF91_0_25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6_15_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40481\,
            in1 => \N__40505\,
            in2 => \N__40497\,
            in3 => \N__40469\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_o5_15_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40493\,
            in1 => \N__42345\,
            in2 => \N__40485\,
            in3 => \N__42567\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__40482\,
            in1 => \N__49841\,
            in2 => \N__49710\,
            in3 => \N__43131\,
            lcout => \elapsed_time_ns_1_RNI2IIF91_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_9_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__42105\,
            in1 => \N__46860\,
            in2 => \_gnd_net_\,
            in3 => \N__42158\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__40617\,
            in1 => \N__49961\,
            in2 => \N__40635\,
            in3 => \N__40539\,
            lcout => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\,
            ltout => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__40470\,
            in1 => \N__49701\,
            in2 => \N__40473\,
            in3 => \N__43176\,
            lcout => \elapsed_time_ns_1_RNI0GIF91_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIA965M1_18_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__40458\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47826\,
            lcout => \elapsed_time_ns_1_RNIA965M1_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9865M1_17_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__47827\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40452\,
            lcout => \elapsed_time_ns_1_RNI9865M1_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8765M1_16_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42456\,
            in2 => \_gnd_net_\,
            in3 => \N__47828\,
            lcout => \elapsed_time_ns_1_RNI8765M1_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001100"
        )
    port map (
            in0 => \N__40563\,
            in1 => \N__40545\,
            in2 => \N__49967\,
            in3 => \N__42678\,
            lcout => \delay_measurement_inst.delay_tr9\,
            ltout => \delay_measurement_inst.delay_tr9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_15_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__48585\,
            in1 => \N__40587\,
            in2 => \N__40548\,
            in3 => \N__40538\,
            lcout => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_21_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__42889\,
            in1 => \N__42868\,
            in2 => \_gnd_net_\,
            in3 => \N__40604\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_17_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__42714\,
            in1 => \N__42974\,
            in2 => \N__42708\,
            in3 => \N__40596\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_390\,
            ltout => \delay_measurement_inst.delay_tr_timer.N_390_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_17_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40530\,
            in3 => \N__40631\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.N_391_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__48586\,
            in1 => \N__49962\,
            in2 => \N__40527\,
            in3 => \N__40616\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6565M1_14_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40524\,
            in3 => \N__40518\,
            lcout => \elapsed_time_ns_1_RNI6565M1_0_14\,
            ltout => \elapsed_time_ns_1_RNI6565M1_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111000"
        )
    port map (
            in0 => \N__43068\,
            in1 => \N__49818\,
            in2 => \N__40521\,
            in3 => \N__47615\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAPC7_21_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__42890\,
            in1 => \N__40605\,
            in2 => \N__40586\,
            in3 => \N__42869\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_382\,
            ltout => \delay_measurement_inst.delay_tr_timer.N_382_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_1_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__42696\,
            in1 => \_gnd_net_\,
            in2 => \N__40620\,
            in3 => \N__42442\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_371\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQVV04_24_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40884\,
            in1 => \N__43220\,
            in2 => \N__43199\,
            in3 => \N__40569\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_356\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__43062\,
            in1 => \N__46344\,
            in2 => \N__42829\,
            in3 => \N__40559\,
            lcout => \delay_measurement_inst.N_363\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4DNE1_16_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__46345\,
            in1 => \N__47735\,
            in2 => \N__43007\,
            in3 => \N__42941\,
            lcout => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42728\,
            in1 => \N__42773\,
            in2 => \N__42755\,
            in3 => \N__42791\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_351\,
            ltout => \delay_measurement_inst.delay_tr_timer.N_351_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_15_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__43024\,
            in1 => \_gnd_net_\,
            in2 => \N__40590\,
            in3 => \N__42672\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIK0B1_23_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__43088\,
            in1 => \N__43109\,
            in2 => \_gnd_net_\,
            in3 => \N__43241\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__42940\,
            in1 => \N__42967\,
            in2 => \N__43006\,
            in3 => \N__47728\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40923\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH8AP1_20_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43124\,
            in1 => \N__43169\,
            in2 => \N__43151\,
            in3 => \N__42908\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_12_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__49576\,
            in1 => \N__42234\,
            in2 => \N__40872\,
            in3 => \N__46822\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49141\,
            ce => \N__48820\,
            sr => \N__48475\
        );

    \phase_controller_inst1.stoper_tr.target_time_16_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__49575\,
            in1 => \N__46484\,
            in2 => \_gnd_net_\,
            in3 => \N__46821\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49141\,
            ce => \N__48820\,
            sr => \N__48475\
        );

    \phase_controller_inst1.stoper_tr.target_time_19_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__46820\,
            in1 => \N__47783\,
            in2 => \_gnd_net_\,
            in3 => \N__49577\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49141\,
            ce => \N__48820\,
            sr => \N__48475\
        );

    \phase_controller_inst1.stoper_tr.target_time_18_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__49578\,
            in1 => \N__42561\,
            in2 => \_gnd_net_\,
            in3 => \N__46819\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49136\,
            ce => \N__48801\,
            sr => \N__48483\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_17_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40733\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49244\,
            ce => \N__44136\,
            sr => \N__48391\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44898\,
            lcout => \current_shift_inst.un4_control_input_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_17_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45424\,
            in1 => \N__46006\,
            in2 => \N__40707\,
            in3 => \N__41252\,
            lcout => \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_17_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40651\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_17_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45427\,
            in1 => \N__46004\,
            in2 => \N__46277\,
            in3 => \N__46236\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_17_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46269\,
            lcout => \current_shift_inst.un4_control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44998\,
            lcout => \current_shift_inst.un4_control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_17_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46007\,
            in1 => \N__45425\,
            in2 => \N__41102\,
            in3 => \N__41203\,
            lcout => \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_17_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45426\,
            in1 => \N__46005\,
            in2 => \N__43700\,
            in3 => \N__43647\,
            lcout => \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43512\,
            in2 => \N__41056\,
            in3 => \N__41049\,
            lcout => \current_shift_inst.un4_control_input1_2\,
            ltout => OPEN,
            carryin => \bfn_17_7_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41028\,
            in2 => \_gnd_net_\,
            in3 => \N__40998\,
            lcout => \current_shift_inst.un4_control_input1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_1\,
            carryout => \current_shift_inst.un4_control_input_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40995\,
            in2 => \_gnd_net_\,
            in3 => \N__40962\,
            lcout => \current_shift_inst.un4_control_input1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_2\,
            carryout => \current_shift_inst.un4_control_input_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40959\,
            in2 => \_gnd_net_\,
            in3 => \N__40926\,
            lcout => \current_shift_inst.un4_control_input1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_3\,
            carryout => \current_shift_inst.un4_control_input_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41265\,
            in2 => \_gnd_net_\,
            in3 => \N__41235\,
            lcout => \current_shift_inst.un4_control_input1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_4\,
            carryout => \current_shift_inst.un4_control_input_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41232\,
            in2 => \_gnd_net_\,
            in3 => \N__41220\,
            lcout => \current_shift_inst.un4_control_input1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_5\,
            carryout => \current_shift_inst.un4_control_input_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41217\,
            in2 => \_gnd_net_\,
            in3 => \N__41184\,
            lcout => \current_shift_inst.un4_control_input1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_6\,
            carryout => \current_shift_inst.un4_control_input_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41181\,
            in2 => \_gnd_net_\,
            in3 => \N__41172\,
            lcout => \current_shift_inst.un4_control_input1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_7\,
            carryout => \current_shift_inst.un4_control_input_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41169\,
            in2 => \_gnd_net_\,
            in3 => \N__41133\,
            lcout => \current_shift_inst.un4_control_input1_10\,
            ltout => OPEN,
            carryin => \bfn_17_8_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41130\,
            in2 => \_gnd_net_\,
            in3 => \N__41124\,
            lcout => \current_shift_inst.un4_control_input1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_9\,
            carryout => \current_shift_inst.un4_control_input_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41121\,
            in2 => \_gnd_net_\,
            in3 => \N__41109\,
            lcout => \current_shift_inst.un4_control_input1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_10\,
            carryout => \current_shift_inst.un4_control_input_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43521\,
            in3 => \N__41106\,
            lcout => \current_shift_inst.un4_control_input1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_11\,
            carryout => \current_shift_inst.un4_control_input_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41343\,
            in2 => \_gnd_net_\,
            in3 => \N__41337\,
            lcout => \current_shift_inst.un4_control_input1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_12\,
            carryout => \current_shift_inst.un4_control_input_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43344\,
            in2 => \_gnd_net_\,
            in3 => \N__41334\,
            lcout => \current_shift_inst.un4_control_input1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_13\,
            carryout => \current_shift_inst.un4_control_input_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41331\,
            in2 => \_gnd_net_\,
            in3 => \N__41319\,
            lcout => \current_shift_inst.un4_control_input1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_14\,
            carryout => \current_shift_inst.un4_control_input_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41316\,
            in2 => \_gnd_net_\,
            in3 => \N__41307\,
            lcout => \current_shift_inst.un4_control_input1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_15\,
            carryout => \current_shift_inst.un4_control_input_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41304\,
            in2 => \_gnd_net_\,
            in3 => \N__41295\,
            lcout => \current_shift_inst.un4_control_input1_18\,
            ltout => OPEN,
            carryin => \bfn_17_9_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41292\,
            in2 => \_gnd_net_\,
            in3 => \N__41283\,
            lcout => \current_shift_inst.un4_control_input1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_17\,
            carryout => \current_shift_inst.un4_control_input_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41280\,
            in2 => \_gnd_net_\,
            in3 => \N__41271\,
            lcout => \current_shift_inst.un4_control_input1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_18\,
            carryout => \current_shift_inst.un4_control_input_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46200\,
            in2 => \_gnd_net_\,
            in3 => \N__41268\,
            lcout => \current_shift_inst.un4_control_input1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_19\,
            carryout => \current_shift_inst.un4_control_input_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41559\,
            in2 => \_gnd_net_\,
            in3 => \N__41538\,
            lcout => \current_shift_inst.un4_control_input1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_20\,
            carryout => \current_shift_inst.un4_control_input_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41535\,
            in2 => \_gnd_net_\,
            in3 => \N__41526\,
            lcout => \current_shift_inst.un4_control_input1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_21\,
            carryout => \current_shift_inst.un4_control_input_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41523\,
            in2 => \_gnd_net_\,
            in3 => \N__41514\,
            lcout => \current_shift_inst.un4_control_input1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_22\,
            carryout => \current_shift_inst.un4_control_input_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41511\,
            in2 => \_gnd_net_\,
            in3 => \N__41496\,
            lcout => \current_shift_inst.un4_control_input1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_23\,
            carryout => \current_shift_inst.un4_control_input_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41493\,
            in2 => \_gnd_net_\,
            in3 => \N__41454\,
            lcout => \current_shift_inst.un4_control_input1_26\,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41451\,
            in2 => \_gnd_net_\,
            in3 => \N__41409\,
            lcout => \current_shift_inst.un4_control_input1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_25\,
            carryout => \current_shift_inst.un4_control_input_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41406\,
            in2 => \_gnd_net_\,
            in3 => \N__41370\,
            lcout => \current_shift_inst.un4_control_input1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_26\,
            carryout => \current_shift_inst.un4_control_input_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41367\,
            in2 => \_gnd_net_\,
            in3 => \N__41346\,
            lcout => \current_shift_inst.un4_control_input1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_27\,
            carryout => \current_shift_inst.un4_control_input_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41796\,
            in2 => \_gnd_net_\,
            in3 => \N__41787\,
            lcout => \current_shift_inst.un4_control_input1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_28\,
            carryout => \current_shift_inst.un4_control_input1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41784\,
            lcout => \current_shift_inst.un4_control_input1_31_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45266\,
            in1 => \N__45942\,
            in2 => \N__41780\,
            in3 => \N__41734\,
            lcout => \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__45941\,
            in1 => \N__45267\,
            in2 => \N__41709\,
            in3 => \N__41656\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41637\,
            in2 => \N__41612\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_11_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44093\,
            in2 => \N__44070\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45888\,
            in2 => \N__41595\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41586\,
            in2 => \N__45993\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45892\,
            in2 => \N__41574\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41847\,
            in2 => \N__45994\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45896\,
            in2 => \N__43359\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41838\,
            in2 => \N__45995\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45751\,
            in2 => \N__43281\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_12_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41829\,
            in2 => \N__45907\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45755\,
            in2 => \N__44757\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41817\,
            in2 => \N__45908\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45759\,
            in2 => \N__41808\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43440\,
            in2 => \N__45909\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45763\,
            in2 => \N__46029\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43713\,
            in2 => \N__45910\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45911\,
            in2 => \N__43536\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_13_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46122\,
            in2 => \N__45996\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45915\,
            in2 => \N__44178\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44610\,
            in2 => \N__45997\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45919\,
            in2 => \N__45072\,
            in3 => \N__41874\,
            lcout => \current_shift_inst.un38_control_input_0_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41871\,
            in2 => \N__45998\,
            in3 => \N__41850\,
            lcout => \current_shift_inst.un38_control_input_0_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45923\,
            in2 => \N__42078\,
            in3 => \N__42051\,
            lcout => \current_shift_inst.un38_control_input_0_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44940\,
            in2 => \N__45999\,
            in3 => \N__42036\,
            lcout => \current_shift_inst.un38_control_input_0_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45927\,
            in2 => \N__42033\,
            in3 => \N__42009\,
            lcout => \current_shift_inst.un38_control_input_0_s1_24\,
            ltout => OPEN,
            carryin => \bfn_17_14_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42006\,
            in2 => \N__46000\,
            in3 => \N__41988\,
            lcout => \current_shift_inst.un38_control_input_0_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45931\,
            in2 => \N__41985\,
            in3 => \N__41961\,
            lcout => \current_shift_inst.un38_control_input_0_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41958\,
            in2 => \N__46001\,
            in3 => \N__41934\,
            lcout => \current_shift_inst.un38_control_input_0_s1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45935\,
            in2 => \N__41931\,
            in3 => \N__41904\,
            lcout => \current_shift_inst.un38_control_input_0_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44841\,
            in2 => \N__46002\,
            in3 => \N__41889\,
            lcout => \current_shift_inst.un38_control_input_0_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45939\,
            in2 => \N__43869\,
            in3 => \N__42288\,
            lcout => \current_shift_inst.un38_control_input_0_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__45940\,
            in1 => \N__45403\,
            in2 => \_gnd_net_\,
            in3 => \N__42285\,
            lcout => \current_shift_inst.un38_control_input_0_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__49861\,
            in1 => \N__49686\,
            in2 => \N__42253\,
            in3 => \N__42795\,
            lcout => \elapsed_time_ns_1_RNIP7HF91_0_10\,
            ltout => \elapsed_time_ns_1_RNIP7HF91_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_2_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42225\,
            in1 => \N__42199\,
            in2 => \N__42183\,
            in3 => \N__42321\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_6_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42169\,
            in2 => \N__42132\,
            in3 => \N__42127\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_6_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111010"
        )
    port map (
            in0 => \N__42388\,
            in1 => \N__46867\,
            in2 => \N__42087\,
            in3 => \N__46727\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC8TA1_3_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111101100"
        )
    port map (
            in0 => \N__49863\,
            in1 => \N__47842\,
            in2 => \N__42660\,
            in3 => \N__46427\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK8NQL1_3_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42084\,
            in3 => \N__47668\,
            lcout => \elapsed_time_ns_1_RNIK8NQL1_0_3\,
            ltout => \elapsed_time_ns_1_RNIK8NQL1_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2_1_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42081\,
            in3 => \N__46399\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__46400\,
            in1 => \N__49862\,
            in2 => \N__49709\,
            in3 => \N__50013\,
            lcout => \elapsed_time_ns_1_RNIAE2591_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__49679\,
            in1 => \N__49814\,
            in2 => \N__42363\,
            in3 => \N__42894\,
            lcout => \elapsed_time_ns_1_RNIRAIF91_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110100"
        )
    port map (
            in0 => \N__42449\,
            in1 => \N__48584\,
            in2 => \N__42423\,
            in3 => \N__49951\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\,
            ltout => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__46874\,
            in1 => \N__43038\,
            in2 => \N__42414\,
            in3 => \N__49816\,
            lcout => \elapsed_time_ns_1_RNIUCHF91_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBA65M1_19_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47841\,
            in2 => \_gnd_net_\,
            in3 => \N__47715\,
            lcout => \elapsed_time_ns_1_RNIBA65M1_0_19\,
            ltout => \elapsed_time_ns_1_RNIBA65M1_0_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_9_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__42554\,
            in1 => \N__42515\,
            in2 => \N__42411\,
            in3 => \N__46472\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__49813\,
            in1 => \N__42372\,
            in2 => \N__42918\,
            in3 => \N__49678\,
            lcout => \elapsed_time_ns_1_RNIQ9IF91_0_20\,
            ltout => \elapsed_time_ns_1_RNIQ9IF91_0_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7_15_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42599\,
            in1 => \N__42467\,
            in2 => \N__42366\,
            in3 => \N__42356\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__49815\,
            in1 => \N__42777\,
            in2 => \N__42335\,
            in3 => \N__49680\,
            lcout => \elapsed_time_ns_1_RNIQ8HF91_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__49682\,
            in1 => \N__49820\,
            in2 => \N__42603\,
            in3 => \N__43110\,
            lcout => \elapsed_time_ns_1_RNI3JIF91_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__49819\,
            in1 => \N__42588\,
            in2 => \N__43248\,
            in3 => \N__49681\,
            lcout => \elapsed_time_ns_1_RNITCIF91_0_23\,
            ltout => \elapsed_time_ns_1_RNITCIF91_0_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_15_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42582\,
            in3 => \N__42578\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__50416\,
            in1 => \N__42639\,
            in2 => \N__49864\,
            in3 => \N__49684\,
            lcout => \elapsed_time_ns_1_RNICG2591_0_4\,
            ltout => \elapsed_time_ns_1_RNICG2591_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3_2_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__47766\,
            in1 => \N__42555\,
            in2 => \N__42528\,
            in3 => \N__46536\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_2_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__42516\,
            in1 => \N__42485\,
            in2 => \N__42474\,
            in3 => \N__46473\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__49683\,
            in1 => \N__49821\,
            in2 => \N__42471\,
            in3 => \N__43089\,
            lcout => \elapsed_time_ns_1_RNIRBJF91_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__46537\,
            in1 => \N__42621\,
            in2 => \N__49865\,
            in3 => \N__49685\,
            lcout => \elapsed_time_ns_1_RNIDH2591_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101100"
        )
    port map (
            in0 => \N__43008\,
            in1 => \N__46480\,
            in2 => \N__49886\,
            in3 => \N__47626\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNINAPP_2_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__42653\,
            in1 => \N__50009\,
            in2 => \N__42830\,
            in3 => \N__43066\,
            lcout => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42617\,
            in2 => \_gnd_net_\,
            in3 => \N__42635\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_344\,
            ltout => \delay_measurement_inst.delay_tr_timer.N_344_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42652\,
            in1 => \N__50008\,
            in2 => \N__42699\,
            in3 => \N__50054\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_347\,
            ltout => \delay_measurement_inst.delay_tr_timer.N_347_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQMF21_6_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010000000"
        )
    port map (
            in0 => \N__42825\,
            in1 => \N__46346\,
            in2 => \N__42690\,
            in3 => \N__42671\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.N_373_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNID68O3_15_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101010"
        )
    port map (
            in0 => \N__43037\,
            in1 => \N__43067\,
            in2 => \N__42687\,
            in3 => \N__42684\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_353\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47897\,
            in2 => \_gnd_net_\,
            in3 => \N__45032\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_348\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46594\,
            in2 => \N__50081\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_17_19_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__49165\,
            ce => \N__49985\,
            sr => \N__48446\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46570\,
            in2 => \N__50036\,
            in3 => \N__42624\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__49165\,
            ce => \N__49985\,
            sr => \N__48446\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47077\,
            in2 => \N__46599\,
            in3 => \N__42606\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__49165\,
            ce => \N__49985\,
            sr => \N__48446\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47053\,
            in2 => \N__46575\,
            in3 => \N__42843\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__49165\,
            ce => \N__49985\,
            sr => \N__48446\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47029\,
            in2 => \N__47082\,
            in3 => \N__42840\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__49165\,
            ce => \N__49985\,
            sr => \N__48446\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47005\,
            in2 => \N__47058\,
            in3 => \N__42837\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__49165\,
            ce => \N__49985\,
            sr => \N__48446\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46981\,
            in2 => \N__47034\,
            in3 => \N__42798\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__49165\,
            ce => \N__49985\,
            sr => \N__48446\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46957\,
            in2 => \N__47010\,
            in3 => \N__42780\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__49165\,
            ce => \N__49985\,
            sr => \N__48446\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46933\,
            in2 => \N__46986\,
            in3 => \N__42762\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_17_20_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__49157\,
            ce => \N__49986\,
            sr => \N__48456\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46909\,
            in2 => \N__46962\,
            in3 => \N__42738\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__49157\,
            ce => \N__49986\,
            sr => \N__48456\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47293\,
            in2 => \N__46938\,
            in3 => \N__42717\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__49157\,
            ce => \N__49986\,
            sr => \N__48456\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47269\,
            in2 => \N__46914\,
            in3 => \N__43041\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__49157\,
            ce => \N__49986\,
            sr => \N__48456\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47245\,
            in2 => \N__47298\,
            in3 => \N__43011\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__49157\,
            ce => \N__49986\,
            sr => \N__48456\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47221\,
            in2 => \N__47274\,
            in3 => \N__42981\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__49157\,
            ce => \N__49986\,
            sr => \N__48456\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47197\,
            in2 => \N__47250\,
            in3 => \N__42951\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__49157\,
            ce => \N__49986\,
            sr => \N__48456\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47173\,
            in2 => \N__47226\,
            in3 => \N__42924\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__49157\,
            ce => \N__49986\,
            sr => \N__48456\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47149\,
            in2 => \N__47202\,
            in3 => \N__42921\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_17_21_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__49152\,
            ce => \N__49987\,
            sr => \N__48463\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47125\,
            in2 => \N__47178\,
            in3 => \N__42897\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__49152\,
            ce => \N__49987\,
            sr => \N__48463\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47101\,
            in2 => \N__47154\,
            in3 => \N__42873\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__49152\,
            ce => \N__49987\,
            sr => \N__48463\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47476\,
            in2 => \N__47130\,
            in3 => \N__42846\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__49152\,
            ce => \N__49987\,
            sr => \N__48463\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47452\,
            in2 => \N__47106\,
            in3 => \N__43230\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__49152\,
            ce => \N__49987\,
            sr => \N__48463\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47428\,
            in2 => \N__47481\,
            in3 => \N__43206\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__49152\,
            ce => \N__49987\,
            sr => \N__48463\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47404\,
            in2 => \N__47457\,
            in3 => \N__43179\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__49152\,
            ce => \N__49987\,
            sr => \N__48463\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47380\,
            in2 => \N__47433\,
            in3 => \N__43158\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__49152\,
            ce => \N__49987\,
            sr => \N__48463\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47356\,
            in2 => \N__47409\,
            in3 => \N__43134\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_17_22_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__49147\,
            ce => \N__49989\,
            sr => \N__48469\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47332\,
            in2 => \N__47385\,
            in3 => \N__43113\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__49147\,
            ce => \N__49989\,
            sr => \N__48469\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_17_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47312\,
            in2 => \N__47361\,
            in3 => \N__43092\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__49147\,
            ce => \N__49989\,
            sr => \N__48469\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47957\,
            in2 => \N__47337\,
            in3 => \N__43071\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__49147\,
            ce => \N__49989\,
            sr => \N__48469\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43611\,
            lcout => \delay_measurement_inst.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49147\,
            ce => \N__49989\,
            sr => \N__48469\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_18_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46009\,
            in1 => \N__45431\,
            in2 => \N__43608\,
            in3 => \N__43552\,
            lcout => \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43693\,
            lcout => \current_shift_inst.un4_control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43914\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_18_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46008\,
            in1 => \N__45430\,
            in2 => \N__43502\,
            in3 => \N__43457\,
            lcout => \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_18_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45428\,
            in1 => \N__46010\,
            in2 => \N__43421\,
            in3 => \N__43378\,
            lcout => \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_18_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46105\,
            lcout => \current_shift_inst.un4_control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_18_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__45429\,
            in1 => \N__46011\,
            in2 => \N__43338\,
            in3 => \N__43314\,
            lcout => \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__45413\,
            in1 => \N__43931\,
            in2 => \N__44103\,
            in3 => \N__43916\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44163\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49236\,
            ce => \N__44135\,
            sr => \N__48392\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__43917\,
            in1 => \N__45414\,
            in2 => \N__43932\,
            in3 => \N__44102\,
            lcout => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__44054\,
            in1 => \N__43927\,
            in2 => \_gnd_net_\,
            in3 => \N__43915\,
            lcout => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45415\,
            in2 => \_gnd_net_\,
            in3 => \N__43816\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__45416\,
            in1 => \N__43818\,
            in2 => \N__43854\,
            in3 => \N__45992\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \N__43850\,
            in1 => \N__45417\,
            in2 => \N__46014\,
            in3 => \N__43817\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__45954\,
            in1 => \N__45434\,
            in2 => \N__43782\,
            in3 => \N__43732\,
            lcout => \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45433\,
            in1 => \N__45953\,
            in2 => \N__43701\,
            in3 => \N__43646\,
            lcout => \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__45948\,
            in1 => \N__45436\,
            in2 => \N__45002\,
            in3 => \N__44957\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44917\,
            in2 => \_gnd_net_\,
            in3 => \N__44589\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__44899\,
            in1 => \N__45437\,
            in2 => \N__46003\,
            in3 => \N__44857\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45432\,
            in1 => \N__45952\,
            in2 => \N__44825\,
            in3 => \N__44774\,
            lcout => \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44745\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45435\,
            in1 => \N__45955\,
            in2 => \N__44675\,
            in3 => \N__44627\,
            lcout => \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44588\,
            in1 => \N__44269\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__45947\,
            in1 => \N__45439\,
            in2 => \N__44243\,
            in3 => \N__44216\,
            lcout => \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45442\,
            in1 => \N__45943\,
            in2 => \N__46281\,
            in3 => \N__46232\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45101\,
            lcout => \current_shift_inst.un4_control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__45946\,
            in1 => \N__45440\,
            in2 => \N__46194\,
            in3 => \N__46139\,
            lcout => \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__45438\,
            in1 => \N__45945\,
            in2 => \N__46113\,
            in3 => \N__46052\,
            lcout => \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__45944\,
            in1 => \N__45441\,
            in2 => \N__45126\,
            in3 => \N__45102\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_3_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__46428\,
            in1 => \N__49383\,
            in2 => \N__46386\,
            in3 => \N__50384\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49210\,
            ce => \N__48821\,
            sr => \N__48402\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__49893\,
            in1 => \N__47527\,
            in2 => \N__45042\,
            in3 => \N__49705\,
            lcout => \elapsed_time_ns_1_RNIFJ2591_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_8_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__50348\,
            in1 => \N__49538\,
            in2 => \_gnd_net_\,
            in3 => \N__47885\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49199\,
            ce => \N__50284\,
            sr => \N__48407\
        );

    \phase_controller_inst2.stoper_tr.target_time_5_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__49367\,
            in1 => \N__50349\,
            in2 => \N__49579\,
            in3 => \N__46547\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49199\,
            ce => \N__50284\,
            sr => \N__48407\
        );

    \phase_controller_inst2.stoper_tr.target_time_3_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111010101010"
        )
    port map (
            in0 => \N__46382\,
            in1 => \N__49368\,
            in2 => \N__50383\,
            in3 => \N__46423\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49199\,
            ce => \N__50284\,
            sr => \N__48407\
        );

    \phase_controller_inst2.stoper_tr.target_time_16_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__49537\,
            in1 => \N__46485\,
            in2 => \_gnd_net_\,
            in3 => \N__46818\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49199\,
            ce => \N__50284\,
            sr => \N__48407\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_0_2_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011111111"
        )
    port map (
            in0 => \N__46368\,
            in1 => \N__46422\,
            in2 => \N__46299\,
            in3 => \N__46401\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_3_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010101010"
        )
    port map (
            in0 => \N__49464\,
            in1 => \N__46294\,
            in2 => \N__46808\,
            in3 => \N__46367\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5_1_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__46366\,
            in1 => \N__46772\,
            in2 => \N__46298\,
            in3 => \N__46356\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101110"
        )
    port map (
            in0 => \N__47662\,
            in1 => \N__46630\,
            in2 => \N__49905\,
            in3 => \N__46350\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNINBNQL1_6_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__46326\,
            in3 => \N__47846\,
            lcout => \elapsed_time_ns_1_RNINBNQL1_0_6\,
            ltout => \elapsed_time_ns_1_RNINBNQL1_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_2_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__47881\,
            in1 => \N__47520\,
            in2 => \N__46323\,
            in3 => \N__46310\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_6_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46868\,
            in2 => \N__46827\,
            in3 => \N__46768\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_6_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010000000101"
        )
    port map (
            in0 => \N__49465\,
            in1 => \N__46631\,
            in2 => \N__46671\,
            in3 => \N__50385\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49194\,
            ce => \N__50280\,
            sr => \N__48414\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__49364\,
            in1 => \N__50394\,
            in2 => \N__49607\,
            in3 => \N__50420\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49188\,
            ce => \N__48811\,
            sr => \N__48420\
        );

    \phase_controller_inst1.stoper_tr.target_time_2_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001010100"
        )
    port map (
            in0 => \N__50447\,
            in1 => \N__49366\,
            in2 => \N__50400\,
            in3 => \N__49606\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49188\,
            ce => \N__48811\,
            sr => \N__48420\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__49365\,
            in1 => \N__50395\,
            in2 => \N__49608\,
            in3 => \N__46632\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49188\,
            ce => \N__48811\,
            sr => \N__48420\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48083\,
            in1 => \N__50074\,
            in2 => \_gnd_net_\,
            in3 => \N__46605\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_18_18_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__49181\,
            ce => \N__47934\,
            sr => \N__48429\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48061\,
            in1 => \N__50029\,
            in2 => \_gnd_net_\,
            in3 => \N__46602\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__49181\,
            ce => \N__47934\,
            sr => \N__48429\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48084\,
            in1 => \N__46595\,
            in2 => \_gnd_net_\,
            in3 => \N__46578\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__49181\,
            ce => \N__47934\,
            sr => \N__48429\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48062\,
            in1 => \N__46571\,
            in2 => \_gnd_net_\,
            in3 => \N__46554\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__49181\,
            ce => \N__47934\,
            sr => \N__48429\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48085\,
            in1 => \N__47078\,
            in2 => \_gnd_net_\,
            in3 => \N__47061\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__49181\,
            ce => \N__47934\,
            sr => \N__48429\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48063\,
            in1 => \N__47054\,
            in2 => \_gnd_net_\,
            in3 => \N__47037\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__49181\,
            ce => \N__47934\,
            sr => \N__48429\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48086\,
            in1 => \N__47030\,
            in2 => \_gnd_net_\,
            in3 => \N__47013\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__49181\,
            ce => \N__47934\,
            sr => \N__48429\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48064\,
            in1 => \N__47006\,
            in2 => \_gnd_net_\,
            in3 => \N__46989\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__49181\,
            ce => \N__47934\,
            sr => \N__48429\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48068\,
            in1 => \N__46982\,
            in2 => \_gnd_net_\,
            in3 => \N__46965\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_18_19_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__49173\,
            ce => \N__47945\,
            sr => \N__48435\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48076\,
            in1 => \N__46958\,
            in2 => \_gnd_net_\,
            in3 => \N__46941\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__49173\,
            ce => \N__47945\,
            sr => \N__48435\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48065\,
            in1 => \N__46934\,
            in2 => \_gnd_net_\,
            in3 => \N__46917\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__49173\,
            ce => \N__47945\,
            sr => \N__48435\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48073\,
            in1 => \N__46910\,
            in2 => \_gnd_net_\,
            in3 => \N__46893\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__49173\,
            ce => \N__47945\,
            sr => \N__48435\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48066\,
            in1 => \N__47294\,
            in2 => \_gnd_net_\,
            in3 => \N__47277\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__49173\,
            ce => \N__47945\,
            sr => \N__48435\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48074\,
            in1 => \N__47270\,
            in2 => \_gnd_net_\,
            in3 => \N__47253\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__49173\,
            ce => \N__47945\,
            sr => \N__48435\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48067\,
            in1 => \N__47246\,
            in2 => \_gnd_net_\,
            in3 => \N__47229\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__49173\,
            ce => \N__47945\,
            sr => \N__48435\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48075\,
            in1 => \N__47222\,
            in2 => \_gnd_net_\,
            in3 => \N__47205\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__49173\,
            ce => \N__47945\,
            sr => \N__48435\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48087\,
            in1 => \N__47198\,
            in2 => \_gnd_net_\,
            in3 => \N__47181\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_18_20_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__49166\,
            ce => \N__47944\,
            sr => \N__48447\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48069\,
            in1 => \N__47174\,
            in2 => \_gnd_net_\,
            in3 => \N__47157\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__49166\,
            ce => \N__47944\,
            sr => \N__48447\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48088\,
            in1 => \N__47150\,
            in2 => \_gnd_net_\,
            in3 => \N__47133\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__49166\,
            ce => \N__47944\,
            sr => \N__48447\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48070\,
            in1 => \N__47126\,
            in2 => \_gnd_net_\,
            in3 => \N__47109\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__49166\,
            ce => \N__47944\,
            sr => \N__48447\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48089\,
            in1 => \N__47102\,
            in2 => \_gnd_net_\,
            in3 => \N__47085\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__49166\,
            ce => \N__47944\,
            sr => \N__48447\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48071\,
            in1 => \N__47477\,
            in2 => \_gnd_net_\,
            in3 => \N__47460\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__49166\,
            ce => \N__47944\,
            sr => \N__48447\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48090\,
            in1 => \N__47453\,
            in2 => \_gnd_net_\,
            in3 => \N__47436\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__49166\,
            ce => \N__47944\,
            sr => \N__48447\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_18_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48072\,
            in1 => \N__47429\,
            in2 => \_gnd_net_\,
            in3 => \N__47412\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__49166\,
            ce => \N__47944\,
            sr => \N__48447\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48077\,
            in1 => \N__47405\,
            in2 => \_gnd_net_\,
            in3 => \N__47388\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_18_21_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__49158\,
            ce => \N__47946\,
            sr => \N__48457\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48081\,
            in1 => \N__47381\,
            in2 => \_gnd_net_\,
            in3 => \N__47364\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__49158\,
            ce => \N__47946\,
            sr => \N__48457\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48078\,
            in1 => \N__47357\,
            in2 => \_gnd_net_\,
            in3 => \N__47340\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__49158\,
            ce => \N__47946\,
            sr => \N__48457\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_18_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48082\,
            in1 => \N__47333\,
            in2 => \_gnd_net_\,
            in3 => \N__47316\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__49158\,
            ce => \N__47946\,
            sr => \N__48457\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48079\,
            in1 => \N__47313\,
            in2 => \_gnd_net_\,
            in3 => \N__47301\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__49158\,
            ce => \N__47946\,
            sr => \N__48457\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_18_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__47958\,
            in1 => \N__48080\,
            in2 => \_gnd_net_\,
            in3 => \N__47961\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49158\,
            ce => \N__47946\,
            sr => \N__48457\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_20_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__47871\,
            in1 => \N__49900\,
            in2 => \N__47907\,
            in3 => \N__49716\,
            lcout => \elapsed_time_ns_1_RNIGK2591_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII6NQL1_1_LC_20_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47544\,
            in2 => \_gnd_net_\,
            in3 => \N__47847\,
            lcout => \elapsed_time_ns_1_RNII6NQL1_0_1\,
            ltout => \elapsed_time_ns_1_RNII6NQL1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_1_LC_20_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101010"
        )
    port map (
            in0 => \N__49451\,
            in1 => \_gnd_net_\,
            in2 => \N__47787\,
            in3 => \N__50359\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_20_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110010"
        )
    port map (
            in0 => \N__47782\,
            in1 => \N__49888\,
            in2 => \N__47701\,
            in3 => \N__47742\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_20_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101001110"
        )
    port map (
            in0 => \N__49889\,
            in1 => \N__49315\,
            in2 => \N__50058\,
            in3 => \N__47690\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_7_LC_20_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__47537\,
            in1 => \N__49458\,
            in2 => \_gnd_net_\,
            in3 => \N__50391\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49205\,
            ce => \N__50286\,
            sr => \N__48415\
        );

    \phase_controller_inst2.stoper_tr.target_time_1_LC_20_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__49372\,
            in1 => \N__49316\,
            in2 => \N__49281\,
            in3 => \N__49298\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49205\,
            ce => \N__50286\,
            sr => \N__48415\
        );

    \phase_controller_inst2.stoper_tr.target_time_2_LC_20_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001010100"
        )
    port map (
            in0 => \N__50451\,
            in1 => \N__49374\,
            in2 => \N__50399\,
            in3 => \N__49459\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49205\,
            ce => \N__50286\,
            sr => \N__48415\
        );

    \phase_controller_inst2.stoper_tr.target_time_4_LC_20_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__49373\,
            in1 => \N__49460\,
            in2 => \N__50427\,
            in3 => \N__50390\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49205\,
            ce => \N__50286\,
            sr => \N__48415\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_20_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50082\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49195\,
            ce => \N__49988\,
            sr => \N__48430\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_20_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50037\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49195\,
            ce => \N__49988\,
            sr => \N__48430\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_21_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__49963\,
            in1 => \N__49904\,
            in2 => \N__49498\,
            in3 => \N__49715\,
            lcout => \elapsed_time_ns_1_RNISCJF91_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_1_LC_21_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__49381\,
            in1 => \N__49317\,
            in2 => \N__49299\,
            in3 => \N__49280\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49212\,
            ce => \N__48822\,
            sr => \N__48421\
        );
end \INTERFACE\;
